magic
tech sky130A
magscale 1 2
timestamp 1647558357
<< obsli1 >>
rect 1104 2159 10856 77809
<< obsm1 >>
rect 14 1028 10856 77840
<< metal2 >>
rect 5998 79200 6054 80000
<< obsm2 >>
rect 18 79144 5942 79529
rect 6110 79144 10284 79529
rect 18 167 10284 79144
<< metal3 >>
rect 0 79568 800 79688
rect 11200 79432 12000 79552
rect 0 79160 800 79280
rect 0 78752 800 78872
rect 11200 78616 12000 78736
rect 0 78344 800 78464
rect 0 77936 800 78056
rect 11200 77936 12000 78056
rect 0 77528 800 77648
rect 0 77120 800 77240
rect 11200 77120 12000 77240
rect 0 76576 800 76696
rect 0 76168 800 76288
rect 11200 76304 12000 76424
rect 0 75760 800 75880
rect 11200 75624 12000 75744
rect 0 75352 800 75472
rect 0 74944 800 75064
rect 11200 74808 12000 74928
rect 0 74536 800 74656
rect 0 74128 800 74248
rect 11200 73992 12000 74112
rect 0 73720 800 73840
rect 0 73176 800 73296
rect 11200 73312 12000 73432
rect 0 72768 800 72888
rect 0 72360 800 72480
rect 11200 72496 12000 72616
rect 0 71952 800 72072
rect 0 71544 800 71664
rect 11200 71680 12000 71800
rect 0 71136 800 71256
rect 11200 71000 12000 71120
rect 0 70728 800 70848
rect 0 70320 800 70440
rect 11200 70184 12000 70304
rect 0 69776 800 69896
rect 0 69368 800 69488
rect 11200 69368 12000 69488
rect 0 68960 800 69080
rect 0 68552 800 68672
rect 11200 68688 12000 68808
rect 0 68144 800 68264
rect 0 67736 800 67856
rect 11200 67872 12000 67992
rect 0 67328 800 67448
rect 0 66920 800 67040
rect 11200 67056 12000 67176
rect 0 66376 800 66496
rect 11200 66376 12000 66496
rect 0 65968 800 66088
rect 0 65560 800 65680
rect 11200 65560 12000 65680
rect 0 65152 800 65272
rect 0 64744 800 64864
rect 11200 64744 12000 64864
rect 0 64336 800 64456
rect 0 63928 800 64048
rect 11200 64064 12000 64184
rect 0 63520 800 63640
rect 11200 63248 12000 63368
rect 0 62976 800 63096
rect 0 62568 800 62688
rect 11200 62432 12000 62552
rect 0 62160 800 62280
rect 0 61752 800 61872
rect 11200 61752 12000 61872
rect 0 61344 800 61464
rect 0 60936 800 61056
rect 11200 60936 12000 61056
rect 0 60528 800 60648
rect 0 60120 800 60240
rect 11200 60256 12000 60376
rect 0 59576 800 59696
rect 11200 59440 12000 59560
rect 0 59168 800 59288
rect 0 58760 800 58880
rect 11200 58624 12000 58744
rect 0 58352 800 58472
rect 0 57944 800 58064
rect 11200 57944 12000 58064
rect 0 57536 800 57656
rect 0 57128 800 57248
rect 11200 57128 12000 57248
rect 0 56584 800 56704
rect 0 56176 800 56296
rect 11200 56312 12000 56432
rect 0 55768 800 55888
rect 11200 55632 12000 55752
rect 0 55360 800 55480
rect 0 54952 800 55072
rect 11200 54816 12000 54936
rect 0 54544 800 54664
rect 0 54136 800 54256
rect 11200 54000 12000 54120
rect 0 53728 800 53848
rect 0 53184 800 53304
rect 11200 53320 12000 53440
rect 0 52776 800 52896
rect 0 52368 800 52488
rect 11200 52504 12000 52624
rect 0 51960 800 52080
rect 0 51552 800 51672
rect 11200 51688 12000 51808
rect 0 51144 800 51264
rect 11200 51008 12000 51128
rect 0 50736 800 50856
rect 0 50328 800 50448
rect 11200 50192 12000 50312
rect 0 49784 800 49904
rect 0 49376 800 49496
rect 11200 49376 12000 49496
rect 0 48968 800 49088
rect 0 48560 800 48680
rect 11200 48696 12000 48816
rect 0 48152 800 48272
rect 0 47744 800 47864
rect 11200 47880 12000 48000
rect 0 47336 800 47456
rect 0 46928 800 47048
rect 11200 47064 12000 47184
rect 0 46384 800 46504
rect 11200 46384 12000 46504
rect 0 45976 800 46096
rect 0 45568 800 45688
rect 11200 45568 12000 45688
rect 0 45160 800 45280
rect 0 44752 800 44872
rect 11200 44752 12000 44872
rect 0 44344 800 44464
rect 0 43936 800 44056
rect 11200 44072 12000 44192
rect 0 43528 800 43648
rect 11200 43256 12000 43376
rect 0 42984 800 43104
rect 0 42576 800 42696
rect 11200 42440 12000 42560
rect 0 42168 800 42288
rect 0 41760 800 41880
rect 11200 41760 12000 41880
rect 0 41352 800 41472
rect 0 40944 800 41064
rect 11200 40944 12000 41064
rect 0 40536 800 40656
rect 0 40128 800 40248
rect 11200 40264 12000 40384
rect 0 39584 800 39704
rect 11200 39448 12000 39568
rect 0 39176 800 39296
rect 0 38768 800 38888
rect 11200 38632 12000 38752
rect 0 38360 800 38480
rect 0 37952 800 38072
rect 11200 37952 12000 38072
rect 0 37544 800 37664
rect 0 37136 800 37256
rect 11200 37136 12000 37256
rect 0 36592 800 36712
rect 0 36184 800 36304
rect 11200 36320 12000 36440
rect 0 35776 800 35896
rect 11200 35640 12000 35760
rect 0 35368 800 35488
rect 0 34960 800 35080
rect 11200 34824 12000 34944
rect 0 34552 800 34672
rect 0 34144 800 34264
rect 11200 34008 12000 34128
rect 0 33736 800 33856
rect 0 33192 800 33312
rect 11200 33328 12000 33448
rect 0 32784 800 32904
rect 0 32376 800 32496
rect 11200 32512 12000 32632
rect 0 31968 800 32088
rect 0 31560 800 31680
rect 11200 31696 12000 31816
rect 0 31152 800 31272
rect 11200 31016 12000 31136
rect 0 30744 800 30864
rect 0 30336 800 30456
rect 11200 30200 12000 30320
rect 0 29792 800 29912
rect 0 29384 800 29504
rect 11200 29384 12000 29504
rect 0 28976 800 29096
rect 0 28568 800 28688
rect 11200 28704 12000 28824
rect 0 28160 800 28280
rect 0 27752 800 27872
rect 11200 27888 12000 28008
rect 0 27344 800 27464
rect 0 26936 800 27056
rect 11200 27072 12000 27192
rect 0 26392 800 26512
rect 11200 26392 12000 26512
rect 0 25984 800 26104
rect 0 25576 800 25696
rect 11200 25576 12000 25696
rect 0 25168 800 25288
rect 0 24760 800 24880
rect 11200 24760 12000 24880
rect 0 24352 800 24472
rect 0 23944 800 24064
rect 11200 24080 12000 24200
rect 0 23536 800 23656
rect 11200 23264 12000 23384
rect 0 22992 800 23112
rect 0 22584 800 22704
rect 11200 22448 12000 22568
rect 0 22176 800 22296
rect 0 21768 800 21888
rect 11200 21768 12000 21888
rect 0 21360 800 21480
rect 0 20952 800 21072
rect 11200 20952 12000 21072
rect 0 20544 800 20664
rect 0 20136 800 20256
rect 11200 20272 12000 20392
rect 0 19592 800 19712
rect 11200 19456 12000 19576
rect 0 19184 800 19304
rect 0 18776 800 18896
rect 11200 18640 12000 18760
rect 0 18368 800 18488
rect 0 17960 800 18080
rect 11200 17960 12000 18080
rect 0 17552 800 17672
rect 0 17144 800 17264
rect 11200 17144 12000 17264
rect 0 16600 800 16720
rect 0 16192 800 16312
rect 11200 16328 12000 16448
rect 0 15784 800 15904
rect 11200 15648 12000 15768
rect 0 15376 800 15496
rect 0 14968 800 15088
rect 11200 14832 12000 14952
rect 0 14560 800 14680
rect 0 14152 800 14272
rect 11200 14016 12000 14136
rect 0 13744 800 13864
rect 0 13200 800 13320
rect 11200 13336 12000 13456
rect 0 12792 800 12912
rect 0 12384 800 12504
rect 11200 12520 12000 12640
rect 0 11976 800 12096
rect 0 11568 800 11688
rect 11200 11704 12000 11824
rect 0 11160 800 11280
rect 11200 11024 12000 11144
rect 0 10752 800 10872
rect 0 10344 800 10464
rect 11200 10208 12000 10328
rect 0 9800 800 9920
rect 0 9392 800 9512
rect 11200 9392 12000 9512
rect 0 8984 800 9104
rect 0 8576 800 8696
rect 11200 8712 12000 8832
rect 0 8168 800 8288
rect 0 7760 800 7880
rect 11200 7896 12000 8016
rect 0 7352 800 7472
rect 0 6944 800 7064
rect 11200 7080 12000 7200
rect 0 6400 800 6520
rect 11200 6400 12000 6520
rect 0 5992 800 6112
rect 0 5584 800 5704
rect 11200 5584 12000 5704
rect 0 5176 800 5296
rect 0 4768 800 4888
rect 11200 4768 12000 4888
rect 0 4360 800 4480
rect 0 3952 800 4072
rect 11200 4088 12000 4208
rect 0 3544 800 3664
rect 11200 3272 12000 3392
rect 0 3000 800 3120
rect 0 2592 800 2712
rect 11200 2456 12000 2576
rect 0 2184 800 2304
rect 0 1776 800 1896
rect 11200 1776 12000 1896
rect 0 1368 800 1488
rect 0 960 800 1080
rect 11200 960 12000 1080
rect 0 552 800 672
rect 0 144 800 264
rect 11200 280 12000 400
<< obsm3 >>
rect 880 79488 11120 79525
rect 13 79360 11120 79488
rect 880 79352 11120 79360
rect 880 79080 11200 79352
rect 13 78952 11200 79080
rect 880 78816 11200 78952
rect 880 78672 11120 78816
rect 13 78544 11120 78672
rect 880 78536 11120 78544
rect 880 78264 11200 78536
rect 13 78136 11200 78264
rect 880 77856 11120 78136
rect 13 77728 11200 77856
rect 880 77448 11200 77728
rect 13 77320 11200 77448
rect 880 77040 11120 77320
rect 13 76776 11200 77040
rect 880 76504 11200 76776
rect 880 76496 11120 76504
rect 13 76368 11120 76496
rect 880 76224 11120 76368
rect 880 76088 11200 76224
rect 13 75960 11200 76088
rect 880 75824 11200 75960
rect 880 75680 11120 75824
rect 13 75552 11120 75680
rect 880 75544 11120 75552
rect 880 75272 11200 75544
rect 13 75144 11200 75272
rect 880 75008 11200 75144
rect 880 74864 11120 75008
rect 13 74736 11120 74864
rect 880 74728 11120 74736
rect 880 74456 11200 74728
rect 13 74328 11200 74456
rect 880 74192 11200 74328
rect 880 74048 11120 74192
rect 13 73920 11120 74048
rect 880 73912 11120 73920
rect 880 73640 11200 73912
rect 13 73512 11200 73640
rect 13 73376 11120 73512
rect 880 73232 11120 73376
rect 880 73096 11200 73232
rect 13 72968 11200 73096
rect 880 72696 11200 72968
rect 880 72688 11120 72696
rect 13 72560 11120 72688
rect 880 72416 11120 72560
rect 880 72280 11200 72416
rect 13 72152 11200 72280
rect 880 71880 11200 72152
rect 880 71872 11120 71880
rect 13 71744 11120 71872
rect 880 71600 11120 71744
rect 880 71464 11200 71600
rect 13 71336 11200 71464
rect 880 71200 11200 71336
rect 880 71056 11120 71200
rect 13 70928 11120 71056
rect 880 70920 11120 70928
rect 880 70648 11200 70920
rect 13 70520 11200 70648
rect 880 70384 11200 70520
rect 880 70240 11120 70384
rect 13 70104 11120 70240
rect 13 69976 11200 70104
rect 880 69696 11200 69976
rect 13 69568 11200 69696
rect 880 69288 11120 69568
rect 13 69160 11200 69288
rect 880 68888 11200 69160
rect 880 68880 11120 68888
rect 13 68752 11120 68880
rect 880 68608 11120 68752
rect 880 68472 11200 68608
rect 13 68344 11200 68472
rect 880 68072 11200 68344
rect 880 68064 11120 68072
rect 13 67936 11120 68064
rect 880 67792 11120 67936
rect 880 67656 11200 67792
rect 13 67528 11200 67656
rect 880 67256 11200 67528
rect 880 67248 11120 67256
rect 13 67120 11120 67248
rect 880 66976 11120 67120
rect 880 66840 11200 66976
rect 13 66576 11200 66840
rect 880 66296 11120 66576
rect 13 66168 11200 66296
rect 880 65888 11200 66168
rect 13 65760 11200 65888
rect 880 65480 11120 65760
rect 13 65352 11200 65480
rect 880 65072 11200 65352
rect 13 64944 11200 65072
rect 880 64664 11120 64944
rect 13 64536 11200 64664
rect 880 64264 11200 64536
rect 880 64256 11120 64264
rect 13 64128 11120 64256
rect 880 63984 11120 64128
rect 880 63848 11200 63984
rect 13 63720 11200 63848
rect 880 63448 11200 63720
rect 880 63440 11120 63448
rect 13 63176 11120 63440
rect 880 63168 11120 63176
rect 880 62896 11200 63168
rect 13 62768 11200 62896
rect 880 62632 11200 62768
rect 880 62488 11120 62632
rect 13 62360 11120 62488
rect 880 62352 11120 62360
rect 880 62080 11200 62352
rect 13 61952 11200 62080
rect 880 61672 11120 61952
rect 13 61544 11200 61672
rect 880 61264 11200 61544
rect 13 61136 11200 61264
rect 880 60856 11120 61136
rect 13 60728 11200 60856
rect 880 60456 11200 60728
rect 880 60448 11120 60456
rect 13 60320 11120 60448
rect 880 60176 11120 60320
rect 880 60040 11200 60176
rect 13 59776 11200 60040
rect 880 59640 11200 59776
rect 880 59496 11120 59640
rect 13 59368 11120 59496
rect 880 59360 11120 59368
rect 880 59088 11200 59360
rect 13 58960 11200 59088
rect 880 58824 11200 58960
rect 880 58680 11120 58824
rect 13 58552 11120 58680
rect 880 58544 11120 58552
rect 880 58272 11200 58544
rect 13 58144 11200 58272
rect 880 57864 11120 58144
rect 13 57736 11200 57864
rect 880 57456 11200 57736
rect 13 57328 11200 57456
rect 880 57048 11120 57328
rect 13 56784 11200 57048
rect 880 56512 11200 56784
rect 880 56504 11120 56512
rect 13 56376 11120 56504
rect 880 56232 11120 56376
rect 880 56096 11200 56232
rect 13 55968 11200 56096
rect 880 55832 11200 55968
rect 880 55688 11120 55832
rect 13 55560 11120 55688
rect 880 55552 11120 55560
rect 880 55280 11200 55552
rect 13 55152 11200 55280
rect 880 55016 11200 55152
rect 880 54872 11120 55016
rect 13 54744 11120 54872
rect 880 54736 11120 54744
rect 880 54464 11200 54736
rect 13 54336 11200 54464
rect 880 54200 11200 54336
rect 880 54056 11120 54200
rect 13 53928 11120 54056
rect 880 53920 11120 53928
rect 880 53648 11200 53920
rect 13 53520 11200 53648
rect 13 53384 11120 53520
rect 880 53240 11120 53384
rect 880 53104 11200 53240
rect 13 52976 11200 53104
rect 880 52704 11200 52976
rect 880 52696 11120 52704
rect 13 52568 11120 52696
rect 880 52424 11120 52568
rect 880 52288 11200 52424
rect 13 52160 11200 52288
rect 880 51888 11200 52160
rect 880 51880 11120 51888
rect 13 51752 11120 51880
rect 880 51608 11120 51752
rect 880 51472 11200 51608
rect 13 51344 11200 51472
rect 880 51208 11200 51344
rect 880 51064 11120 51208
rect 13 50936 11120 51064
rect 880 50928 11120 50936
rect 880 50656 11200 50928
rect 13 50528 11200 50656
rect 880 50392 11200 50528
rect 880 50248 11120 50392
rect 13 50112 11120 50248
rect 13 49984 11200 50112
rect 880 49704 11200 49984
rect 13 49576 11200 49704
rect 880 49296 11120 49576
rect 13 49168 11200 49296
rect 880 48896 11200 49168
rect 880 48888 11120 48896
rect 13 48760 11120 48888
rect 880 48616 11120 48760
rect 880 48480 11200 48616
rect 13 48352 11200 48480
rect 880 48080 11200 48352
rect 880 48072 11120 48080
rect 13 47944 11120 48072
rect 880 47800 11120 47944
rect 880 47664 11200 47800
rect 13 47536 11200 47664
rect 880 47264 11200 47536
rect 880 47256 11120 47264
rect 13 47128 11120 47256
rect 880 46984 11120 47128
rect 880 46848 11200 46984
rect 13 46584 11200 46848
rect 880 46304 11120 46584
rect 13 46176 11200 46304
rect 880 45896 11200 46176
rect 13 45768 11200 45896
rect 880 45488 11120 45768
rect 13 45360 11200 45488
rect 880 45080 11200 45360
rect 13 44952 11200 45080
rect 880 44672 11120 44952
rect 13 44544 11200 44672
rect 880 44272 11200 44544
rect 880 44264 11120 44272
rect 13 44136 11120 44264
rect 880 43992 11120 44136
rect 880 43856 11200 43992
rect 13 43728 11200 43856
rect 880 43456 11200 43728
rect 880 43448 11120 43456
rect 13 43184 11120 43448
rect 880 43176 11120 43184
rect 880 42904 11200 43176
rect 13 42776 11200 42904
rect 880 42640 11200 42776
rect 880 42496 11120 42640
rect 13 42368 11120 42496
rect 880 42360 11120 42368
rect 880 42088 11200 42360
rect 13 41960 11200 42088
rect 880 41680 11120 41960
rect 13 41552 11200 41680
rect 880 41272 11200 41552
rect 13 41144 11200 41272
rect 880 40864 11120 41144
rect 13 40736 11200 40864
rect 880 40464 11200 40736
rect 880 40456 11120 40464
rect 13 40328 11120 40456
rect 880 40184 11120 40328
rect 880 40048 11200 40184
rect 13 39784 11200 40048
rect 880 39648 11200 39784
rect 880 39504 11120 39648
rect 13 39376 11120 39504
rect 880 39368 11120 39376
rect 880 39096 11200 39368
rect 13 38968 11200 39096
rect 880 38832 11200 38968
rect 880 38688 11120 38832
rect 13 38560 11120 38688
rect 880 38552 11120 38560
rect 880 38280 11200 38552
rect 13 38152 11200 38280
rect 880 37872 11120 38152
rect 13 37744 11200 37872
rect 880 37464 11200 37744
rect 13 37336 11200 37464
rect 880 37056 11120 37336
rect 13 36792 11200 37056
rect 880 36520 11200 36792
rect 880 36512 11120 36520
rect 13 36384 11120 36512
rect 880 36240 11120 36384
rect 880 36104 11200 36240
rect 13 35976 11200 36104
rect 880 35840 11200 35976
rect 880 35696 11120 35840
rect 13 35568 11120 35696
rect 880 35560 11120 35568
rect 880 35288 11200 35560
rect 13 35160 11200 35288
rect 880 35024 11200 35160
rect 880 34880 11120 35024
rect 13 34752 11120 34880
rect 880 34744 11120 34752
rect 880 34472 11200 34744
rect 13 34344 11200 34472
rect 880 34208 11200 34344
rect 880 34064 11120 34208
rect 13 33936 11120 34064
rect 880 33928 11120 33936
rect 880 33656 11200 33928
rect 13 33528 11200 33656
rect 13 33392 11120 33528
rect 880 33248 11120 33392
rect 880 33112 11200 33248
rect 13 32984 11200 33112
rect 880 32712 11200 32984
rect 880 32704 11120 32712
rect 13 32576 11120 32704
rect 880 32432 11120 32576
rect 880 32296 11200 32432
rect 13 32168 11200 32296
rect 880 31896 11200 32168
rect 880 31888 11120 31896
rect 13 31760 11120 31888
rect 880 31616 11120 31760
rect 880 31480 11200 31616
rect 13 31352 11200 31480
rect 880 31216 11200 31352
rect 880 31072 11120 31216
rect 13 30944 11120 31072
rect 880 30936 11120 30944
rect 880 30664 11200 30936
rect 13 30536 11200 30664
rect 880 30400 11200 30536
rect 880 30256 11120 30400
rect 13 30120 11120 30256
rect 13 29992 11200 30120
rect 880 29712 11200 29992
rect 13 29584 11200 29712
rect 880 29304 11120 29584
rect 13 29176 11200 29304
rect 880 28904 11200 29176
rect 880 28896 11120 28904
rect 13 28768 11120 28896
rect 880 28624 11120 28768
rect 880 28488 11200 28624
rect 13 28360 11200 28488
rect 880 28088 11200 28360
rect 880 28080 11120 28088
rect 13 27952 11120 28080
rect 880 27808 11120 27952
rect 880 27672 11200 27808
rect 13 27544 11200 27672
rect 880 27272 11200 27544
rect 880 27264 11120 27272
rect 13 27136 11120 27264
rect 880 26992 11120 27136
rect 880 26856 11200 26992
rect 13 26592 11200 26856
rect 880 26312 11120 26592
rect 13 26184 11200 26312
rect 880 25904 11200 26184
rect 13 25776 11200 25904
rect 880 25496 11120 25776
rect 13 25368 11200 25496
rect 880 25088 11200 25368
rect 13 24960 11200 25088
rect 880 24680 11120 24960
rect 13 24552 11200 24680
rect 880 24280 11200 24552
rect 880 24272 11120 24280
rect 13 24144 11120 24272
rect 880 24000 11120 24144
rect 880 23864 11200 24000
rect 13 23736 11200 23864
rect 880 23464 11200 23736
rect 880 23456 11120 23464
rect 13 23192 11120 23456
rect 880 23184 11120 23192
rect 880 22912 11200 23184
rect 13 22784 11200 22912
rect 880 22648 11200 22784
rect 880 22504 11120 22648
rect 13 22376 11120 22504
rect 880 22368 11120 22376
rect 880 22096 11200 22368
rect 13 21968 11200 22096
rect 880 21688 11120 21968
rect 13 21560 11200 21688
rect 880 21280 11200 21560
rect 13 21152 11200 21280
rect 880 20872 11120 21152
rect 13 20744 11200 20872
rect 880 20472 11200 20744
rect 880 20464 11120 20472
rect 13 20336 11120 20464
rect 880 20192 11120 20336
rect 880 20056 11200 20192
rect 13 19792 11200 20056
rect 880 19656 11200 19792
rect 880 19512 11120 19656
rect 13 19384 11120 19512
rect 880 19376 11120 19384
rect 880 19104 11200 19376
rect 13 18976 11200 19104
rect 880 18840 11200 18976
rect 880 18696 11120 18840
rect 13 18568 11120 18696
rect 880 18560 11120 18568
rect 880 18288 11200 18560
rect 13 18160 11200 18288
rect 880 17880 11120 18160
rect 13 17752 11200 17880
rect 880 17472 11200 17752
rect 13 17344 11200 17472
rect 880 17064 11120 17344
rect 13 16800 11200 17064
rect 880 16528 11200 16800
rect 880 16520 11120 16528
rect 13 16392 11120 16520
rect 880 16248 11120 16392
rect 880 16112 11200 16248
rect 13 15984 11200 16112
rect 880 15848 11200 15984
rect 880 15704 11120 15848
rect 13 15576 11120 15704
rect 880 15568 11120 15576
rect 880 15296 11200 15568
rect 13 15168 11200 15296
rect 880 15032 11200 15168
rect 880 14888 11120 15032
rect 13 14760 11120 14888
rect 880 14752 11120 14760
rect 880 14480 11200 14752
rect 13 14352 11200 14480
rect 880 14216 11200 14352
rect 880 14072 11120 14216
rect 13 13944 11120 14072
rect 880 13936 11120 13944
rect 880 13664 11200 13936
rect 13 13536 11200 13664
rect 13 13400 11120 13536
rect 880 13256 11120 13400
rect 880 13120 11200 13256
rect 13 12992 11200 13120
rect 880 12720 11200 12992
rect 880 12712 11120 12720
rect 13 12584 11120 12712
rect 880 12440 11120 12584
rect 880 12304 11200 12440
rect 13 12176 11200 12304
rect 880 11904 11200 12176
rect 880 11896 11120 11904
rect 13 11768 11120 11896
rect 880 11624 11120 11768
rect 880 11488 11200 11624
rect 13 11360 11200 11488
rect 880 11224 11200 11360
rect 880 11080 11120 11224
rect 13 10952 11120 11080
rect 880 10944 11120 10952
rect 880 10672 11200 10944
rect 13 10544 11200 10672
rect 880 10408 11200 10544
rect 880 10264 11120 10408
rect 13 10128 11120 10264
rect 13 10000 11200 10128
rect 880 9720 11200 10000
rect 13 9592 11200 9720
rect 880 9312 11120 9592
rect 13 9184 11200 9312
rect 880 8912 11200 9184
rect 880 8904 11120 8912
rect 13 8776 11120 8904
rect 880 8632 11120 8776
rect 880 8496 11200 8632
rect 13 8368 11200 8496
rect 880 8096 11200 8368
rect 880 8088 11120 8096
rect 13 7960 11120 8088
rect 880 7816 11120 7960
rect 880 7680 11200 7816
rect 13 7552 11200 7680
rect 880 7280 11200 7552
rect 880 7272 11120 7280
rect 13 7144 11120 7272
rect 880 7000 11120 7144
rect 880 6864 11200 7000
rect 13 6600 11200 6864
rect 880 6320 11120 6600
rect 13 6192 11200 6320
rect 880 5912 11200 6192
rect 13 5784 11200 5912
rect 880 5504 11120 5784
rect 13 5376 11200 5504
rect 880 5096 11200 5376
rect 13 4968 11200 5096
rect 880 4688 11120 4968
rect 13 4560 11200 4688
rect 880 4288 11200 4560
rect 880 4280 11120 4288
rect 13 4152 11120 4280
rect 880 4008 11120 4152
rect 880 3872 11200 4008
rect 13 3744 11200 3872
rect 880 3472 11200 3744
rect 880 3464 11120 3472
rect 13 3200 11120 3464
rect 880 3192 11120 3200
rect 880 2920 11200 3192
rect 13 2792 11200 2920
rect 880 2656 11200 2792
rect 880 2512 11120 2656
rect 13 2384 11120 2512
rect 880 2376 11120 2384
rect 880 2104 11200 2376
rect 13 1976 11200 2104
rect 880 1696 11120 1976
rect 13 1568 11200 1696
rect 880 1288 11200 1568
rect 13 1160 11200 1288
rect 880 880 11120 1160
rect 13 752 11200 880
rect 880 480 11200 752
rect 880 472 11120 480
rect 13 344 11120 472
rect 880 200 11120 344
rect 880 171 11200 200
<< metal4 >>
rect 2576 2128 2896 77840
rect 4208 2128 4528 77840
rect 5840 2128 6160 77840
rect 7472 2128 7792 77840
rect 9104 2128 9424 77840
<< obsm4 >>
rect 243 5203 2496 74765
rect 2976 5203 4128 74765
rect 4608 5203 5760 74765
rect 6240 5203 6381 74765
<< labels >>
rlabel metal4 s 2576 2128 2896 77840 6 vccd1
port 1 nsew power input
rlabel metal4 s 5840 2128 6160 77840 6 vccd1
port 1 nsew power input
rlabel metal4 s 9104 2128 9424 77840 6 vccd1
port 1 nsew power input
rlabel metal4 s 4208 2128 4528 77840 6 vssd1
port 2 nsew ground input
rlabel metal4 s 7472 2128 7792 77840 6 vssd1
port 2 nsew ground input
rlabel metal3 s 0 79568 800 79688 6 wb_clk_i
port 3 nsew signal input
rlabel metal2 s 5998 79200 6054 80000 6 wb_rst_i
port 4 nsew signal input
rlabel metal3 s 11200 79432 12000 79552 6 wbm_a_ack_i
port 5 nsew signal input
rlabel metal3 s 11200 5584 12000 5704 6 wbm_a_adr_o[0]
port 6 nsew signal output
rlabel metal3 s 11200 13336 12000 13456 6 wbm_a_adr_o[10]
port 7 nsew signal output
rlabel metal3 s 11200 14016 12000 14136 6 wbm_a_adr_o[11]
port 8 nsew signal output
rlabel metal3 s 11200 14832 12000 14952 6 wbm_a_adr_o[12]
port 9 nsew signal output
rlabel metal3 s 11200 15648 12000 15768 6 wbm_a_adr_o[13]
port 10 nsew signal output
rlabel metal3 s 11200 16328 12000 16448 6 wbm_a_adr_o[14]
port 11 nsew signal output
rlabel metal3 s 11200 17144 12000 17264 6 wbm_a_adr_o[15]
port 12 nsew signal output
rlabel metal3 s 11200 17960 12000 18080 6 wbm_a_adr_o[16]
port 13 nsew signal output
rlabel metal3 s 11200 18640 12000 18760 6 wbm_a_adr_o[17]
port 14 nsew signal output
rlabel metal3 s 11200 19456 12000 19576 6 wbm_a_adr_o[18]
port 15 nsew signal output
rlabel metal3 s 11200 20272 12000 20392 6 wbm_a_adr_o[19]
port 16 nsew signal output
rlabel metal3 s 11200 6400 12000 6520 6 wbm_a_adr_o[1]
port 17 nsew signal output
rlabel metal3 s 11200 20952 12000 21072 6 wbm_a_adr_o[20]
port 18 nsew signal output
rlabel metal3 s 11200 21768 12000 21888 6 wbm_a_adr_o[21]
port 19 nsew signal output
rlabel metal3 s 11200 22448 12000 22568 6 wbm_a_adr_o[22]
port 20 nsew signal output
rlabel metal3 s 11200 23264 12000 23384 6 wbm_a_adr_o[23]
port 21 nsew signal output
rlabel metal3 s 11200 24080 12000 24200 6 wbm_a_adr_o[24]
port 22 nsew signal output
rlabel metal3 s 11200 24760 12000 24880 6 wbm_a_adr_o[25]
port 23 nsew signal output
rlabel metal3 s 11200 25576 12000 25696 6 wbm_a_adr_o[26]
port 24 nsew signal output
rlabel metal3 s 11200 26392 12000 26512 6 wbm_a_adr_o[27]
port 25 nsew signal output
rlabel metal3 s 11200 27072 12000 27192 6 wbm_a_adr_o[28]
port 26 nsew signal output
rlabel metal3 s 11200 27888 12000 28008 6 wbm_a_adr_o[29]
port 27 nsew signal output
rlabel metal3 s 11200 7080 12000 7200 6 wbm_a_adr_o[2]
port 28 nsew signal output
rlabel metal3 s 11200 28704 12000 28824 6 wbm_a_adr_o[30]
port 29 nsew signal output
rlabel metal3 s 11200 29384 12000 29504 6 wbm_a_adr_o[31]
port 30 nsew signal output
rlabel metal3 s 11200 7896 12000 8016 6 wbm_a_adr_o[3]
port 31 nsew signal output
rlabel metal3 s 11200 8712 12000 8832 6 wbm_a_adr_o[4]
port 32 nsew signal output
rlabel metal3 s 11200 9392 12000 9512 6 wbm_a_adr_o[5]
port 33 nsew signal output
rlabel metal3 s 11200 10208 12000 10328 6 wbm_a_adr_o[6]
port 34 nsew signal output
rlabel metal3 s 11200 11024 12000 11144 6 wbm_a_adr_o[7]
port 35 nsew signal output
rlabel metal3 s 11200 11704 12000 11824 6 wbm_a_adr_o[8]
port 36 nsew signal output
rlabel metal3 s 11200 12520 12000 12640 6 wbm_a_adr_o[9]
port 37 nsew signal output
rlabel metal3 s 11200 960 12000 1080 6 wbm_a_cyc_o
port 38 nsew signal output
rlabel metal3 s 11200 54816 12000 54936 6 wbm_a_dat_i[0]
port 39 nsew signal input
rlabel metal3 s 11200 62432 12000 62552 6 wbm_a_dat_i[10]
port 40 nsew signal input
rlabel metal3 s 11200 63248 12000 63368 6 wbm_a_dat_i[11]
port 41 nsew signal input
rlabel metal3 s 11200 64064 12000 64184 6 wbm_a_dat_i[12]
port 42 nsew signal input
rlabel metal3 s 11200 64744 12000 64864 6 wbm_a_dat_i[13]
port 43 nsew signal input
rlabel metal3 s 11200 65560 12000 65680 6 wbm_a_dat_i[14]
port 44 nsew signal input
rlabel metal3 s 11200 66376 12000 66496 6 wbm_a_dat_i[15]
port 45 nsew signal input
rlabel metal3 s 11200 67056 12000 67176 6 wbm_a_dat_i[16]
port 46 nsew signal input
rlabel metal3 s 11200 67872 12000 67992 6 wbm_a_dat_i[17]
port 47 nsew signal input
rlabel metal3 s 11200 68688 12000 68808 6 wbm_a_dat_i[18]
port 48 nsew signal input
rlabel metal3 s 11200 69368 12000 69488 6 wbm_a_dat_i[19]
port 49 nsew signal input
rlabel metal3 s 11200 55632 12000 55752 6 wbm_a_dat_i[1]
port 50 nsew signal input
rlabel metal3 s 11200 70184 12000 70304 6 wbm_a_dat_i[20]
port 51 nsew signal input
rlabel metal3 s 11200 71000 12000 71120 6 wbm_a_dat_i[21]
port 52 nsew signal input
rlabel metal3 s 11200 71680 12000 71800 6 wbm_a_dat_i[22]
port 53 nsew signal input
rlabel metal3 s 11200 72496 12000 72616 6 wbm_a_dat_i[23]
port 54 nsew signal input
rlabel metal3 s 11200 73312 12000 73432 6 wbm_a_dat_i[24]
port 55 nsew signal input
rlabel metal3 s 11200 73992 12000 74112 6 wbm_a_dat_i[25]
port 56 nsew signal input
rlabel metal3 s 11200 74808 12000 74928 6 wbm_a_dat_i[26]
port 57 nsew signal input
rlabel metal3 s 11200 75624 12000 75744 6 wbm_a_dat_i[27]
port 58 nsew signal input
rlabel metal3 s 11200 76304 12000 76424 6 wbm_a_dat_i[28]
port 59 nsew signal input
rlabel metal3 s 11200 77120 12000 77240 6 wbm_a_dat_i[29]
port 60 nsew signal input
rlabel metal3 s 11200 56312 12000 56432 6 wbm_a_dat_i[2]
port 61 nsew signal input
rlabel metal3 s 11200 77936 12000 78056 6 wbm_a_dat_i[30]
port 62 nsew signal input
rlabel metal3 s 11200 78616 12000 78736 6 wbm_a_dat_i[31]
port 63 nsew signal input
rlabel metal3 s 11200 57128 12000 57248 6 wbm_a_dat_i[3]
port 64 nsew signal input
rlabel metal3 s 11200 57944 12000 58064 6 wbm_a_dat_i[4]
port 65 nsew signal input
rlabel metal3 s 11200 58624 12000 58744 6 wbm_a_dat_i[5]
port 66 nsew signal input
rlabel metal3 s 11200 59440 12000 59560 6 wbm_a_dat_i[6]
port 67 nsew signal input
rlabel metal3 s 11200 60256 12000 60376 6 wbm_a_dat_i[7]
port 68 nsew signal input
rlabel metal3 s 11200 60936 12000 61056 6 wbm_a_dat_i[8]
port 69 nsew signal input
rlabel metal3 s 11200 61752 12000 61872 6 wbm_a_dat_i[9]
port 70 nsew signal input
rlabel metal3 s 11200 30200 12000 30320 6 wbm_a_dat_o[0]
port 71 nsew signal output
rlabel metal3 s 11200 37952 12000 38072 6 wbm_a_dat_o[10]
port 72 nsew signal output
rlabel metal3 s 11200 38632 12000 38752 6 wbm_a_dat_o[11]
port 73 nsew signal output
rlabel metal3 s 11200 39448 12000 39568 6 wbm_a_dat_o[12]
port 74 nsew signal output
rlabel metal3 s 11200 40264 12000 40384 6 wbm_a_dat_o[13]
port 75 nsew signal output
rlabel metal3 s 11200 40944 12000 41064 6 wbm_a_dat_o[14]
port 76 nsew signal output
rlabel metal3 s 11200 41760 12000 41880 6 wbm_a_dat_o[15]
port 77 nsew signal output
rlabel metal3 s 11200 42440 12000 42560 6 wbm_a_dat_o[16]
port 78 nsew signal output
rlabel metal3 s 11200 43256 12000 43376 6 wbm_a_dat_o[17]
port 79 nsew signal output
rlabel metal3 s 11200 44072 12000 44192 6 wbm_a_dat_o[18]
port 80 nsew signal output
rlabel metal3 s 11200 44752 12000 44872 6 wbm_a_dat_o[19]
port 81 nsew signal output
rlabel metal3 s 11200 31016 12000 31136 6 wbm_a_dat_o[1]
port 82 nsew signal output
rlabel metal3 s 11200 45568 12000 45688 6 wbm_a_dat_o[20]
port 83 nsew signal output
rlabel metal3 s 11200 46384 12000 46504 6 wbm_a_dat_o[21]
port 84 nsew signal output
rlabel metal3 s 11200 47064 12000 47184 6 wbm_a_dat_o[22]
port 85 nsew signal output
rlabel metal3 s 11200 47880 12000 48000 6 wbm_a_dat_o[23]
port 86 nsew signal output
rlabel metal3 s 11200 48696 12000 48816 6 wbm_a_dat_o[24]
port 87 nsew signal output
rlabel metal3 s 11200 49376 12000 49496 6 wbm_a_dat_o[25]
port 88 nsew signal output
rlabel metal3 s 11200 50192 12000 50312 6 wbm_a_dat_o[26]
port 89 nsew signal output
rlabel metal3 s 11200 51008 12000 51128 6 wbm_a_dat_o[27]
port 90 nsew signal output
rlabel metal3 s 11200 51688 12000 51808 6 wbm_a_dat_o[28]
port 91 nsew signal output
rlabel metal3 s 11200 52504 12000 52624 6 wbm_a_dat_o[29]
port 92 nsew signal output
rlabel metal3 s 11200 31696 12000 31816 6 wbm_a_dat_o[2]
port 93 nsew signal output
rlabel metal3 s 11200 53320 12000 53440 6 wbm_a_dat_o[30]
port 94 nsew signal output
rlabel metal3 s 11200 54000 12000 54120 6 wbm_a_dat_o[31]
port 95 nsew signal output
rlabel metal3 s 11200 32512 12000 32632 6 wbm_a_dat_o[3]
port 96 nsew signal output
rlabel metal3 s 11200 33328 12000 33448 6 wbm_a_dat_o[4]
port 97 nsew signal output
rlabel metal3 s 11200 34008 12000 34128 6 wbm_a_dat_o[5]
port 98 nsew signal output
rlabel metal3 s 11200 34824 12000 34944 6 wbm_a_dat_o[6]
port 99 nsew signal output
rlabel metal3 s 11200 35640 12000 35760 6 wbm_a_dat_o[7]
port 100 nsew signal output
rlabel metal3 s 11200 36320 12000 36440 6 wbm_a_dat_o[8]
port 101 nsew signal output
rlabel metal3 s 11200 37136 12000 37256 6 wbm_a_dat_o[9]
port 102 nsew signal output
rlabel metal3 s 11200 2456 12000 2576 6 wbm_a_sel_o[0]
port 103 nsew signal output
rlabel metal3 s 11200 3272 12000 3392 6 wbm_a_sel_o[1]
port 104 nsew signal output
rlabel metal3 s 11200 4088 12000 4208 6 wbm_a_sel_o[2]
port 105 nsew signal output
rlabel metal3 s 11200 4768 12000 4888 6 wbm_a_sel_o[3]
port 106 nsew signal output
rlabel metal3 s 11200 280 12000 400 6 wbm_a_stb_o
port 107 nsew signal output
rlabel metal3 s 11200 1776 12000 1896 6 wbm_a_we_o
port 108 nsew signal output
rlabel metal3 s 0 79160 800 79280 6 wbm_b_ack_i
port 109 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 wbm_b_adr_o[0]
port 110 nsew signal output
rlabel metal3 s 0 51552 800 51672 6 wbm_b_adr_o[10]
port 111 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 wbm_b_adr_o[1]
port 112 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 wbm_b_adr_o[2]
port 113 nsew signal output
rlabel metal3 s 0 48560 800 48680 6 wbm_b_adr_o[3]
port 114 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 wbm_b_adr_o[4]
port 115 nsew signal output
rlabel metal3 s 0 49376 800 49496 6 wbm_b_adr_o[5]
port 116 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 wbm_b_adr_o[6]
port 117 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 wbm_b_adr_o[7]
port 118 nsew signal output
rlabel metal3 s 0 50736 800 50856 6 wbm_b_adr_o[8]
port 119 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 wbm_b_adr_o[9]
port 120 nsew signal output
rlabel metal3 s 0 44752 800 44872 6 wbm_b_cyc_o
port 121 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 wbm_b_dat_i[0]
port 122 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 wbm_b_dat_i[10]
port 123 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 wbm_b_dat_i[11]
port 124 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 wbm_b_dat_i[12]
port 125 nsew signal input
rlabel metal3 s 0 71136 800 71256 6 wbm_b_dat_i[13]
port 126 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 wbm_b_dat_i[14]
port 127 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 wbm_b_dat_i[15]
port 128 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 wbm_b_dat_i[16]
port 129 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 wbm_b_dat_i[17]
port 130 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 wbm_b_dat_i[18]
port 131 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 wbm_b_dat_i[19]
port 132 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 wbm_b_dat_i[1]
port 133 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 wbm_b_dat_i[20]
port 134 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 wbm_b_dat_i[21]
port 135 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 wbm_b_dat_i[22]
port 136 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 wbm_b_dat_i[23]
port 137 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 wbm_b_dat_i[24]
port 138 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 wbm_b_dat_i[25]
port 139 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 wbm_b_dat_i[26]
port 140 nsew signal input
rlabel metal3 s 0 77120 800 77240 6 wbm_b_dat_i[27]
port 141 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 wbm_b_dat_i[28]
port 142 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 wbm_b_dat_i[29]
port 143 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 wbm_b_dat_i[2]
port 144 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 wbm_b_dat_i[30]
port 145 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 wbm_b_dat_i[31]
port 146 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 wbm_b_dat_i[3]
port 147 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 wbm_b_dat_i[4]
port 148 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 wbm_b_dat_i[5]
port 149 nsew signal input
rlabel metal3 s 0 68144 800 68264 6 wbm_b_dat_i[6]
port 150 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 wbm_b_dat_i[7]
port 151 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 wbm_b_dat_i[8]
port 152 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 wbm_b_dat_i[9]
port 153 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 wbm_b_dat_o[0]
port 154 nsew signal output
rlabel metal3 s 0 56176 800 56296 6 wbm_b_dat_o[10]
port 155 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 wbm_b_dat_o[11]
port 156 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 wbm_b_dat_o[12]
port 157 nsew signal output
rlabel metal3 s 0 57536 800 57656 6 wbm_b_dat_o[13]
port 158 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 wbm_b_dat_o[14]
port 159 nsew signal output
rlabel metal3 s 0 58352 800 58472 6 wbm_b_dat_o[15]
port 160 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 wbm_b_dat_o[16]
port 161 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 wbm_b_dat_o[17]
port 162 nsew signal output
rlabel metal3 s 0 59576 800 59696 6 wbm_b_dat_o[18]
port 163 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 wbm_b_dat_o[19]
port 164 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 wbm_b_dat_o[1]
port 165 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 wbm_b_dat_o[20]
port 166 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 wbm_b_dat_o[21]
port 167 nsew signal output
rlabel metal3 s 0 61344 800 61464 6 wbm_b_dat_o[22]
port 168 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 wbm_b_dat_o[23]
port 169 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 wbm_b_dat_o[24]
port 170 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 wbm_b_dat_o[25]
port 171 nsew signal output
rlabel metal3 s 0 62976 800 63096 6 wbm_b_dat_o[26]
port 172 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 wbm_b_dat_o[27]
port 173 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 wbm_b_dat_o[28]
port 174 nsew signal output
rlabel metal3 s 0 64336 800 64456 6 wbm_b_dat_o[29]
port 175 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 wbm_b_dat_o[2]
port 176 nsew signal output
rlabel metal3 s 0 64744 800 64864 6 wbm_b_dat_o[30]
port 177 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 wbm_b_dat_o[31]
port 178 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 wbm_b_dat_o[3]
port 179 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 wbm_b_dat_o[4]
port 180 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 wbm_b_dat_o[5]
port 181 nsew signal output
rlabel metal3 s 0 54544 800 54664 6 wbm_b_dat_o[6]
port 182 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 wbm_b_dat_o[7]
port 183 nsew signal output
rlabel metal3 s 0 55360 800 55480 6 wbm_b_dat_o[8]
port 184 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 wbm_b_dat_o[9]
port 185 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 wbm_b_sel_o[0]
port 186 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 wbm_b_sel_o[1]
port 187 nsew signal output
rlabel metal3 s 0 46384 800 46504 6 wbm_b_sel_o[2]
port 188 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 wbm_b_sel_o[3]
port 189 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 wbm_b_stb_o
port 190 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 wbm_b_we_o
port 191 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 wbs_ack_o
port 192 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 wbs_adr_i[0]
port 193 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 wbs_adr_i[10]
port 194 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 wbs_adr_i[11]
port 195 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 wbs_adr_i[12]
port 196 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 wbs_adr_i[13]
port 197 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 wbs_adr_i[14]
port 198 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 wbs_adr_i[15]
port 199 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 wbs_adr_i[16]
port 200 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 wbs_adr_i[17]
port 201 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 wbs_adr_i[18]
port 202 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 wbs_adr_i[19]
port 203 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 wbs_adr_i[1]
port 204 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_adr_i[20]
port 205 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 wbs_adr_i[21]
port 206 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 wbs_adr_i[22]
port 207 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 wbs_adr_i[23]
port 208 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 wbs_adr_i[24]
port 209 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 wbs_adr_i[25]
port 210 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 wbs_adr_i[26]
port 211 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 wbs_adr_i[27]
port 212 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 wbs_adr_i[28]
port 213 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 wbs_adr_i[29]
port 214 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 wbs_adr_i[2]
port 215 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 wbs_adr_i[30]
port 216 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 wbs_adr_i[31]
port 217 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 wbs_adr_i[3]
port 218 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 wbs_adr_i[4]
port 219 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 wbs_adr_i[5]
port 220 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 wbs_adr_i[6]
port 221 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 wbs_adr_i[7]
port 222 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 wbs_adr_i[8]
port 223 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 wbs_adr_i[9]
port 224 nsew signal input
rlabel metal3 s 0 552 800 672 6 wbs_cyc_i
port 225 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 wbs_dat_i[0]
port 226 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 wbs_dat_i[10]
port 227 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 wbs_dat_i[11]
port 228 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 wbs_dat_i[12]
port 229 nsew signal input
rlabel metal3 s 0 22176 800 22296 6 wbs_dat_i[13]
port 230 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 wbs_dat_i[14]
port 231 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 wbs_dat_i[15]
port 232 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 wbs_dat_i[16]
port 233 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 wbs_dat_i[17]
port 234 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 wbs_dat_i[18]
port 235 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 wbs_dat_i[19]
port 236 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 wbs_dat_i[1]
port 237 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 wbs_dat_i[20]
port 238 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 wbs_dat_i[21]
port 239 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 wbs_dat_i[22]
port 240 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 wbs_dat_i[23]
port 241 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 wbs_dat_i[24]
port 242 nsew signal input
rlabel metal3 s 0 27344 800 27464 6 wbs_dat_i[25]
port 243 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 wbs_dat_i[26]
port 244 nsew signal input
rlabel metal3 s 0 28160 800 28280 6 wbs_dat_i[27]
port 245 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 wbs_dat_i[28]
port 246 nsew signal input
rlabel metal3 s 0 28976 800 29096 6 wbs_dat_i[29]
port 247 nsew signal input
rlabel metal3 s 0 17552 800 17672 6 wbs_dat_i[2]
port 248 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 wbs_dat_i[30]
port 249 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 wbs_dat_i[31]
port 250 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 wbs_dat_i[3]
port 251 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 wbs_dat_i[4]
port 252 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 wbs_dat_i[5]
port 253 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 wbs_dat_i[6]
port 254 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 wbs_dat_i[7]
port 255 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 wbs_dat_i[8]
port 256 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 wbs_dat_i[9]
port 257 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 wbs_dat_o[0]
port 258 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 wbs_dat_o[10]
port 259 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 wbs_dat_o[11]
port 260 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_o[12]
port 261 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 wbs_dat_o[13]
port 262 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 wbs_dat_o[14]
port 263 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 wbs_dat_o[15]
port 264 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 wbs_dat_o[16]
port 265 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 wbs_dat_o[17]
port 266 nsew signal output
rlabel metal3 s 0 37952 800 38072 6 wbs_dat_o[18]
port 267 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 wbs_dat_o[19]
port 268 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 wbs_dat_o[1]
port 269 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 wbs_dat_o[20]
port 270 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 wbs_dat_o[21]
port 271 nsew signal output
rlabel metal3 s 0 39584 800 39704 6 wbs_dat_o[22]
port 272 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 wbs_dat_o[23]
port 273 nsew signal output
rlabel metal3 s 0 40536 800 40656 6 wbs_dat_o[24]
port 274 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 wbs_dat_o[25]
port 275 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 wbs_dat_o[26]
port 276 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 wbs_dat_o[27]
port 277 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 wbs_dat_o[28]
port 278 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 wbs_dat_o[29]
port 279 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 wbs_dat_o[2]
port 280 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 wbs_dat_o[30]
port 281 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 wbs_dat_o[31]
port 282 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 wbs_dat_o[3]
port 283 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 wbs_dat_o[4]
port 284 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 wbs_dat_o[5]
port 285 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 wbs_dat_o[6]
port 286 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 wbs_dat_o[7]
port 287 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 wbs_dat_o[8]
port 288 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 wbs_dat_o[9]
port 289 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 wbs_sel_i[0]
port 290 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 wbs_sel_i[1]
port 291 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wbs_sel_i[2]
port 292 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 wbs_sel_i[3]
port 293 nsew signal input
rlabel metal3 s 0 144 800 264 6 wbs_stb_i
port 294 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wbs_we_i
port 295 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1837948
string GDS_FILE /openlane/designs/wb_bridge/runs/RUN_2022.03.17_23.03.05/results/finishing/wb_bridge_2way.magic.gds
string GDS_START 131198
<< end >>

