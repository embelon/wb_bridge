VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_bridge_2way
  CLASS BLOCK ;
  FOREIGN wb_bridge_2way ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 400.000 ;
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 12.880 10.640 14.480 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.200 10.640 30.800 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.520 10.640 47.120 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.360 10.640 38.960 389.200 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 396.000 30.270 400.000 ;
    END
  END wb_rst_i
  PIN wbm_a_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 397.160 60.000 397.760 ;
    END
  END wbm_a_ack_i
  PIN wbm_a_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 27.920 60.000 28.520 ;
    END
  END wbm_a_adr_o[0]
  PIN wbm_a_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 66.680 60.000 67.280 ;
    END
  END wbm_a_adr_o[10]
  PIN wbm_a_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 70.080 60.000 70.680 ;
    END
  END wbm_a_adr_o[11]
  PIN wbm_a_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 74.160 60.000 74.760 ;
    END
  END wbm_a_adr_o[12]
  PIN wbm_a_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 78.240 60.000 78.840 ;
    END
  END wbm_a_adr_o[13]
  PIN wbm_a_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 81.640 60.000 82.240 ;
    END
  END wbm_a_adr_o[14]
  PIN wbm_a_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 85.720 60.000 86.320 ;
    END
  END wbm_a_adr_o[15]
  PIN wbm_a_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 89.800 60.000 90.400 ;
    END
  END wbm_a_adr_o[16]
  PIN wbm_a_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 93.200 60.000 93.800 ;
    END
  END wbm_a_adr_o[17]
  PIN wbm_a_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 97.280 60.000 97.880 ;
    END
  END wbm_a_adr_o[18]
  PIN wbm_a_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 101.360 60.000 101.960 ;
    END
  END wbm_a_adr_o[19]
  PIN wbm_a_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 32.000 60.000 32.600 ;
    END
  END wbm_a_adr_o[1]
  PIN wbm_a_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 104.760 60.000 105.360 ;
    END
  END wbm_a_adr_o[20]
  PIN wbm_a_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 108.840 60.000 109.440 ;
    END
  END wbm_a_adr_o[21]
  PIN wbm_a_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 112.240 60.000 112.840 ;
    END
  END wbm_a_adr_o[22]
  PIN wbm_a_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 116.320 60.000 116.920 ;
    END
  END wbm_a_adr_o[23]
  PIN wbm_a_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 120.400 60.000 121.000 ;
    END
  END wbm_a_adr_o[24]
  PIN wbm_a_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 123.800 60.000 124.400 ;
    END
  END wbm_a_adr_o[25]
  PIN wbm_a_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 127.880 60.000 128.480 ;
    END
  END wbm_a_adr_o[26]
  PIN wbm_a_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 131.960 60.000 132.560 ;
    END
  END wbm_a_adr_o[27]
  PIN wbm_a_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 135.360 60.000 135.960 ;
    END
  END wbm_a_adr_o[28]
  PIN wbm_a_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 139.440 60.000 140.040 ;
    END
  END wbm_a_adr_o[29]
  PIN wbm_a_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 35.400 60.000 36.000 ;
    END
  END wbm_a_adr_o[2]
  PIN wbm_a_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 143.520 60.000 144.120 ;
    END
  END wbm_a_adr_o[30]
  PIN wbm_a_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 146.920 60.000 147.520 ;
    END
  END wbm_a_adr_o[31]
  PIN wbm_a_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 39.480 60.000 40.080 ;
    END
  END wbm_a_adr_o[3]
  PIN wbm_a_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 43.560 60.000 44.160 ;
    END
  END wbm_a_adr_o[4]
  PIN wbm_a_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 46.960 60.000 47.560 ;
    END
  END wbm_a_adr_o[5]
  PIN wbm_a_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 51.040 60.000 51.640 ;
    END
  END wbm_a_adr_o[6]
  PIN wbm_a_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 55.120 60.000 55.720 ;
    END
  END wbm_a_adr_o[7]
  PIN wbm_a_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 58.520 60.000 59.120 ;
    END
  END wbm_a_adr_o[8]
  PIN wbm_a_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 62.600 60.000 63.200 ;
    END
  END wbm_a_adr_o[9]
  PIN wbm_a_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 4.800 60.000 5.400 ;
    END
  END wbm_a_cyc_o
  PIN wbm_a_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 274.080 60.000 274.680 ;
    END
  END wbm_a_dat_i[0]
  PIN wbm_a_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 312.160 60.000 312.760 ;
    END
  END wbm_a_dat_i[10]
  PIN wbm_a_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 316.240 60.000 316.840 ;
    END
  END wbm_a_dat_i[11]
  PIN wbm_a_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 320.320 60.000 320.920 ;
    END
  END wbm_a_dat_i[12]
  PIN wbm_a_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 323.720 60.000 324.320 ;
    END
  END wbm_a_dat_i[13]
  PIN wbm_a_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 327.800 60.000 328.400 ;
    END
  END wbm_a_dat_i[14]
  PIN wbm_a_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 331.880 60.000 332.480 ;
    END
  END wbm_a_dat_i[15]
  PIN wbm_a_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 335.280 60.000 335.880 ;
    END
  END wbm_a_dat_i[16]
  PIN wbm_a_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 339.360 60.000 339.960 ;
    END
  END wbm_a_dat_i[17]
  PIN wbm_a_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 343.440 60.000 344.040 ;
    END
  END wbm_a_dat_i[18]
  PIN wbm_a_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 346.840 60.000 347.440 ;
    END
  END wbm_a_dat_i[19]
  PIN wbm_a_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 278.160 60.000 278.760 ;
    END
  END wbm_a_dat_i[1]
  PIN wbm_a_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 350.920 60.000 351.520 ;
    END
  END wbm_a_dat_i[20]
  PIN wbm_a_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 355.000 60.000 355.600 ;
    END
  END wbm_a_dat_i[21]
  PIN wbm_a_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 358.400 60.000 359.000 ;
    END
  END wbm_a_dat_i[22]
  PIN wbm_a_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 362.480 60.000 363.080 ;
    END
  END wbm_a_dat_i[23]
  PIN wbm_a_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 366.560 60.000 367.160 ;
    END
  END wbm_a_dat_i[24]
  PIN wbm_a_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 369.960 60.000 370.560 ;
    END
  END wbm_a_dat_i[25]
  PIN wbm_a_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 374.040 60.000 374.640 ;
    END
  END wbm_a_dat_i[26]
  PIN wbm_a_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 378.120 60.000 378.720 ;
    END
  END wbm_a_dat_i[27]
  PIN wbm_a_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 381.520 60.000 382.120 ;
    END
  END wbm_a_dat_i[28]
  PIN wbm_a_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 385.600 60.000 386.200 ;
    END
  END wbm_a_dat_i[29]
  PIN wbm_a_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 281.560 60.000 282.160 ;
    END
  END wbm_a_dat_i[2]
  PIN wbm_a_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 389.680 60.000 390.280 ;
    END
  END wbm_a_dat_i[30]
  PIN wbm_a_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 393.080 60.000 393.680 ;
    END
  END wbm_a_dat_i[31]
  PIN wbm_a_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 285.640 60.000 286.240 ;
    END
  END wbm_a_dat_i[3]
  PIN wbm_a_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 289.720 60.000 290.320 ;
    END
  END wbm_a_dat_i[4]
  PIN wbm_a_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 293.120 60.000 293.720 ;
    END
  END wbm_a_dat_i[5]
  PIN wbm_a_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 297.200 60.000 297.800 ;
    END
  END wbm_a_dat_i[6]
  PIN wbm_a_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 301.280 60.000 301.880 ;
    END
  END wbm_a_dat_i[7]
  PIN wbm_a_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 304.680 60.000 305.280 ;
    END
  END wbm_a_dat_i[8]
  PIN wbm_a_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 308.760 60.000 309.360 ;
    END
  END wbm_a_dat_i[9]
  PIN wbm_a_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 151.000 60.000 151.600 ;
    END
  END wbm_a_dat_o[0]
  PIN wbm_a_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 189.760 60.000 190.360 ;
    END
  END wbm_a_dat_o[10]
  PIN wbm_a_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 193.160 60.000 193.760 ;
    END
  END wbm_a_dat_o[11]
  PIN wbm_a_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 197.240 60.000 197.840 ;
    END
  END wbm_a_dat_o[12]
  PIN wbm_a_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 201.320 60.000 201.920 ;
    END
  END wbm_a_dat_o[13]
  PIN wbm_a_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 204.720 60.000 205.320 ;
    END
  END wbm_a_dat_o[14]
  PIN wbm_a_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 208.800 60.000 209.400 ;
    END
  END wbm_a_dat_o[15]
  PIN wbm_a_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 212.200 60.000 212.800 ;
    END
  END wbm_a_dat_o[16]
  PIN wbm_a_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 216.280 60.000 216.880 ;
    END
  END wbm_a_dat_o[17]
  PIN wbm_a_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 220.360 60.000 220.960 ;
    END
  END wbm_a_dat_o[18]
  PIN wbm_a_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 223.760 60.000 224.360 ;
    END
  END wbm_a_dat_o[19]
  PIN wbm_a_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 155.080 60.000 155.680 ;
    END
  END wbm_a_dat_o[1]
  PIN wbm_a_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 227.840 60.000 228.440 ;
    END
  END wbm_a_dat_o[20]
  PIN wbm_a_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 231.920 60.000 232.520 ;
    END
  END wbm_a_dat_o[21]
  PIN wbm_a_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 235.320 60.000 235.920 ;
    END
  END wbm_a_dat_o[22]
  PIN wbm_a_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 239.400 60.000 240.000 ;
    END
  END wbm_a_dat_o[23]
  PIN wbm_a_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 243.480 60.000 244.080 ;
    END
  END wbm_a_dat_o[24]
  PIN wbm_a_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 246.880 60.000 247.480 ;
    END
  END wbm_a_dat_o[25]
  PIN wbm_a_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 250.960 60.000 251.560 ;
    END
  END wbm_a_dat_o[26]
  PIN wbm_a_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 255.040 60.000 255.640 ;
    END
  END wbm_a_dat_o[27]
  PIN wbm_a_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 258.440 60.000 259.040 ;
    END
  END wbm_a_dat_o[28]
  PIN wbm_a_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 262.520 60.000 263.120 ;
    END
  END wbm_a_dat_o[29]
  PIN wbm_a_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 158.480 60.000 159.080 ;
    END
  END wbm_a_dat_o[2]
  PIN wbm_a_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 266.600 60.000 267.200 ;
    END
  END wbm_a_dat_o[30]
  PIN wbm_a_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 270.000 60.000 270.600 ;
    END
  END wbm_a_dat_o[31]
  PIN wbm_a_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 162.560 60.000 163.160 ;
    END
  END wbm_a_dat_o[3]
  PIN wbm_a_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 166.640 60.000 167.240 ;
    END
  END wbm_a_dat_o[4]
  PIN wbm_a_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 170.040 60.000 170.640 ;
    END
  END wbm_a_dat_o[5]
  PIN wbm_a_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 174.120 60.000 174.720 ;
    END
  END wbm_a_dat_o[6]
  PIN wbm_a_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 178.200 60.000 178.800 ;
    END
  END wbm_a_dat_o[7]
  PIN wbm_a_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 181.600 60.000 182.200 ;
    END
  END wbm_a_dat_o[8]
  PIN wbm_a_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 185.680 60.000 186.280 ;
    END
  END wbm_a_dat_o[9]
  PIN wbm_a_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 12.280 60.000 12.880 ;
    END
  END wbm_a_sel_o[0]
  PIN wbm_a_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 16.360 60.000 16.960 ;
    END
  END wbm_a_sel_o[1]
  PIN wbm_a_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 20.440 60.000 21.040 ;
    END
  END wbm_a_sel_o[2]
  PIN wbm_a_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 23.840 60.000 24.440 ;
    END
  END wbm_a_sel_o[3]
  PIN wbm_a_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 1.400 60.000 2.000 ;
    END
  END wbm_a_stb_o
  PIN wbm_a_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 8.880 60.000 9.480 ;
    END
  END wbm_a_we_o
  PIN wbm_b_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END wbm_b_ack_i
  PIN wbm_b_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END wbm_b_adr_o[0]
  PIN wbm_b_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END wbm_b_adr_o[10]
  PIN wbm_b_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END wbm_b_adr_o[1]
  PIN wbm_b_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END wbm_b_adr_o[2]
  PIN wbm_b_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END wbm_b_adr_o[3]
  PIN wbm_b_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END wbm_b_adr_o[4]
  PIN wbm_b_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END wbm_b_adr_o[5]
  PIN wbm_b_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END wbm_b_adr_o[6]
  PIN wbm_b_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END wbm_b_adr_o[7]
  PIN wbm_b_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END wbm_b_adr_o[8]
  PIN wbm_b_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END wbm_b_adr_o[9]
  PIN wbm_b_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END wbm_b_cyc_o
  PIN wbm_b_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END wbm_b_dat_i[0]
  PIN wbm_b_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END wbm_b_dat_i[10]
  PIN wbm_b_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END wbm_b_dat_i[11]
  PIN wbm_b_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END wbm_b_dat_i[12]
  PIN wbm_b_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END wbm_b_dat_i[13]
  PIN wbm_b_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END wbm_b_dat_i[14]
  PIN wbm_b_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END wbm_b_dat_i[15]
  PIN wbm_b_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END wbm_b_dat_i[16]
  PIN wbm_b_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END wbm_b_dat_i[17]
  PIN wbm_b_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END wbm_b_dat_i[18]
  PIN wbm_b_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END wbm_b_dat_i[19]
  PIN wbm_b_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END wbm_b_dat_i[1]
  PIN wbm_b_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END wbm_b_dat_i[20]
  PIN wbm_b_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END wbm_b_dat_i[21]
  PIN wbm_b_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END wbm_b_dat_i[22]
  PIN wbm_b_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END wbm_b_dat_i[23]
  PIN wbm_b_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END wbm_b_dat_i[24]
  PIN wbm_b_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END wbm_b_dat_i[25]
  PIN wbm_b_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END wbm_b_dat_i[26]
  PIN wbm_b_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END wbm_b_dat_i[27]
  PIN wbm_b_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END wbm_b_dat_i[28]
  PIN wbm_b_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END wbm_b_dat_i[29]
  PIN wbm_b_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END wbm_b_dat_i[2]
  PIN wbm_b_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END wbm_b_dat_i[30]
  PIN wbm_b_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END wbm_b_dat_i[31]
  PIN wbm_b_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END wbm_b_dat_i[3]
  PIN wbm_b_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END wbm_b_dat_i[4]
  PIN wbm_b_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END wbm_b_dat_i[5]
  PIN wbm_b_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END wbm_b_dat_i[6]
  PIN wbm_b_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END wbm_b_dat_i[7]
  PIN wbm_b_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END wbm_b_dat_i[8]
  PIN wbm_b_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END wbm_b_dat_i[9]
  PIN wbm_b_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END wbm_b_dat_o[0]
  PIN wbm_b_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END wbm_b_dat_o[10]
  PIN wbm_b_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END wbm_b_dat_o[11]
  PIN wbm_b_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END wbm_b_dat_o[12]
  PIN wbm_b_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END wbm_b_dat_o[13]
  PIN wbm_b_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END wbm_b_dat_o[14]
  PIN wbm_b_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END wbm_b_dat_o[15]
  PIN wbm_b_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END wbm_b_dat_o[16]
  PIN wbm_b_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END wbm_b_dat_o[17]
  PIN wbm_b_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END wbm_b_dat_o[18]
  PIN wbm_b_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END wbm_b_dat_o[19]
  PIN wbm_b_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END wbm_b_dat_o[1]
  PIN wbm_b_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END wbm_b_dat_o[20]
  PIN wbm_b_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END wbm_b_dat_o[21]
  PIN wbm_b_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END wbm_b_dat_o[22]
  PIN wbm_b_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END wbm_b_dat_o[23]
  PIN wbm_b_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END wbm_b_dat_o[24]
  PIN wbm_b_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END wbm_b_dat_o[25]
  PIN wbm_b_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END wbm_b_dat_o[26]
  PIN wbm_b_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.960 4.000 319.560 ;
    END
  END wbm_b_dat_o[27]
  PIN wbm_b_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END wbm_b_dat_o[28]
  PIN wbm_b_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END wbm_b_dat_o[29]
  PIN wbm_b_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END wbm_b_dat_o[2]
  PIN wbm_b_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END wbm_b_dat_o[30]
  PIN wbm_b_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END wbm_b_dat_o[31]
  PIN wbm_b_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END wbm_b_dat_o[3]
  PIN wbm_b_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END wbm_b_dat_o[4]
  PIN wbm_b_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END wbm_b_dat_o[5]
  PIN wbm_b_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END wbm_b_dat_o[6]
  PIN wbm_b_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END wbm_b_dat_o[7]
  PIN wbm_b_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END wbm_b_dat_o[8]
  PIN wbm_b_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END wbm_b_dat_o[9]
  PIN wbm_b_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END wbm_b_sel_o[0]
  PIN wbm_b_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END wbm_b_sel_o[1]
  PIN wbm_b_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END wbm_b_sel_o[2]
  PIN wbm_b_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END wbm_b_sel_o[3]
  PIN wbm_b_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END wbm_b_stb_o
  PIN wbm_b_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END wbm_b_we_o
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 54.280 389.045 ;
      LAYER met1 ;
        RECT 0.070 5.140 54.280 389.200 ;
      LAYER met2 ;
        RECT 0.100 395.720 29.710 398.325 ;
        RECT 30.550 395.720 51.420 398.325 ;
        RECT 0.100 4.280 51.420 395.720 ;
        RECT 0.100 0.835 29.710 4.280 ;
        RECT 30.550 0.835 51.420 4.280 ;
      LAYER met3 ;
        RECT 4.400 398.160 56.000 398.305 ;
        RECT 4.400 397.440 55.600 398.160 ;
        RECT 0.270 396.800 55.600 397.440 ;
        RECT 4.400 396.760 55.600 396.800 ;
        RECT 4.400 395.400 56.000 396.760 ;
        RECT 0.270 394.760 56.000 395.400 ;
        RECT 4.400 394.080 56.000 394.760 ;
        RECT 4.400 393.360 55.600 394.080 ;
        RECT 0.270 392.720 55.600 393.360 ;
        RECT 4.400 392.680 55.600 392.720 ;
        RECT 4.400 391.320 56.000 392.680 ;
        RECT 0.270 390.680 56.000 391.320 ;
        RECT 4.400 389.280 55.600 390.680 ;
        RECT 0.270 388.640 56.000 389.280 ;
        RECT 4.400 387.240 56.000 388.640 ;
        RECT 0.270 386.600 56.000 387.240 ;
        RECT 0.270 385.920 55.600 386.600 ;
        RECT 4.400 385.200 55.600 385.920 ;
        RECT 4.400 384.520 56.000 385.200 ;
        RECT 0.270 383.880 56.000 384.520 ;
        RECT 4.400 382.520 56.000 383.880 ;
        RECT 4.400 382.480 55.600 382.520 ;
        RECT 0.270 381.840 55.600 382.480 ;
        RECT 4.400 381.120 55.600 381.840 ;
        RECT 4.400 380.440 56.000 381.120 ;
        RECT 0.270 379.800 56.000 380.440 ;
        RECT 4.400 379.120 56.000 379.800 ;
        RECT 4.400 378.400 55.600 379.120 ;
        RECT 0.270 377.760 55.600 378.400 ;
        RECT 4.400 377.720 55.600 377.760 ;
        RECT 4.400 376.360 56.000 377.720 ;
        RECT 0.270 375.720 56.000 376.360 ;
        RECT 4.400 375.040 56.000 375.720 ;
        RECT 4.400 374.320 55.600 375.040 ;
        RECT 0.270 373.680 55.600 374.320 ;
        RECT 4.400 373.640 55.600 373.680 ;
        RECT 4.400 372.280 56.000 373.640 ;
        RECT 0.270 370.960 56.000 372.280 ;
        RECT 4.400 369.560 55.600 370.960 ;
        RECT 0.270 368.920 56.000 369.560 ;
        RECT 4.400 367.560 56.000 368.920 ;
        RECT 4.400 367.520 55.600 367.560 ;
        RECT 0.270 366.880 55.600 367.520 ;
        RECT 4.400 366.160 55.600 366.880 ;
        RECT 4.400 365.480 56.000 366.160 ;
        RECT 0.270 364.840 56.000 365.480 ;
        RECT 4.400 363.480 56.000 364.840 ;
        RECT 4.400 363.440 55.600 363.480 ;
        RECT 0.270 362.800 55.600 363.440 ;
        RECT 4.400 362.080 55.600 362.800 ;
        RECT 4.400 361.400 56.000 362.080 ;
        RECT 0.270 360.760 56.000 361.400 ;
        RECT 4.400 359.400 56.000 360.760 ;
        RECT 4.400 359.360 55.600 359.400 ;
        RECT 0.270 358.720 55.600 359.360 ;
        RECT 4.400 358.000 55.600 358.720 ;
        RECT 4.400 357.320 56.000 358.000 ;
        RECT 0.270 356.000 56.000 357.320 ;
        RECT 4.400 354.600 55.600 356.000 ;
        RECT 0.270 353.960 56.000 354.600 ;
        RECT 4.400 352.560 56.000 353.960 ;
        RECT 0.270 351.920 56.000 352.560 ;
        RECT 4.400 350.520 55.600 351.920 ;
        RECT 0.270 349.880 56.000 350.520 ;
        RECT 4.400 348.480 56.000 349.880 ;
        RECT 0.270 347.840 56.000 348.480 ;
        RECT 4.400 346.440 55.600 347.840 ;
        RECT 0.270 345.800 56.000 346.440 ;
        RECT 4.400 344.440 56.000 345.800 ;
        RECT 4.400 344.400 55.600 344.440 ;
        RECT 0.270 343.760 55.600 344.400 ;
        RECT 4.400 343.040 55.600 343.760 ;
        RECT 4.400 342.360 56.000 343.040 ;
        RECT 0.270 341.040 56.000 342.360 ;
        RECT 4.400 340.360 56.000 341.040 ;
        RECT 4.400 339.640 55.600 340.360 ;
        RECT 0.270 339.000 55.600 339.640 ;
        RECT 4.400 338.960 55.600 339.000 ;
        RECT 4.400 337.600 56.000 338.960 ;
        RECT 0.270 336.960 56.000 337.600 ;
        RECT 4.400 336.280 56.000 336.960 ;
        RECT 4.400 335.560 55.600 336.280 ;
        RECT 0.270 334.920 55.600 335.560 ;
        RECT 4.400 334.880 55.600 334.920 ;
        RECT 4.400 333.520 56.000 334.880 ;
        RECT 0.270 332.880 56.000 333.520 ;
        RECT 4.400 331.480 55.600 332.880 ;
        RECT 0.270 330.840 56.000 331.480 ;
        RECT 4.400 329.440 56.000 330.840 ;
        RECT 0.270 328.800 56.000 329.440 ;
        RECT 4.400 327.400 55.600 328.800 ;
        RECT 0.270 326.080 56.000 327.400 ;
        RECT 4.400 324.720 56.000 326.080 ;
        RECT 4.400 324.680 55.600 324.720 ;
        RECT 0.270 324.040 55.600 324.680 ;
        RECT 4.400 323.320 55.600 324.040 ;
        RECT 4.400 322.640 56.000 323.320 ;
        RECT 0.270 322.000 56.000 322.640 ;
        RECT 4.400 321.320 56.000 322.000 ;
        RECT 4.400 320.600 55.600 321.320 ;
        RECT 0.270 319.960 55.600 320.600 ;
        RECT 4.400 319.920 55.600 319.960 ;
        RECT 4.400 318.560 56.000 319.920 ;
        RECT 0.270 317.920 56.000 318.560 ;
        RECT 4.400 317.240 56.000 317.920 ;
        RECT 4.400 316.520 55.600 317.240 ;
        RECT 0.270 315.880 55.600 316.520 ;
        RECT 4.400 315.840 55.600 315.880 ;
        RECT 4.400 314.480 56.000 315.840 ;
        RECT 0.270 313.840 56.000 314.480 ;
        RECT 4.400 313.160 56.000 313.840 ;
        RECT 4.400 312.440 55.600 313.160 ;
        RECT 0.270 311.760 55.600 312.440 ;
        RECT 0.270 311.120 56.000 311.760 ;
        RECT 4.400 309.760 56.000 311.120 ;
        RECT 4.400 309.720 55.600 309.760 ;
        RECT 0.270 309.080 55.600 309.720 ;
        RECT 4.400 308.360 55.600 309.080 ;
        RECT 4.400 307.680 56.000 308.360 ;
        RECT 0.270 307.040 56.000 307.680 ;
        RECT 4.400 305.680 56.000 307.040 ;
        RECT 4.400 305.640 55.600 305.680 ;
        RECT 0.270 305.000 55.600 305.640 ;
        RECT 4.400 304.280 55.600 305.000 ;
        RECT 4.400 303.600 56.000 304.280 ;
        RECT 0.270 302.960 56.000 303.600 ;
        RECT 4.400 302.280 56.000 302.960 ;
        RECT 4.400 301.560 55.600 302.280 ;
        RECT 0.270 300.920 55.600 301.560 ;
        RECT 4.400 300.880 55.600 300.920 ;
        RECT 4.400 299.520 56.000 300.880 ;
        RECT 0.270 298.880 56.000 299.520 ;
        RECT 4.400 298.200 56.000 298.880 ;
        RECT 4.400 297.480 55.600 298.200 ;
        RECT 0.270 296.800 55.600 297.480 ;
        RECT 0.270 296.160 56.000 296.800 ;
        RECT 4.400 294.760 56.000 296.160 ;
        RECT 0.270 294.120 56.000 294.760 ;
        RECT 4.400 292.720 55.600 294.120 ;
        RECT 0.270 292.080 56.000 292.720 ;
        RECT 4.400 290.720 56.000 292.080 ;
        RECT 4.400 290.680 55.600 290.720 ;
        RECT 0.270 290.040 55.600 290.680 ;
        RECT 4.400 289.320 55.600 290.040 ;
        RECT 4.400 288.640 56.000 289.320 ;
        RECT 0.270 288.000 56.000 288.640 ;
        RECT 4.400 286.640 56.000 288.000 ;
        RECT 4.400 286.600 55.600 286.640 ;
        RECT 0.270 285.960 55.600 286.600 ;
        RECT 4.400 285.240 55.600 285.960 ;
        RECT 4.400 284.560 56.000 285.240 ;
        RECT 0.270 283.920 56.000 284.560 ;
        RECT 4.400 282.560 56.000 283.920 ;
        RECT 4.400 282.520 55.600 282.560 ;
        RECT 0.270 281.200 55.600 282.520 ;
        RECT 4.400 281.160 55.600 281.200 ;
        RECT 4.400 279.800 56.000 281.160 ;
        RECT 0.270 279.160 56.000 279.800 ;
        RECT 4.400 277.760 55.600 279.160 ;
        RECT 0.270 277.120 56.000 277.760 ;
        RECT 4.400 275.720 56.000 277.120 ;
        RECT 0.270 275.080 56.000 275.720 ;
        RECT 4.400 273.680 55.600 275.080 ;
        RECT 0.270 273.040 56.000 273.680 ;
        RECT 4.400 271.640 56.000 273.040 ;
        RECT 0.270 271.000 56.000 271.640 ;
        RECT 4.400 269.600 55.600 271.000 ;
        RECT 0.270 268.960 56.000 269.600 ;
        RECT 4.400 267.600 56.000 268.960 ;
        RECT 4.400 267.560 55.600 267.600 ;
        RECT 0.270 266.240 55.600 267.560 ;
        RECT 4.400 266.200 55.600 266.240 ;
        RECT 4.400 264.840 56.000 266.200 ;
        RECT 0.270 264.200 56.000 264.840 ;
        RECT 4.400 263.520 56.000 264.200 ;
        RECT 4.400 262.800 55.600 263.520 ;
        RECT 0.270 262.160 55.600 262.800 ;
        RECT 4.400 262.120 55.600 262.160 ;
        RECT 4.400 260.760 56.000 262.120 ;
        RECT 0.270 260.120 56.000 260.760 ;
        RECT 4.400 259.440 56.000 260.120 ;
        RECT 4.400 258.720 55.600 259.440 ;
        RECT 0.270 258.080 55.600 258.720 ;
        RECT 4.400 258.040 55.600 258.080 ;
        RECT 4.400 256.680 56.000 258.040 ;
        RECT 0.270 256.040 56.000 256.680 ;
        RECT 4.400 254.640 55.600 256.040 ;
        RECT 0.270 254.000 56.000 254.640 ;
        RECT 4.400 252.600 56.000 254.000 ;
        RECT 0.270 251.960 56.000 252.600 ;
        RECT 0.270 251.280 55.600 251.960 ;
        RECT 4.400 250.560 55.600 251.280 ;
        RECT 4.400 249.880 56.000 250.560 ;
        RECT 0.270 249.240 56.000 249.880 ;
        RECT 4.400 247.880 56.000 249.240 ;
        RECT 4.400 247.840 55.600 247.880 ;
        RECT 0.270 247.200 55.600 247.840 ;
        RECT 4.400 246.480 55.600 247.200 ;
        RECT 4.400 245.800 56.000 246.480 ;
        RECT 0.270 245.160 56.000 245.800 ;
        RECT 4.400 244.480 56.000 245.160 ;
        RECT 4.400 243.760 55.600 244.480 ;
        RECT 0.270 243.120 55.600 243.760 ;
        RECT 4.400 243.080 55.600 243.120 ;
        RECT 4.400 241.720 56.000 243.080 ;
        RECT 0.270 241.080 56.000 241.720 ;
        RECT 4.400 240.400 56.000 241.080 ;
        RECT 4.400 239.680 55.600 240.400 ;
        RECT 0.270 239.040 55.600 239.680 ;
        RECT 4.400 239.000 55.600 239.040 ;
        RECT 4.400 237.640 56.000 239.000 ;
        RECT 0.270 236.320 56.000 237.640 ;
        RECT 4.400 234.920 55.600 236.320 ;
        RECT 0.270 234.280 56.000 234.920 ;
        RECT 4.400 232.920 56.000 234.280 ;
        RECT 4.400 232.880 55.600 232.920 ;
        RECT 0.270 232.240 55.600 232.880 ;
        RECT 4.400 231.520 55.600 232.240 ;
        RECT 4.400 230.840 56.000 231.520 ;
        RECT 0.270 230.200 56.000 230.840 ;
        RECT 4.400 228.840 56.000 230.200 ;
        RECT 4.400 228.800 55.600 228.840 ;
        RECT 0.270 228.160 55.600 228.800 ;
        RECT 4.400 227.440 55.600 228.160 ;
        RECT 4.400 226.760 56.000 227.440 ;
        RECT 0.270 226.120 56.000 226.760 ;
        RECT 4.400 224.760 56.000 226.120 ;
        RECT 4.400 224.720 55.600 224.760 ;
        RECT 0.270 224.080 55.600 224.720 ;
        RECT 4.400 223.360 55.600 224.080 ;
        RECT 4.400 222.680 56.000 223.360 ;
        RECT 0.270 221.360 56.000 222.680 ;
        RECT 4.400 219.960 55.600 221.360 ;
        RECT 0.270 219.320 56.000 219.960 ;
        RECT 4.400 217.920 56.000 219.320 ;
        RECT 0.270 217.280 56.000 217.920 ;
        RECT 4.400 215.880 55.600 217.280 ;
        RECT 0.270 215.240 56.000 215.880 ;
        RECT 4.400 213.840 56.000 215.240 ;
        RECT 0.270 213.200 56.000 213.840 ;
        RECT 4.400 211.800 55.600 213.200 ;
        RECT 0.270 211.160 56.000 211.800 ;
        RECT 4.400 209.800 56.000 211.160 ;
        RECT 4.400 209.760 55.600 209.800 ;
        RECT 0.270 209.120 55.600 209.760 ;
        RECT 4.400 208.400 55.600 209.120 ;
        RECT 4.400 207.720 56.000 208.400 ;
        RECT 0.270 206.400 56.000 207.720 ;
        RECT 4.400 205.720 56.000 206.400 ;
        RECT 4.400 205.000 55.600 205.720 ;
        RECT 0.270 204.360 55.600 205.000 ;
        RECT 4.400 204.320 55.600 204.360 ;
        RECT 4.400 202.960 56.000 204.320 ;
        RECT 0.270 202.320 56.000 202.960 ;
        RECT 4.400 200.920 55.600 202.320 ;
        RECT 0.270 200.280 56.000 200.920 ;
        RECT 4.400 198.880 56.000 200.280 ;
        RECT 0.270 198.240 56.000 198.880 ;
        RECT 4.400 196.840 55.600 198.240 ;
        RECT 0.270 196.200 56.000 196.840 ;
        RECT 4.400 194.800 56.000 196.200 ;
        RECT 0.270 194.160 56.000 194.800 ;
        RECT 0.270 193.480 55.600 194.160 ;
        RECT 4.400 192.760 55.600 193.480 ;
        RECT 4.400 192.080 56.000 192.760 ;
        RECT 0.270 191.440 56.000 192.080 ;
        RECT 4.400 190.760 56.000 191.440 ;
        RECT 4.400 190.040 55.600 190.760 ;
        RECT 0.270 189.400 55.600 190.040 ;
        RECT 4.400 189.360 55.600 189.400 ;
        RECT 4.400 188.000 56.000 189.360 ;
        RECT 0.270 187.360 56.000 188.000 ;
        RECT 4.400 186.680 56.000 187.360 ;
        RECT 4.400 185.960 55.600 186.680 ;
        RECT 0.270 185.320 55.600 185.960 ;
        RECT 4.400 185.280 55.600 185.320 ;
        RECT 4.400 183.920 56.000 185.280 ;
        RECT 0.270 183.280 56.000 183.920 ;
        RECT 4.400 182.600 56.000 183.280 ;
        RECT 4.400 181.880 55.600 182.600 ;
        RECT 0.270 181.240 55.600 181.880 ;
        RECT 4.400 181.200 55.600 181.240 ;
        RECT 4.400 179.840 56.000 181.200 ;
        RECT 0.270 179.200 56.000 179.840 ;
        RECT 0.270 178.520 55.600 179.200 ;
        RECT 4.400 177.800 55.600 178.520 ;
        RECT 4.400 177.120 56.000 177.800 ;
        RECT 0.270 176.480 56.000 177.120 ;
        RECT 4.400 175.120 56.000 176.480 ;
        RECT 4.400 175.080 55.600 175.120 ;
        RECT 0.270 174.440 55.600 175.080 ;
        RECT 4.400 173.720 55.600 174.440 ;
        RECT 4.400 173.040 56.000 173.720 ;
        RECT 0.270 172.400 56.000 173.040 ;
        RECT 4.400 171.040 56.000 172.400 ;
        RECT 4.400 171.000 55.600 171.040 ;
        RECT 0.270 170.360 55.600 171.000 ;
        RECT 4.400 169.640 55.600 170.360 ;
        RECT 4.400 168.960 56.000 169.640 ;
        RECT 0.270 168.320 56.000 168.960 ;
        RECT 4.400 167.640 56.000 168.320 ;
        RECT 4.400 166.920 55.600 167.640 ;
        RECT 0.270 166.280 55.600 166.920 ;
        RECT 4.400 166.240 55.600 166.280 ;
        RECT 4.400 164.880 56.000 166.240 ;
        RECT 0.270 163.560 56.000 164.880 ;
        RECT 4.400 162.160 55.600 163.560 ;
        RECT 0.270 161.520 56.000 162.160 ;
        RECT 4.400 160.120 56.000 161.520 ;
        RECT 0.270 159.480 56.000 160.120 ;
        RECT 4.400 158.080 55.600 159.480 ;
        RECT 0.270 157.440 56.000 158.080 ;
        RECT 4.400 156.080 56.000 157.440 ;
        RECT 4.400 156.040 55.600 156.080 ;
        RECT 0.270 155.400 55.600 156.040 ;
        RECT 4.400 154.680 55.600 155.400 ;
        RECT 4.400 154.000 56.000 154.680 ;
        RECT 0.270 153.360 56.000 154.000 ;
        RECT 4.400 152.000 56.000 153.360 ;
        RECT 4.400 151.960 55.600 152.000 ;
        RECT 0.270 151.320 55.600 151.960 ;
        RECT 4.400 150.600 55.600 151.320 ;
        RECT 4.400 149.920 56.000 150.600 ;
        RECT 0.270 148.600 56.000 149.920 ;
        RECT 4.400 147.920 56.000 148.600 ;
        RECT 4.400 147.200 55.600 147.920 ;
        RECT 0.270 146.560 55.600 147.200 ;
        RECT 4.400 146.520 55.600 146.560 ;
        RECT 4.400 145.160 56.000 146.520 ;
        RECT 0.270 144.520 56.000 145.160 ;
        RECT 4.400 143.120 55.600 144.520 ;
        RECT 0.270 142.480 56.000 143.120 ;
        RECT 4.400 141.080 56.000 142.480 ;
        RECT 0.270 140.440 56.000 141.080 ;
        RECT 4.400 139.040 55.600 140.440 ;
        RECT 0.270 138.400 56.000 139.040 ;
        RECT 4.400 137.000 56.000 138.400 ;
        RECT 0.270 136.360 56.000 137.000 ;
        RECT 4.400 134.960 55.600 136.360 ;
        RECT 0.270 133.640 56.000 134.960 ;
        RECT 4.400 132.960 56.000 133.640 ;
        RECT 4.400 132.240 55.600 132.960 ;
        RECT 0.270 131.600 55.600 132.240 ;
        RECT 4.400 131.560 55.600 131.600 ;
        RECT 4.400 130.200 56.000 131.560 ;
        RECT 0.270 129.560 56.000 130.200 ;
        RECT 4.400 128.880 56.000 129.560 ;
        RECT 4.400 128.160 55.600 128.880 ;
        RECT 0.270 127.520 55.600 128.160 ;
        RECT 4.400 127.480 55.600 127.520 ;
        RECT 4.400 126.120 56.000 127.480 ;
        RECT 0.270 125.480 56.000 126.120 ;
        RECT 4.400 124.800 56.000 125.480 ;
        RECT 4.400 124.080 55.600 124.800 ;
        RECT 0.270 123.440 55.600 124.080 ;
        RECT 4.400 123.400 55.600 123.440 ;
        RECT 4.400 122.040 56.000 123.400 ;
        RECT 0.270 121.400 56.000 122.040 ;
        RECT 4.400 120.000 55.600 121.400 ;
        RECT 0.270 118.680 56.000 120.000 ;
        RECT 4.400 117.320 56.000 118.680 ;
        RECT 4.400 117.280 55.600 117.320 ;
        RECT 0.270 116.640 55.600 117.280 ;
        RECT 4.400 115.920 55.600 116.640 ;
        RECT 4.400 115.240 56.000 115.920 ;
        RECT 0.270 114.600 56.000 115.240 ;
        RECT 4.400 113.240 56.000 114.600 ;
        RECT 4.400 113.200 55.600 113.240 ;
        RECT 0.270 112.560 55.600 113.200 ;
        RECT 4.400 111.840 55.600 112.560 ;
        RECT 4.400 111.160 56.000 111.840 ;
        RECT 0.270 110.520 56.000 111.160 ;
        RECT 4.400 109.840 56.000 110.520 ;
        RECT 4.400 109.120 55.600 109.840 ;
        RECT 0.270 108.480 55.600 109.120 ;
        RECT 4.400 108.440 55.600 108.480 ;
        RECT 4.400 107.080 56.000 108.440 ;
        RECT 0.270 106.440 56.000 107.080 ;
        RECT 4.400 105.760 56.000 106.440 ;
        RECT 4.400 105.040 55.600 105.760 ;
        RECT 0.270 104.360 55.600 105.040 ;
        RECT 0.270 103.720 56.000 104.360 ;
        RECT 4.400 102.360 56.000 103.720 ;
        RECT 4.400 102.320 55.600 102.360 ;
        RECT 0.270 101.680 55.600 102.320 ;
        RECT 4.400 100.960 55.600 101.680 ;
        RECT 4.400 100.280 56.000 100.960 ;
        RECT 0.270 99.640 56.000 100.280 ;
        RECT 4.400 98.280 56.000 99.640 ;
        RECT 4.400 98.240 55.600 98.280 ;
        RECT 0.270 97.600 55.600 98.240 ;
        RECT 4.400 96.880 55.600 97.600 ;
        RECT 4.400 96.200 56.000 96.880 ;
        RECT 0.270 95.560 56.000 96.200 ;
        RECT 4.400 94.200 56.000 95.560 ;
        RECT 4.400 94.160 55.600 94.200 ;
        RECT 0.270 93.520 55.600 94.160 ;
        RECT 4.400 92.800 55.600 93.520 ;
        RECT 4.400 92.120 56.000 92.800 ;
        RECT 0.270 91.480 56.000 92.120 ;
        RECT 4.400 90.800 56.000 91.480 ;
        RECT 4.400 90.080 55.600 90.800 ;
        RECT 0.270 89.400 55.600 90.080 ;
        RECT 0.270 88.760 56.000 89.400 ;
        RECT 4.400 87.360 56.000 88.760 ;
        RECT 0.270 86.720 56.000 87.360 ;
        RECT 4.400 85.320 55.600 86.720 ;
        RECT 0.270 84.680 56.000 85.320 ;
        RECT 4.400 83.280 56.000 84.680 ;
        RECT 0.270 82.640 56.000 83.280 ;
        RECT 4.400 81.240 55.600 82.640 ;
        RECT 0.270 80.600 56.000 81.240 ;
        RECT 4.400 79.240 56.000 80.600 ;
        RECT 4.400 79.200 55.600 79.240 ;
        RECT 0.270 78.560 55.600 79.200 ;
        RECT 4.400 77.840 55.600 78.560 ;
        RECT 4.400 77.160 56.000 77.840 ;
        RECT 0.270 76.520 56.000 77.160 ;
        RECT 4.400 75.160 56.000 76.520 ;
        RECT 4.400 75.120 55.600 75.160 ;
        RECT 0.270 73.800 55.600 75.120 ;
        RECT 4.400 73.760 55.600 73.800 ;
        RECT 4.400 72.400 56.000 73.760 ;
        RECT 0.270 71.760 56.000 72.400 ;
        RECT 4.400 71.080 56.000 71.760 ;
        RECT 4.400 70.360 55.600 71.080 ;
        RECT 0.270 69.720 55.600 70.360 ;
        RECT 4.400 69.680 55.600 69.720 ;
        RECT 4.400 68.320 56.000 69.680 ;
        RECT 0.270 67.680 56.000 68.320 ;
        RECT 4.400 66.280 55.600 67.680 ;
        RECT 0.270 65.640 56.000 66.280 ;
        RECT 4.400 64.240 56.000 65.640 ;
        RECT 0.270 63.600 56.000 64.240 ;
        RECT 4.400 62.200 55.600 63.600 ;
        RECT 0.270 61.560 56.000 62.200 ;
        RECT 4.400 60.160 56.000 61.560 ;
        RECT 0.270 59.520 56.000 60.160 ;
        RECT 0.270 58.840 55.600 59.520 ;
        RECT 4.400 58.120 55.600 58.840 ;
        RECT 4.400 57.440 56.000 58.120 ;
        RECT 0.270 56.800 56.000 57.440 ;
        RECT 4.400 56.120 56.000 56.800 ;
        RECT 4.400 55.400 55.600 56.120 ;
        RECT 0.270 54.760 55.600 55.400 ;
        RECT 4.400 54.720 55.600 54.760 ;
        RECT 4.400 53.360 56.000 54.720 ;
        RECT 0.270 52.720 56.000 53.360 ;
        RECT 4.400 52.040 56.000 52.720 ;
        RECT 4.400 51.320 55.600 52.040 ;
        RECT 0.270 50.680 55.600 51.320 ;
        RECT 4.400 50.640 55.600 50.680 ;
        RECT 4.400 49.280 56.000 50.640 ;
        RECT 0.270 48.640 56.000 49.280 ;
        RECT 4.400 47.960 56.000 48.640 ;
        RECT 4.400 47.240 55.600 47.960 ;
        RECT 0.270 46.600 55.600 47.240 ;
        RECT 4.400 46.560 55.600 46.600 ;
        RECT 4.400 45.200 56.000 46.560 ;
        RECT 0.270 44.560 56.000 45.200 ;
        RECT 0.270 43.880 55.600 44.560 ;
        RECT 4.400 43.160 55.600 43.880 ;
        RECT 4.400 42.480 56.000 43.160 ;
        RECT 0.270 41.840 56.000 42.480 ;
        RECT 4.400 40.480 56.000 41.840 ;
        RECT 4.400 40.440 55.600 40.480 ;
        RECT 0.270 39.800 55.600 40.440 ;
        RECT 4.400 39.080 55.600 39.800 ;
        RECT 4.400 38.400 56.000 39.080 ;
        RECT 0.270 37.760 56.000 38.400 ;
        RECT 4.400 36.400 56.000 37.760 ;
        RECT 4.400 36.360 55.600 36.400 ;
        RECT 0.270 35.720 55.600 36.360 ;
        RECT 4.400 35.000 55.600 35.720 ;
        RECT 4.400 34.320 56.000 35.000 ;
        RECT 0.270 33.680 56.000 34.320 ;
        RECT 4.400 33.000 56.000 33.680 ;
        RECT 4.400 32.280 55.600 33.000 ;
        RECT 0.270 31.640 55.600 32.280 ;
        RECT 4.400 31.600 55.600 31.640 ;
        RECT 4.400 30.240 56.000 31.600 ;
        RECT 0.270 28.920 56.000 30.240 ;
        RECT 4.400 27.520 55.600 28.920 ;
        RECT 0.270 26.880 56.000 27.520 ;
        RECT 4.400 25.480 56.000 26.880 ;
        RECT 0.270 24.840 56.000 25.480 ;
        RECT 4.400 23.440 55.600 24.840 ;
        RECT 0.270 22.800 56.000 23.440 ;
        RECT 4.400 21.440 56.000 22.800 ;
        RECT 4.400 21.400 55.600 21.440 ;
        RECT 0.270 20.760 55.600 21.400 ;
        RECT 4.400 20.040 55.600 20.760 ;
        RECT 4.400 19.360 56.000 20.040 ;
        RECT 0.270 18.720 56.000 19.360 ;
        RECT 4.400 17.360 56.000 18.720 ;
        RECT 4.400 17.320 55.600 17.360 ;
        RECT 0.270 16.680 55.600 17.320 ;
        RECT 4.400 15.960 55.600 16.680 ;
        RECT 4.400 15.280 56.000 15.960 ;
        RECT 0.270 13.960 56.000 15.280 ;
        RECT 4.400 13.280 56.000 13.960 ;
        RECT 4.400 12.560 55.600 13.280 ;
        RECT 0.270 11.920 55.600 12.560 ;
        RECT 4.400 11.880 55.600 11.920 ;
        RECT 4.400 10.520 56.000 11.880 ;
        RECT 0.270 9.880 56.000 10.520 ;
        RECT 4.400 8.480 55.600 9.880 ;
        RECT 0.270 7.840 56.000 8.480 ;
        RECT 4.400 6.440 56.000 7.840 ;
        RECT 0.270 5.800 56.000 6.440 ;
        RECT 4.400 4.400 55.600 5.800 ;
        RECT 0.270 3.760 56.000 4.400 ;
        RECT 4.400 2.400 56.000 3.760 ;
        RECT 4.400 2.360 55.600 2.400 ;
        RECT 0.270 1.720 55.600 2.360 ;
        RECT 4.400 1.000 55.600 1.720 ;
        RECT 4.400 0.855 56.000 1.000 ;
      LAYER met4 ;
        RECT 0.295 23.975 12.480 375.185 ;
        RECT 14.880 23.975 20.640 375.185 ;
        RECT 23.040 23.975 28.800 375.185 ;
        RECT 31.200 23.975 36.960 375.185 ;
        RECT 39.360 23.975 42.025 375.185 ;
  END
END wb_bridge_2way
END LIBRARY

