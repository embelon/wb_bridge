magic
tech sky130A
magscale 1 2
timestamp 1647472436
<< viali >>
rect 2145 77673 2179 77707
rect 1409 77469 1443 77503
rect 2329 77469 2363 77503
rect 2973 77469 3007 77503
rect 3985 77469 4019 77503
rect 4629 77469 4663 77503
rect 9413 77469 9447 77503
rect 9965 77469 9999 77503
rect 10149 77401 10183 77435
rect 1593 77333 1627 77367
rect 2789 77333 2823 77367
rect 3801 77333 3835 77367
rect 4445 77333 4479 77367
rect 9229 77333 9263 77367
rect 4445 77129 4479 77163
rect 1685 77061 1719 77095
rect 1409 76993 1443 77027
rect 1593 76993 1627 77027
rect 1829 76993 1863 77027
rect 2697 76993 2731 77027
rect 3341 76993 3375 77027
rect 3985 76993 4019 77027
rect 4629 76993 4663 77027
rect 9413 76993 9447 77027
rect 9873 76993 9907 77027
rect 9229 76857 9263 76891
rect 1961 76789 1995 76823
rect 2513 76789 2547 76823
rect 3157 76789 3191 76823
rect 3801 76789 3835 76823
rect 10057 76789 10091 76823
rect 2789 76517 2823 76551
rect 9965 76517 9999 76551
rect 1593 76381 1627 76415
rect 2237 76381 2271 76415
rect 2657 76381 2691 76415
rect 3985 76381 4019 76415
rect 10149 76381 10183 76415
rect 2421 76313 2455 76347
rect 2513 76313 2547 76347
rect 1409 76245 1443 76279
rect 3801 76245 3835 76279
rect 1409 76041 1443 76075
rect 9965 76041 9999 76075
rect 2990 75973 3024 76007
rect 1593 75905 1627 75939
rect 2421 75905 2455 75939
rect 2605 75905 2639 75939
rect 2697 75905 2731 75939
rect 2794 75905 2828 75939
rect 3709 75905 3743 75939
rect 10149 75905 10183 75939
rect 3525 75701 3559 75735
rect 2513 75429 2547 75463
rect 9965 75429 9999 75463
rect 1961 75293 1995 75327
rect 2334 75293 2368 75327
rect 10149 75293 10183 75327
rect 2145 75225 2179 75259
rect 2237 75225 2271 75259
rect 1685 74885 1719 74919
rect 1409 74817 1443 74851
rect 1593 74817 1627 74851
rect 1829 74817 1863 74851
rect 2697 74817 2731 74851
rect 2513 74681 2547 74715
rect 1961 74613 1995 74647
rect 2513 74341 2547 74375
rect 9965 74341 9999 74375
rect 1961 74205 1995 74239
rect 2334 74205 2368 74239
rect 10149 74205 10183 74239
rect 2145 74137 2179 74171
rect 2237 74137 2271 74171
rect 1593 73729 1627 73763
rect 2237 73729 2271 73763
rect 2881 73729 2915 73763
rect 10149 73729 10183 73763
rect 1409 73525 1443 73559
rect 2053 73525 2087 73559
rect 2697 73525 2731 73559
rect 9965 73525 9999 73559
rect 1593 73117 1627 73151
rect 1409 72981 1443 73015
rect 1593 72709 1627 72743
rect 1685 72709 1719 72743
rect 1409 72641 1443 72675
rect 1829 72641 1863 72675
rect 2513 72641 2547 72675
rect 2697 72641 2731 72675
rect 2789 72641 2823 72675
rect 2933 72641 2967 72675
rect 10149 72641 10183 72675
rect 1961 72505 1995 72539
rect 3065 72437 3099 72471
rect 9965 72437 9999 72471
rect 9965 72233 9999 72267
rect 2697 72165 2731 72199
rect 1593 72029 1627 72063
rect 2237 72029 2271 72063
rect 2881 72029 2915 72063
rect 10149 72029 10183 72063
rect 1409 71893 1443 71927
rect 2053 71893 2087 71927
rect 1685 71621 1719 71655
rect 2697 71621 2731 71655
rect 2789 71621 2823 71655
rect 1409 71553 1443 71587
rect 1593 71553 1627 71587
rect 1829 71553 1863 71587
rect 2513 71553 2547 71587
rect 2933 71553 2967 71587
rect 3082 71553 3116 71587
rect 10149 71553 10183 71587
rect 9965 71417 9999 71451
rect 1961 71349 1995 71383
rect 1593 70941 1627 70975
rect 1409 70805 1443 70839
rect 1978 70601 2012 70635
rect 1593 70533 1627 70567
rect 1685 70533 1719 70567
rect 1409 70465 1443 70499
rect 1829 70465 1863 70499
rect 2697 70465 2731 70499
rect 10149 70465 10183 70499
rect 9965 70329 9999 70363
rect 2513 70261 2547 70295
rect 1593 69853 1627 69887
rect 2237 69853 2271 69887
rect 2881 69853 2915 69887
rect 10149 69853 10183 69887
rect 1409 69717 1443 69751
rect 2053 69717 2087 69751
rect 2697 69717 2731 69751
rect 9965 69717 9999 69751
rect 1685 69445 1719 69479
rect 1409 69377 1443 69411
rect 1593 69377 1627 69411
rect 1829 69377 1863 69411
rect 2697 69377 2731 69411
rect 1961 69241 1995 69275
rect 2513 69173 2547 69207
rect 9965 68969 9999 69003
rect 2881 68901 2915 68935
rect 1593 68765 1627 68799
rect 2329 68765 2363 68799
rect 2749 68765 2783 68799
rect 10149 68765 10183 68799
rect 2513 68697 2547 68731
rect 2605 68697 2639 68731
rect 1409 68629 1443 68663
rect 1685 68289 1719 68323
rect 10149 68289 10183 68323
rect 1409 68221 1443 68255
rect 9965 68085 9999 68119
rect 1409 67677 1443 67711
rect 1685 67677 1719 67711
rect 2881 67201 2915 67235
rect 10149 67201 10183 67235
rect 1409 67133 1443 67167
rect 1685 67133 1719 67167
rect 2697 67065 2731 67099
rect 9965 66997 9999 67031
rect 1961 66725 1995 66759
rect 1409 66589 1443 66623
rect 1829 66589 1863 66623
rect 2513 66589 2547 66623
rect 10149 66589 10183 66623
rect 1593 66521 1627 66555
rect 1686 66521 1720 66555
rect 2697 66453 2731 66487
rect 9965 66453 9999 66487
rect 1777 66181 1811 66215
rect 1501 66113 1535 66147
rect 1685 66113 1719 66147
rect 1874 66113 1908 66147
rect 2605 66113 2639 66147
rect 10149 66113 10183 66147
rect 2053 65977 2087 66011
rect 2789 65909 2823 65943
rect 9965 65909 9999 65943
rect 1593 65501 1627 65535
rect 2053 65501 2087 65535
rect 2329 65501 2363 65535
rect 2473 65501 2507 65535
rect 3801 65501 3835 65535
rect 2237 65433 2271 65467
rect 1409 65365 1443 65399
rect 2622 65365 2656 65399
rect 3985 65365 4019 65399
rect 1978 65093 2012 65127
rect 2697 65093 2731 65127
rect 2789 65093 2823 65127
rect 1409 65025 1443 65059
rect 1593 65025 1627 65059
rect 1685 65025 1719 65059
rect 1782 65025 1816 65059
rect 2513 65025 2547 65059
rect 2881 65025 2915 65059
rect 3525 65025 3559 65059
rect 10149 65025 10183 65059
rect 3709 64957 3743 64991
rect 3065 64889 3099 64923
rect 9965 64889 9999 64923
rect 2513 64549 2547 64583
rect 1961 64413 1995 64447
rect 2237 64413 2271 64447
rect 2381 64413 2415 64447
rect 3801 64413 3835 64447
rect 10149 64413 10183 64447
rect 2145 64345 2179 64379
rect 3985 64277 4019 64311
rect 9965 64277 9999 64311
rect 3801 64005 3835 64039
rect 1409 63937 1443 63971
rect 2605 63937 2639 63971
rect 3525 63937 3559 63971
rect 2881 63869 2915 63903
rect 1593 63733 1627 63767
rect 2329 63461 2363 63495
rect 3065 63461 3099 63495
rect 1409 63325 1443 63359
rect 2145 63325 2179 63359
rect 2881 63325 2915 63359
rect 10149 63325 10183 63359
rect 1593 63189 1627 63223
rect 9965 63189 9999 63223
rect 1409 62849 1443 62883
rect 2145 62849 2179 62883
rect 10149 62849 10183 62883
rect 1593 62645 1627 62679
rect 2329 62645 2363 62679
rect 9965 62645 9999 62679
rect 2513 62373 2547 62407
rect 1961 62237 1995 62271
rect 2237 62237 2271 62271
rect 2381 62237 2415 62271
rect 10149 62237 10183 62271
rect 2145 62169 2179 62203
rect 9965 62101 9999 62135
rect 1409 61761 1443 61795
rect 1593 61761 1627 61795
rect 1685 61761 1719 61795
rect 1782 61761 1816 61795
rect 2605 61761 2639 61795
rect 3525 61761 3559 61795
rect 2789 61693 2823 61727
rect 3709 61625 3743 61659
rect 1961 61557 1995 61591
rect 9965 61353 9999 61387
rect 1961 61285 1995 61319
rect 1409 61149 1443 61183
rect 1782 61149 1816 61183
rect 2513 61149 2547 61183
rect 10149 61149 10183 61183
rect 1593 61081 1627 61115
rect 1685 61081 1719 61115
rect 2697 61013 2731 61047
rect 1409 60673 1443 60707
rect 2145 60673 2179 60707
rect 2881 60673 2915 60707
rect 10149 60673 10183 60707
rect 3065 60537 3099 60571
rect 1593 60469 1627 60503
rect 2329 60469 2363 60503
rect 9965 60469 9999 60503
rect 2237 60061 2271 60095
rect 2789 60061 2823 60095
rect 2605 59925 2639 59959
rect 1593 59653 1627 59687
rect 1685 59653 1719 59687
rect 2329 59653 2363 59687
rect 2421 59653 2455 59687
rect 1409 59585 1443 59619
rect 1782 59585 1816 59619
rect 2145 59585 2179 59619
rect 2565 59585 2599 59619
rect 10149 59585 10183 59619
rect 1961 59381 1995 59415
rect 2697 59381 2731 59415
rect 9965 59381 9999 59415
rect 1409 59177 1443 59211
rect 2605 59109 2639 59143
rect 1593 58973 1627 59007
rect 2053 58973 2087 59007
rect 2329 58973 2363 59007
rect 2473 58973 2507 59007
rect 3801 58973 3835 59007
rect 10149 58973 10183 59007
rect 2237 58905 2271 58939
rect 3985 58837 4019 58871
rect 9965 58837 9999 58871
rect 2881 58633 2915 58667
rect 1409 58497 1443 58531
rect 2697 58497 2731 58531
rect 3341 58497 3375 58531
rect 9597 58497 9631 58531
rect 2513 58429 2547 58463
rect 9321 58429 9355 58463
rect 3525 58361 3559 58395
rect 1593 58293 1627 58327
rect 1409 57885 1443 57919
rect 2145 57885 2179 57919
rect 1593 57749 1627 57783
rect 2329 57749 2363 57783
rect 1685 57477 1719 57511
rect 1409 57409 1443 57443
rect 1593 57409 1627 57443
rect 1829 57409 1863 57443
rect 9597 57409 9631 57443
rect 9321 57341 9355 57375
rect 1961 57205 1995 57239
rect 2513 57001 2547 57035
rect 1961 56933 1995 56967
rect 9597 56865 9631 56899
rect 1409 56797 1443 56831
rect 1685 56797 1719 56831
rect 1782 56797 1816 56831
rect 2697 56797 2731 56831
rect 9321 56797 9355 56831
rect 1593 56729 1627 56763
rect 1593 56457 1627 56491
rect 3617 56457 3651 56491
rect 1409 56321 1443 56355
rect 2145 56321 2179 56355
rect 2881 56321 2915 56355
rect 3801 56321 3835 56355
rect 10149 56321 10183 56355
rect 3065 56185 3099 56219
rect 2329 56117 2363 56151
rect 9965 56117 9999 56151
rect 1409 55709 1443 55743
rect 2145 55709 2179 55743
rect 2881 55709 2915 55743
rect 3065 55709 3099 55743
rect 3801 55709 3835 55743
rect 3985 55709 4019 55743
rect 10149 55709 10183 55743
rect 1593 55573 1627 55607
rect 2329 55573 2363 55607
rect 3249 55573 3283 55607
rect 4169 55573 4203 55607
rect 9965 55573 9999 55607
rect 2789 55369 2823 55403
rect 3617 55369 3651 55403
rect 4445 55369 4479 55403
rect 1409 55233 1443 55267
rect 2605 55233 2639 55267
rect 3433 55233 3467 55267
rect 4261 55233 4295 55267
rect 10149 55233 10183 55267
rect 2421 55165 2455 55199
rect 3249 55165 3283 55199
rect 4077 55165 4111 55199
rect 1593 55029 1627 55063
rect 9965 55029 9999 55063
rect 1961 54757 1995 54791
rect 1409 54621 1443 54655
rect 1686 54621 1720 54655
rect 1823 54621 1857 54655
rect 2513 54621 2547 54655
rect 9505 54621 9539 54655
rect 10149 54621 10183 54655
rect 1593 54553 1627 54587
rect 2697 54485 2731 54519
rect 9321 54485 9355 54519
rect 9965 54485 9999 54519
rect 1409 54145 1443 54179
rect 1593 54145 1627 54179
rect 1685 54145 1719 54179
rect 1782 54145 1816 54179
rect 2513 54145 2547 54179
rect 9873 54145 9907 54179
rect 10057 54009 10091 54043
rect 1961 53941 1995 53975
rect 2697 53941 2731 53975
rect 1409 53533 1443 53567
rect 2145 53533 2179 53567
rect 9873 53533 9907 53567
rect 1593 53397 1627 53431
rect 2329 53397 2363 53431
rect 10057 53397 10091 53431
rect 1409 53057 1443 53091
rect 9873 53057 9907 53091
rect 1593 52853 1627 52887
rect 10057 52853 10091 52887
rect 2145 52649 2179 52683
rect 1409 52445 1443 52479
rect 2329 52445 2363 52479
rect 1593 52309 1627 52343
rect 3065 52105 3099 52139
rect 1409 51969 1443 52003
rect 2145 51969 2179 52003
rect 2881 51969 2915 52003
rect 9873 51969 9907 52003
rect 1593 51833 1627 51867
rect 2329 51765 2363 51799
rect 10057 51765 10091 51799
rect 2513 51561 2547 51595
rect 2973 51561 3007 51595
rect 1409 51357 1443 51391
rect 2237 51357 2271 51391
rect 2329 51357 2363 51391
rect 3157 51357 3191 51391
rect 9873 51357 9907 51391
rect 1593 51221 1627 51255
rect 10057 51221 10091 51255
rect 2881 51017 2915 51051
rect 9965 51017 9999 51051
rect 1593 50949 1627 50983
rect 1681 50949 1715 50983
rect 1409 50881 1443 50915
rect 1777 50881 1811 50915
rect 2697 50881 2731 50915
rect 3525 50881 3559 50915
rect 10149 50881 10183 50915
rect 2513 50813 2547 50847
rect 3341 50813 3375 50847
rect 1961 50677 1995 50711
rect 3709 50677 3743 50711
rect 1409 50269 1443 50303
rect 1593 50269 1627 50303
rect 1777 50269 1811 50303
rect 2421 50269 2455 50303
rect 9873 50269 9907 50303
rect 1685 50201 1719 50235
rect 1961 50133 1995 50167
rect 2605 50133 2639 50167
rect 10057 50133 10091 50167
rect 10057 49929 10091 49963
rect 1685 49861 1719 49895
rect 1409 49793 1443 49827
rect 1593 49793 1627 49827
rect 1777 49793 1811 49827
rect 2421 49793 2455 49827
rect 9873 49793 9907 49827
rect 1961 49657 1995 49691
rect 2605 49589 2639 49623
rect 9229 49385 9263 49419
rect 1409 49181 1443 49215
rect 2145 49181 2179 49215
rect 9413 49181 9447 49215
rect 9873 49181 9907 49215
rect 1593 49045 1627 49079
rect 2329 49045 2363 49079
rect 10057 49045 10091 49079
rect 9965 48841 9999 48875
rect 1409 48705 1443 48739
rect 2605 48705 2639 48739
rect 3617 48705 3651 48739
rect 3801 48705 3835 48739
rect 10149 48705 10183 48739
rect 2329 48637 2363 48671
rect 3985 48569 4019 48603
rect 1593 48501 1627 48535
rect 2789 48229 2823 48263
rect 9229 48229 9263 48263
rect 4629 48161 4663 48195
rect 1409 48093 1443 48127
rect 2421 48093 2455 48127
rect 2605 48093 2639 48127
rect 4353 48093 4387 48127
rect 4445 48093 4479 48127
rect 5089 48093 5123 48127
rect 5273 48093 5307 48127
rect 5457 48093 5491 48127
rect 7021 48093 7055 48127
rect 9413 48093 9447 48127
rect 9873 48093 9907 48127
rect 1593 47957 1627 47991
rect 6837 47957 6871 47991
rect 10057 47957 10091 47991
rect 1501 47617 1535 47651
rect 1593 47617 1627 47651
rect 2513 47617 2547 47651
rect 3525 47617 3559 47651
rect 9873 47617 9907 47651
rect 2237 47549 2271 47583
rect 1777 47413 1811 47447
rect 3709 47413 3743 47447
rect 10057 47413 10091 47447
rect 3157 47209 3191 47243
rect 7481 47209 7515 47243
rect 9965 47209 9999 47243
rect 1501 47073 1535 47107
rect 1777 47073 1811 47107
rect 2881 47005 2915 47039
rect 2973 47005 3007 47039
rect 3801 47005 3835 47039
rect 4997 47005 5031 47039
rect 5181 47005 5215 47039
rect 5365 47005 5399 47039
rect 7665 47005 7699 47039
rect 10149 47005 10183 47039
rect 3985 46869 4019 46903
rect 3249 46665 3283 46699
rect 1593 46529 1627 46563
rect 1777 46529 1811 46563
rect 3065 46529 3099 46563
rect 3709 46529 3743 46563
rect 9873 46529 9907 46563
rect 2881 46461 2915 46495
rect 3893 46393 3927 46427
rect 10057 46393 10091 46427
rect 1961 46325 1995 46359
rect 1409 45985 1443 46019
rect 1685 45985 1719 46019
rect 2697 45917 2731 45951
rect 3801 45917 3835 45951
rect 9873 45917 9907 45951
rect 2881 45781 2915 45815
rect 3985 45781 4019 45815
rect 10057 45781 10091 45815
rect 2145 45441 2179 45475
rect 1869 45373 1903 45407
rect 1593 45033 1627 45067
rect 2513 45033 2547 45067
rect 5641 45033 5675 45067
rect 1409 44829 1443 44863
rect 2237 44829 2271 44863
rect 2329 44829 2363 44863
rect 5825 44829 5859 44863
rect 9873 44829 9907 44863
rect 10057 44693 10091 44727
rect 1593 44489 1627 44523
rect 4905 44489 4939 44523
rect 1409 44353 1443 44387
rect 2973 44353 3007 44387
rect 3617 44353 3651 44387
rect 4721 44353 4755 44387
rect 9873 44353 9907 44387
rect 2789 44285 2823 44319
rect 4537 44285 4571 44319
rect 3157 44217 3191 44251
rect 3801 44149 3835 44183
rect 10057 44149 10091 44183
rect 9229 43945 9263 43979
rect 2513 43877 2547 43911
rect 1961 43741 1995 43775
rect 2237 43741 2271 43775
rect 2329 43741 2363 43775
rect 2973 43741 3007 43775
rect 3893 43741 3927 43775
rect 3985 43741 4019 43775
rect 4629 43741 4663 43775
rect 9413 43741 9447 43775
rect 9873 43741 9907 43775
rect 2145 43673 2179 43707
rect 4169 43673 4203 43707
rect 3157 43605 3191 43639
rect 4813 43605 4847 43639
rect 10057 43605 10091 43639
rect 1593 43401 1627 43435
rect 9965 43401 9999 43435
rect 1409 43265 1443 43299
rect 2145 43265 2179 43299
rect 2881 43265 2915 43299
rect 3801 43265 3835 43299
rect 10149 43265 10183 43299
rect 3157 43197 3191 43231
rect 2329 43061 2363 43095
rect 3985 43061 4019 43095
rect 1777 42721 1811 42755
rect 1501 42653 1535 42687
rect 2789 42653 2823 42687
rect 3801 42653 3835 42687
rect 9873 42653 9907 42687
rect 2973 42517 3007 42551
rect 3985 42517 4019 42551
rect 10057 42517 10091 42551
rect 3065 42313 3099 42347
rect 4261 42313 4295 42347
rect 1685 42177 1719 42211
rect 2881 42177 2915 42211
rect 3985 42177 4019 42211
rect 4077 42177 4111 42211
rect 4721 42177 4755 42211
rect 5641 42177 5675 42211
rect 9873 42177 9907 42211
rect 1409 42109 1443 42143
rect 2697 42109 2731 42143
rect 4905 42041 4939 42075
rect 5457 42041 5491 42075
rect 10057 41973 10091 42007
rect 4629 41769 4663 41803
rect 1777 41633 1811 41667
rect 4261 41633 4295 41667
rect 2053 41565 2087 41599
rect 4445 41565 4479 41599
rect 1961 41225 1995 41259
rect 2789 41225 2823 41259
rect 1777 41089 1811 41123
rect 2605 41089 2639 41123
rect 3249 41089 3283 41123
rect 4537 41089 4571 41123
rect 4721 41089 4755 41123
rect 5733 41089 5767 41123
rect 9873 41089 9907 41123
rect 1593 41021 1627 41055
rect 2421 41021 2455 41055
rect 4353 41021 4387 41055
rect 5549 40953 5583 40987
rect 10057 40953 10091 40987
rect 3433 40885 3467 40919
rect 9229 40681 9263 40715
rect 2329 40545 2363 40579
rect 2053 40477 2087 40511
rect 3801 40477 3835 40511
rect 9413 40477 9447 40511
rect 9873 40477 9907 40511
rect 3985 40341 4019 40375
rect 10057 40341 10091 40375
rect 6377 40137 6411 40171
rect 1685 40001 1719 40035
rect 1777 40001 1811 40035
rect 3709 40001 3743 40035
rect 4445 40001 4479 40035
rect 6561 40001 6595 40035
rect 9873 40001 9907 40035
rect 1961 39933 1995 39967
rect 2421 39933 2455 39967
rect 2697 39933 2731 39967
rect 4629 39865 4663 39899
rect 3893 39797 3927 39831
rect 10057 39797 10091 39831
rect 3157 39593 3191 39627
rect 5365 39593 5399 39627
rect 9965 39593 9999 39627
rect 4813 39525 4847 39559
rect 1501 39457 1535 39491
rect 1777 39389 1811 39423
rect 2789 39389 2823 39423
rect 2973 39389 3007 39423
rect 3801 39389 3835 39423
rect 3985 39389 4019 39423
rect 4629 39389 4663 39423
rect 5549 39389 5583 39423
rect 10149 39389 10183 39423
rect 4169 39321 4203 39355
rect 5089 39049 5123 39083
rect 1777 38913 1811 38947
rect 3065 38913 3099 38947
rect 4905 38913 4939 38947
rect 9873 38913 9907 38947
rect 1501 38845 1535 38879
rect 2789 38845 2823 38879
rect 4721 38845 4755 38879
rect 10057 38709 10091 38743
rect 2881 38505 2915 38539
rect 4629 38505 4663 38539
rect 1409 38301 1443 38335
rect 2605 38301 2639 38335
rect 2697 38301 2731 38335
rect 4261 38301 4295 38335
rect 4445 38301 4479 38335
rect 9873 38301 9907 38335
rect 1593 38165 1627 38199
rect 10057 38165 10091 38199
rect 1961 37961 1995 37995
rect 2789 37961 2823 37995
rect 9965 37961 9999 37995
rect 1685 37825 1719 37859
rect 1777 37825 1811 37859
rect 2605 37825 2639 37859
rect 3249 37825 3283 37859
rect 3985 37825 4019 37859
rect 10149 37825 10183 37859
rect 2421 37757 2455 37791
rect 4169 37689 4203 37723
rect 3433 37621 3467 37655
rect 2789 37417 2823 37451
rect 3985 37349 4019 37383
rect 1409 37213 1443 37247
rect 3801 37213 3835 37247
rect 9873 37213 9907 37247
rect 2697 37145 2731 37179
rect 1593 37077 1627 37111
rect 10057 37077 10091 37111
rect 1869 36873 1903 36907
rect 2973 36873 3007 36907
rect 4629 36873 4663 36907
rect 1777 36805 1811 36839
rect 2421 36737 2455 36771
rect 3249 36737 3283 36771
rect 4445 36737 4479 36771
rect 9873 36737 9907 36771
rect 2237 36669 2271 36703
rect 4261 36669 4295 36703
rect 3433 36601 3467 36635
rect 2605 36533 2639 36567
rect 10057 36533 10091 36567
rect 2973 36329 3007 36363
rect 9229 36329 9263 36363
rect 1777 36193 1811 36227
rect 1501 36125 1535 36159
rect 2881 36125 2915 36159
rect 9413 36125 9447 36159
rect 9873 36125 9907 36159
rect 10057 35989 10091 36023
rect 4997 35785 5031 35819
rect 9965 35785 9999 35819
rect 3709 35717 3743 35751
rect 4077 35717 4111 35751
rect 1409 35649 1443 35683
rect 2145 35649 2179 35683
rect 4813 35649 4847 35683
rect 10149 35649 10183 35683
rect 4629 35581 4663 35615
rect 2329 35513 2363 35547
rect 1593 35445 1627 35479
rect 1961 35241 1995 35275
rect 4905 35241 4939 35275
rect 1593 35037 1627 35071
rect 1777 35037 1811 35071
rect 2421 35037 2455 35071
rect 4537 35037 4571 35071
rect 4721 35037 4755 35071
rect 9873 35037 9907 35071
rect 2605 34901 2639 34935
rect 10057 34901 10091 34935
rect 1593 34697 1627 34731
rect 10057 34697 10091 34731
rect 4353 34629 4387 34663
rect 1409 34561 1443 34595
rect 2145 34561 2179 34595
rect 2881 34561 2915 34595
rect 4169 34561 4203 34595
rect 9873 34561 9907 34595
rect 3985 34493 4019 34527
rect 2329 34357 2363 34391
rect 3065 34357 3099 34391
rect 9965 34153 9999 34187
rect 2053 34085 2087 34119
rect 3801 34085 3835 34119
rect 2697 33949 2731 33983
rect 2901 33951 2935 33985
rect 3065 33949 3099 33983
rect 3985 33949 4019 33983
rect 10149 33949 10183 33983
rect 1869 33881 1903 33915
rect 2237 33609 2271 33643
rect 2881 33609 2915 33643
rect 4537 33609 4571 33643
rect 1961 33473 1995 33507
rect 2053 33473 2087 33507
rect 2789 33473 2823 33507
rect 4353 33473 4387 33507
rect 9873 33473 9907 33507
rect 4169 33405 4203 33439
rect 10057 33337 10091 33371
rect 3801 33065 3835 33099
rect 1409 32861 1443 32895
rect 2145 32861 2179 32895
rect 2881 32861 2915 32895
rect 3985 32861 4019 32895
rect 9873 32861 9907 32895
rect 1593 32725 1627 32759
rect 2329 32725 2363 32759
rect 3065 32725 3099 32759
rect 10057 32725 10091 32759
rect 2421 32521 2455 32555
rect 3617 32521 3651 32555
rect 2237 32385 2271 32419
rect 2881 32385 2915 32419
rect 3801 32385 3835 32419
rect 4445 32385 4479 32419
rect 2053 32317 2087 32351
rect 3065 32249 3099 32283
rect 4261 32249 4295 32283
rect 1961 31977 1995 32011
rect 4537 31977 4571 32011
rect 2789 31909 2823 31943
rect 3985 31909 4019 31943
rect 10057 31909 10091 31943
rect 3801 31773 3835 31807
rect 4721 31773 4755 31807
rect 9873 31773 9907 31807
rect 1869 31705 1903 31739
rect 2605 31705 2639 31739
rect 1961 31433 1995 31467
rect 3893 31433 3927 31467
rect 1777 31297 1811 31331
rect 2881 31297 2915 31331
rect 3709 31297 3743 31331
rect 9873 31297 9907 31331
rect 1593 31229 1627 31263
rect 2697 31229 2731 31263
rect 3525 31229 3559 31263
rect 3065 31161 3099 31195
rect 10057 31093 10091 31127
rect 1961 30889 1995 30923
rect 2513 30685 2547 30719
rect 9873 30685 9907 30719
rect 1869 30617 1903 30651
rect 2697 30549 2731 30583
rect 10057 30549 10091 30583
rect 1869 30277 1903 30311
rect 2697 30277 2731 30311
rect 1685 30209 1719 30243
rect 2513 30209 2547 30243
rect 3157 30209 3191 30243
rect 4077 30209 4111 30243
rect 4721 30209 4755 30243
rect 2329 30141 2363 30175
rect 3341 30073 3375 30107
rect 4537 30073 4571 30107
rect 3893 30005 3927 30039
rect 2697 29801 2731 29835
rect 7665 29801 7699 29835
rect 2053 29597 2087 29631
rect 7849 29597 7883 29631
rect 10149 29597 10183 29631
rect 1869 29529 1903 29563
rect 2605 29529 2639 29563
rect 2145 29257 2179 29291
rect 2881 29257 2915 29291
rect 2053 29189 2087 29223
rect 2789 29121 2823 29155
rect 10149 28985 10183 29019
rect 1961 28713 1995 28747
rect 4077 28645 4111 28679
rect 2789 28577 2823 28611
rect 1869 28509 1903 28543
rect 2605 28441 2639 28475
rect 3893 28441 3927 28475
rect 3065 28169 3099 28203
rect 4261 28169 4295 28203
rect 1685 28033 1719 28067
rect 2881 28033 2915 28067
rect 3617 28033 3651 28067
rect 4445 28033 4479 28067
rect 1409 27965 1443 27999
rect 2697 27965 2731 27999
rect 3801 27965 3835 27999
rect 9965 27965 9999 27999
rect 3065 27557 3099 27591
rect 4445 27557 4479 27591
rect 1409 27489 1443 27523
rect 2697 27489 2731 27523
rect 1685 27421 1719 27455
rect 2881 27421 2915 27455
rect 4261 27353 4295 27387
rect 9965 27285 9999 27319
rect 3065 27081 3099 27115
rect 3709 27081 3743 27115
rect 2053 26945 2087 26979
rect 2881 26945 2915 26979
rect 3617 26945 3651 26979
rect 1869 26877 1903 26911
rect 2697 26877 2731 26911
rect 2237 26741 2271 26775
rect 10149 26741 10183 26775
rect 1961 26537 1995 26571
rect 2789 26469 2823 26503
rect 4445 26469 4479 26503
rect 1869 26333 1903 26367
rect 2605 26265 2639 26299
rect 4261 26265 4295 26299
rect 3065 25993 3099 26027
rect 1685 25857 1719 25891
rect 2881 25857 2915 25891
rect 1409 25789 1443 25823
rect 2697 25789 2731 25823
rect 10149 25653 10183 25687
rect 3157 25449 3191 25483
rect 1685 25313 1719 25347
rect 1409 25245 1443 25279
rect 2789 25245 2823 25279
rect 2973 25245 3007 25279
rect 10149 25245 10183 25279
rect 1869 24769 1903 24803
rect 2605 24769 2639 24803
rect 2789 24769 2823 24803
rect 3341 24769 3375 24803
rect 3525 24769 3559 24803
rect 1961 24565 1995 24599
rect 1685 24225 1719 24259
rect 2973 24225 3007 24259
rect 1409 24157 1443 24191
rect 10149 24157 10183 24191
rect 2789 24089 2823 24123
rect 1685 23681 1719 23715
rect 2973 23681 3007 23715
rect 1409 23613 1443 23647
rect 2697 23613 2731 23647
rect 10149 23477 10183 23511
rect 3065 23273 3099 23307
rect 1685 23137 1719 23171
rect 1409 23069 1443 23103
rect 2697 23069 2731 23103
rect 2881 23069 2915 23103
rect 3065 22729 3099 22763
rect 4537 22661 4571 22695
rect 1685 22593 1719 22627
rect 2881 22593 2915 22627
rect 3617 22593 3651 22627
rect 4353 22593 4387 22627
rect 1409 22525 1443 22559
rect 2697 22525 2731 22559
rect 10149 22457 10183 22491
rect 3709 22389 3743 22423
rect 10149 22117 10183 22151
rect 1685 22049 1719 22083
rect 3065 22049 3099 22083
rect 4169 22049 4203 22083
rect 1409 21981 1443 22015
rect 2697 21981 2731 22015
rect 2881 21981 2915 22015
rect 3801 21981 3835 22015
rect 3985 21981 4019 22015
rect 3985 21641 4019 21675
rect 2789 21573 2823 21607
rect 1685 21505 1719 21539
rect 3801 21505 3835 21539
rect 1409 21437 1443 21471
rect 3617 21437 3651 21471
rect 2973 21369 3007 21403
rect 10149 21301 10183 21335
rect 3065 21097 3099 21131
rect 1685 20961 1719 20995
rect 1409 20893 1443 20927
rect 2697 20893 2731 20927
rect 2881 20893 2915 20927
rect 3065 20553 3099 20587
rect 1685 20417 1719 20451
rect 2881 20417 2915 20451
rect 9873 20417 9907 20451
rect 1409 20349 1443 20383
rect 2697 20349 2731 20383
rect 10057 20281 10091 20315
rect 2605 20009 2639 20043
rect 3801 20009 3835 20043
rect 1777 19805 1811 19839
rect 1961 19805 1995 19839
rect 2789 19805 2823 19839
rect 3985 19805 4019 19839
rect 9873 19805 9907 19839
rect 2145 19669 2179 19703
rect 10057 19669 10091 19703
rect 1961 19465 1995 19499
rect 2513 19465 2547 19499
rect 9873 19465 9907 19499
rect 1869 19397 1903 19431
rect 2697 19329 2731 19363
rect 10057 19329 10091 19363
rect 1409 18921 1443 18955
rect 2053 18921 2087 18955
rect 2697 18921 2731 18955
rect 1593 18717 1627 18751
rect 2237 18717 2271 18751
rect 2881 18717 2915 18751
rect 9873 18717 9907 18751
rect 10057 18581 10091 18615
rect 1409 18377 1443 18411
rect 9229 18377 9263 18411
rect 2329 18309 2363 18343
rect 2545 18309 2579 18343
rect 1593 18241 1627 18275
rect 9413 18241 9447 18275
rect 9873 18241 9907 18275
rect 2513 18037 2547 18071
rect 2697 18037 2731 18071
rect 10057 18037 10091 18071
rect 1409 17833 1443 17867
rect 2421 17765 2455 17799
rect 4905 17697 4939 17731
rect 1593 17629 1627 17663
rect 2237 17629 2271 17663
rect 2789 17629 2823 17663
rect 2973 17629 3007 17663
rect 9873 17629 9907 17663
rect 4169 17561 4203 17595
rect 10057 17493 10091 17527
rect 3065 17289 3099 17323
rect 9965 17289 9999 17323
rect 2881 17221 2915 17255
rect 1593 17153 1627 17187
rect 10149 17153 10183 17187
rect 2513 17017 2547 17051
rect 1409 16949 1443 16983
rect 2881 16949 2915 16983
rect 1961 16745 1995 16779
rect 2697 16541 2731 16575
rect 3985 16541 4019 16575
rect 9873 16541 9907 16575
rect 1869 16473 1903 16507
rect 2513 16405 2547 16439
rect 3801 16405 3835 16439
rect 10057 16405 10091 16439
rect 2789 16201 2823 16235
rect 9229 16201 9263 16235
rect 1501 16065 1535 16099
rect 1593 16065 1627 16099
rect 1961 16065 1995 16099
rect 2605 16065 2639 16099
rect 9413 16065 9447 16099
rect 9873 16065 9907 16099
rect 1869 15861 1903 15895
rect 2145 15861 2179 15895
rect 10057 15861 10091 15895
rect 1869 15657 1903 15691
rect 2237 15657 2271 15691
rect 3801 15657 3835 15691
rect 9965 15657 9999 15691
rect 1961 15521 1995 15555
rect 1869 15453 1903 15487
rect 2881 15453 2915 15487
rect 3985 15453 4019 15487
rect 10149 15453 10183 15487
rect 2697 15317 2731 15351
rect 2145 15113 2179 15147
rect 2973 15045 3007 15079
rect 2053 14977 2087 15011
rect 2789 14977 2823 15011
rect 9873 14977 9907 15011
rect 10057 14841 10091 14875
rect 1685 14569 1719 14603
rect 1869 14569 1903 14603
rect 2789 14569 2823 14603
rect 2973 14569 3007 14603
rect 3801 14501 3835 14535
rect 1593 14433 1627 14467
rect 1685 14365 1719 14399
rect 3985 14365 4019 14399
rect 9873 14365 9907 14399
rect 1409 14297 1443 14331
rect 2605 14297 2639 14331
rect 2821 14297 2855 14331
rect 10057 14229 10091 14263
rect 1409 14025 1443 14059
rect 2421 14025 2455 14059
rect 3065 14025 3099 14059
rect 10057 14025 10091 14059
rect 1593 13889 1627 13923
rect 2237 13889 2271 13923
rect 3249 13889 3283 13923
rect 3893 13889 3927 13923
rect 9873 13889 9907 13923
rect 2053 13821 2087 13855
rect 3709 13753 3743 13787
rect 9965 13481 9999 13515
rect 3801 13413 3835 13447
rect 1593 13277 1627 13311
rect 2605 13277 2639 13311
rect 3249 13277 3283 13311
rect 3985 13277 4019 13311
rect 9505 13277 9539 13311
rect 10149 13277 10183 13311
rect 1409 13141 1443 13175
rect 2421 13141 2455 13175
rect 3065 13141 3099 13175
rect 9321 13141 9355 13175
rect 1409 12937 1443 12971
rect 2789 12937 2823 12971
rect 2973 12937 3007 12971
rect 9229 12937 9263 12971
rect 1593 12801 1627 12835
rect 2605 12801 2639 12835
rect 2697 12801 2731 12835
rect 9413 12801 9447 12835
rect 9873 12801 9907 12835
rect 2421 12665 2455 12699
rect 10057 12597 10091 12631
rect 1409 12393 1443 12427
rect 1869 12393 1903 12427
rect 9229 12393 9263 12427
rect 3065 12325 3099 12359
rect 1593 12257 1627 12291
rect 1409 12189 1443 12223
rect 1685 12189 1719 12223
rect 2329 12189 2363 12223
rect 3249 12189 3283 12223
rect 9413 12189 9447 12223
rect 9873 12189 9907 12223
rect 2513 12053 2547 12087
rect 10057 12053 10091 12087
rect 2881 11849 2915 11883
rect 3433 11849 3467 11883
rect 1685 11713 1719 11747
rect 2697 11713 2731 11747
rect 3617 11713 3651 11747
rect 1409 11645 1443 11679
rect 2881 11305 2915 11339
rect 3801 11237 3835 11271
rect 10057 11237 10091 11271
rect 1685 11169 1719 11203
rect 1409 11101 1443 11135
rect 2697 11101 2731 11135
rect 3985 11101 4019 11135
rect 9873 11101 9907 11135
rect 3433 10761 3467 10795
rect 2697 10625 2731 10659
rect 3617 10625 3651 10659
rect 9873 10625 9907 10659
rect 1409 10557 1443 10591
rect 1685 10557 1719 10591
rect 2881 10489 2915 10523
rect 10057 10421 10091 10455
rect 3065 10217 3099 10251
rect 1685 10081 1719 10115
rect 1409 10013 1443 10047
rect 2789 10013 2823 10047
rect 2881 10013 2915 10047
rect 1685 9537 1719 9571
rect 2697 9537 2731 9571
rect 3617 9537 3651 9571
rect 9873 9537 9907 9571
rect 1409 9469 1443 9503
rect 2881 9401 2915 9435
rect 10057 9401 10091 9435
rect 3433 9333 3467 9367
rect 2881 9129 2915 9163
rect 1685 8993 1719 9027
rect 1409 8925 1443 8959
rect 2697 8925 2731 8959
rect 3985 8925 4019 8959
rect 9873 8925 9907 8959
rect 3801 8789 3835 8823
rect 10057 8789 10091 8823
rect 3065 8585 3099 8619
rect 3525 8585 3559 8619
rect 1685 8449 1719 8483
rect 2881 8449 2915 8483
rect 3709 8449 3743 8483
rect 9873 8449 9907 8483
rect 1409 8381 1443 8415
rect 2697 8381 2731 8415
rect 10057 8313 10091 8347
rect 1685 7905 1719 7939
rect 1409 7837 1443 7871
rect 2881 7837 2915 7871
rect 2697 7701 2731 7735
rect 1593 7497 1627 7531
rect 2421 7429 2455 7463
rect 1409 7361 1443 7395
rect 2237 7361 2271 7395
rect 4077 7361 4111 7395
rect 9873 7361 9907 7395
rect 3893 7225 3927 7259
rect 10057 7157 10091 7191
rect 2421 6817 2455 6851
rect 1409 6749 1443 6783
rect 3065 6749 3099 6783
rect 9873 6749 9907 6783
rect 2237 6681 2271 6715
rect 1593 6613 1627 6647
rect 2881 6613 2915 6647
rect 10057 6613 10091 6647
rect 2513 6409 2547 6443
rect 2053 6341 2087 6375
rect 1869 6273 1903 6307
rect 2697 6273 2731 6307
rect 3341 6273 3375 6307
rect 3157 6137 3191 6171
rect 3065 5865 3099 5899
rect 1685 5729 1719 5763
rect 3801 5729 3835 5763
rect 1409 5661 1443 5695
rect 2789 5661 2823 5695
rect 2881 5661 2915 5695
rect 3985 5661 4019 5695
rect 9873 5661 9907 5695
rect 4169 5525 4203 5559
rect 10057 5525 10091 5559
rect 3709 5321 3743 5355
rect 9229 5321 9263 5355
rect 1409 5185 1443 5219
rect 1685 5185 1719 5219
rect 2881 5185 2915 5219
rect 3525 5185 3559 5219
rect 9413 5185 9447 5219
rect 9873 5185 9907 5219
rect 2697 5117 2731 5151
rect 3065 5049 3099 5083
rect 10057 4981 10091 5015
rect 3985 4777 4019 4811
rect 2053 4641 2087 4675
rect 1777 4573 1811 4607
rect 1869 4573 1903 4607
rect 2881 4573 2915 4607
rect 2973 4573 3007 4607
rect 3801 4573 3835 4607
rect 4721 4573 4755 4607
rect 9873 4573 9907 4607
rect 3157 4505 3191 4539
rect 4537 4437 4571 4471
rect 10057 4437 10091 4471
rect 9965 4233 9999 4267
rect 1685 4097 1719 4131
rect 2881 4097 2915 4131
rect 3709 4097 3743 4131
rect 4537 4097 4571 4131
rect 5181 4097 5215 4131
rect 10149 4097 10183 4131
rect 1409 4029 1443 4063
rect 2697 4029 2731 4063
rect 3525 4029 3559 4063
rect 3893 4029 3927 4063
rect 4353 3961 4387 3995
rect 3065 3893 3099 3927
rect 4997 3893 5031 3927
rect 2237 3689 2271 3723
rect 4169 3689 4203 3723
rect 1869 3553 1903 3587
rect 2053 3485 2087 3519
rect 2881 3485 2915 3519
rect 3801 3485 3835 3519
rect 3985 3485 4019 3519
rect 9873 3485 9907 3519
rect 2697 3349 2731 3383
rect 10057 3349 10091 3383
rect 1593 3145 1627 3179
rect 2789 3145 2823 3179
rect 4261 3145 4295 3179
rect 1409 3009 1443 3043
rect 2329 3009 2363 3043
rect 2973 3009 3007 3043
rect 3801 3009 3835 3043
rect 4445 3009 4479 3043
rect 5089 3009 5123 3043
rect 9137 3009 9171 3043
rect 9873 3009 9907 3043
rect 2145 2873 2179 2907
rect 3617 2873 3651 2907
rect 4905 2805 4939 2839
rect 9321 2805 9355 2839
rect 10057 2805 10091 2839
rect 2697 2601 2731 2635
rect 4445 2601 4479 2635
rect 3801 2533 3835 2567
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 2881 2397 2915 2431
rect 3985 2397 4019 2431
rect 4629 2397 4663 2431
rect 5273 2397 5307 2431
rect 9137 2397 9171 2431
rect 9873 2397 9907 2431
rect 5089 2261 5123 2295
rect 9321 2261 9355 2295
rect 10057 2261 10091 2295
<< metal1 >>
rect 1104 77818 10856 77840
rect 1104 77766 2582 77818
rect 2634 77766 2646 77818
rect 2698 77766 2710 77818
rect 2762 77766 2774 77818
rect 2826 77766 2838 77818
rect 2890 77766 5846 77818
rect 5898 77766 5910 77818
rect 5962 77766 5974 77818
rect 6026 77766 6038 77818
rect 6090 77766 6102 77818
rect 6154 77766 9110 77818
rect 9162 77766 9174 77818
rect 9226 77766 9238 77818
rect 9290 77766 9302 77818
rect 9354 77766 9366 77818
rect 9418 77766 10856 77818
rect 1104 77744 10856 77766
rect 2133 77707 2191 77713
rect 2133 77673 2145 77707
rect 2179 77704 2191 77707
rect 3510 77704 3516 77716
rect 2179 77676 3516 77704
rect 2179 77673 2191 77676
rect 2133 77667 2191 77673
rect 3510 77664 3516 77676
rect 3568 77664 3574 77716
rect 2958 77636 2964 77648
rect 2332 77608 2964 77636
rect 1394 77500 1400 77512
rect 1355 77472 1400 77500
rect 1394 77460 1400 77472
rect 1452 77460 1458 77512
rect 2332 77509 2360 77608
rect 2958 77596 2964 77608
rect 3016 77596 3022 77648
rect 2317 77503 2375 77509
rect 2317 77469 2329 77503
rect 2363 77469 2375 77503
rect 2958 77500 2964 77512
rect 2919 77472 2964 77500
rect 2317 77463 2375 77469
rect 2958 77460 2964 77472
rect 3016 77460 3022 77512
rect 3970 77500 3976 77512
rect 3931 77472 3976 77500
rect 3970 77460 3976 77472
rect 4028 77460 4034 77512
rect 4062 77460 4068 77512
rect 4120 77500 4126 77512
rect 4617 77503 4675 77509
rect 4617 77500 4629 77503
rect 4120 77472 4629 77500
rect 4120 77460 4126 77472
rect 4617 77469 4629 77472
rect 4663 77469 4675 77503
rect 9398 77500 9404 77512
rect 9359 77472 9404 77500
rect 4617 77463 4675 77469
rect 9398 77460 9404 77472
rect 9456 77460 9462 77512
rect 9950 77500 9956 77512
rect 9911 77472 9956 77500
rect 9950 77460 9956 77472
rect 10008 77460 10014 77512
rect 7834 77392 7840 77444
rect 7892 77432 7898 77444
rect 10137 77435 10195 77441
rect 10137 77432 10149 77435
rect 7892 77404 10149 77432
rect 7892 77392 7898 77404
rect 10137 77401 10149 77404
rect 10183 77401 10195 77435
rect 10137 77395 10195 77401
rect 1581 77367 1639 77373
rect 1581 77333 1593 77367
rect 1627 77364 1639 77367
rect 2038 77364 2044 77376
rect 1627 77336 2044 77364
rect 1627 77333 1639 77336
rect 1581 77327 1639 77333
rect 2038 77324 2044 77336
rect 2096 77324 2102 77376
rect 2777 77367 2835 77373
rect 2777 77333 2789 77367
rect 2823 77364 2835 77367
rect 2866 77364 2872 77376
rect 2823 77336 2872 77364
rect 2823 77333 2835 77336
rect 2777 77327 2835 77333
rect 2866 77324 2872 77336
rect 2924 77324 2930 77376
rect 3142 77324 3148 77376
rect 3200 77364 3206 77376
rect 3789 77367 3847 77373
rect 3789 77364 3801 77367
rect 3200 77336 3801 77364
rect 3200 77324 3206 77336
rect 3789 77333 3801 77336
rect 3835 77333 3847 77367
rect 3789 77327 3847 77333
rect 3878 77324 3884 77376
rect 3936 77364 3942 77376
rect 4433 77367 4491 77373
rect 4433 77364 4445 77367
rect 3936 77336 4445 77364
rect 3936 77324 3942 77336
rect 4433 77333 4445 77336
rect 4479 77333 4491 77367
rect 4433 77327 4491 77333
rect 8294 77324 8300 77376
rect 8352 77364 8358 77376
rect 9217 77367 9275 77373
rect 9217 77364 9229 77367
rect 8352 77336 9229 77364
rect 8352 77324 8358 77336
rect 9217 77333 9229 77336
rect 9263 77333 9275 77367
rect 9217 77327 9275 77333
rect 1104 77274 10856 77296
rect 1104 77222 4214 77274
rect 4266 77222 4278 77274
rect 4330 77222 4342 77274
rect 4394 77222 4406 77274
rect 4458 77222 4470 77274
rect 4522 77222 7478 77274
rect 7530 77222 7542 77274
rect 7594 77222 7606 77274
rect 7658 77222 7670 77274
rect 7722 77222 7734 77274
rect 7786 77222 10856 77274
rect 1104 77200 10856 77222
rect 4433 77163 4491 77169
rect 4433 77160 4445 77163
rect 1688 77132 4445 77160
rect 1688 77101 1716 77132
rect 4433 77129 4445 77132
rect 4479 77129 4491 77163
rect 4433 77123 4491 77129
rect 1673 77095 1731 77101
rect 1673 77061 1685 77095
rect 1719 77061 1731 77095
rect 1673 77055 1731 77061
rect 3694 77052 3700 77104
rect 3752 77092 3758 77104
rect 3752 77064 4660 77092
rect 3752 77052 3758 77064
rect 1397 77027 1455 77033
rect 1397 76993 1409 77027
rect 1443 76993 1455 77027
rect 1397 76987 1455 76993
rect 1412 76956 1440 76987
rect 1486 76984 1492 77036
rect 1544 77024 1550 77036
rect 1581 77027 1639 77033
rect 1581 77024 1593 77027
rect 1544 76996 1593 77024
rect 1544 76984 1550 76996
rect 1581 76993 1593 76996
rect 1627 76993 1639 77027
rect 1581 76987 1639 76993
rect 1817 77027 1875 77033
rect 1817 76993 1829 77027
rect 1863 77024 1875 77027
rect 2314 77024 2320 77036
rect 1863 76996 2320 77024
rect 1863 76993 1875 76996
rect 1817 76987 1875 76993
rect 2314 76984 2320 76996
rect 2372 76984 2378 77036
rect 2498 76984 2504 77036
rect 2556 77024 2562 77036
rect 2685 77027 2743 77033
rect 2685 77024 2697 77027
rect 2556 76996 2697 77024
rect 2556 76984 2562 76996
rect 2685 76993 2697 76996
rect 2731 76993 2743 77027
rect 3326 77024 3332 77036
rect 3287 76996 3332 77024
rect 2685 76987 2743 76993
rect 3326 76984 3332 76996
rect 3384 76984 3390 77036
rect 3418 76984 3424 77036
rect 3476 77024 3482 77036
rect 4632 77033 4660 77064
rect 3973 77027 4031 77033
rect 3973 77024 3985 77027
rect 3476 76996 3985 77024
rect 3476 76984 3482 76996
rect 3973 76993 3985 76996
rect 4019 76993 4031 77027
rect 3973 76987 4031 76993
rect 4617 77027 4675 77033
rect 4617 76993 4629 77027
rect 4663 76993 4675 77027
rect 4617 76987 4675 76993
rect 9401 77027 9459 77033
rect 9401 76993 9413 77027
rect 9447 77024 9459 77027
rect 9490 77024 9496 77036
rect 9447 76996 9496 77024
rect 9447 76993 9459 76996
rect 9401 76987 9459 76993
rect 9490 76984 9496 76996
rect 9548 76984 9554 77036
rect 9582 76984 9588 77036
rect 9640 77024 9646 77036
rect 9861 77027 9919 77033
rect 9861 77024 9873 77027
rect 9640 76996 9873 77024
rect 9640 76984 9646 76996
rect 9861 76993 9873 76996
rect 9907 76993 9919 77027
rect 9861 76987 9919 76993
rect 1412 76928 2774 76956
rect 2746 76888 2774 76928
rect 3050 76916 3056 76968
rect 3108 76956 3114 76968
rect 3602 76956 3608 76968
rect 3108 76928 3608 76956
rect 3108 76916 3114 76928
rect 3602 76916 3608 76928
rect 3660 76916 3666 76968
rect 9217 76891 9275 76897
rect 9217 76888 9229 76891
rect 2746 76860 9229 76888
rect 9217 76857 9229 76860
rect 9263 76857 9275 76891
rect 9217 76851 9275 76857
rect 1946 76820 1952 76832
rect 1907 76792 1952 76820
rect 1946 76780 1952 76792
rect 2004 76780 2010 76832
rect 2406 76780 2412 76832
rect 2464 76820 2470 76832
rect 2501 76823 2559 76829
rect 2501 76820 2513 76823
rect 2464 76792 2513 76820
rect 2464 76780 2470 76792
rect 2501 76789 2513 76792
rect 2547 76789 2559 76823
rect 2501 76783 2559 76789
rect 3050 76780 3056 76832
rect 3108 76820 3114 76832
rect 3145 76823 3203 76829
rect 3145 76820 3157 76823
rect 3108 76792 3157 76820
rect 3108 76780 3114 76792
rect 3145 76789 3157 76792
rect 3191 76789 3203 76823
rect 3145 76783 3203 76789
rect 3234 76780 3240 76832
rect 3292 76820 3298 76832
rect 3789 76823 3847 76829
rect 3789 76820 3801 76823
rect 3292 76792 3801 76820
rect 3292 76780 3298 76792
rect 3789 76789 3801 76792
rect 3835 76789 3847 76823
rect 3789 76783 3847 76789
rect 9766 76780 9772 76832
rect 9824 76820 9830 76832
rect 10045 76823 10103 76829
rect 10045 76820 10057 76823
rect 9824 76792 10057 76820
rect 9824 76780 9830 76792
rect 10045 76789 10057 76792
rect 10091 76789 10103 76823
rect 10045 76783 10103 76789
rect 1104 76730 10856 76752
rect 1104 76678 2582 76730
rect 2634 76678 2646 76730
rect 2698 76678 2710 76730
rect 2762 76678 2774 76730
rect 2826 76678 2838 76730
rect 2890 76678 5846 76730
rect 5898 76678 5910 76730
rect 5962 76678 5974 76730
rect 6026 76678 6038 76730
rect 6090 76678 6102 76730
rect 6154 76678 9110 76730
rect 9162 76678 9174 76730
rect 9226 76678 9238 76730
rect 9290 76678 9302 76730
rect 9354 76678 9366 76730
rect 9418 76678 10856 76730
rect 1104 76656 10856 76678
rect 2777 76551 2835 76557
rect 2777 76517 2789 76551
rect 2823 76548 2835 76551
rect 3050 76548 3056 76560
rect 2823 76520 3056 76548
rect 2823 76517 2835 76520
rect 2777 76511 2835 76517
rect 3050 76508 3056 76520
rect 3108 76508 3114 76560
rect 9953 76551 10011 76557
rect 9953 76517 9965 76551
rect 9999 76517 10011 76551
rect 9953 76511 10011 76517
rect 9968 76480 9996 76511
rect 2240 76452 9996 76480
rect 1394 76372 1400 76424
rect 1452 76412 1458 76424
rect 2240 76421 2268 76452
rect 1581 76415 1639 76421
rect 1581 76412 1593 76415
rect 1452 76384 1593 76412
rect 1452 76372 1458 76384
rect 1581 76381 1593 76384
rect 1627 76381 1639 76415
rect 1581 76375 1639 76381
rect 2225 76415 2283 76421
rect 2225 76381 2237 76415
rect 2271 76381 2283 76415
rect 2225 76375 2283 76381
rect 2645 76415 2703 76421
rect 2645 76381 2657 76415
rect 2691 76412 2703 76415
rect 2774 76412 2780 76424
rect 2691 76384 2780 76412
rect 2691 76381 2703 76384
rect 2645 76375 2703 76381
rect 2774 76372 2780 76384
rect 2832 76372 2838 76424
rect 3970 76412 3976 76424
rect 3931 76384 3976 76412
rect 3970 76372 3976 76384
rect 4028 76372 4034 76424
rect 10134 76412 10140 76424
rect 10095 76384 10140 76412
rect 10134 76372 10140 76384
rect 10192 76372 10198 76424
rect 2409 76347 2467 76353
rect 2409 76313 2421 76347
rect 2455 76313 2467 76347
rect 2409 76307 2467 76313
rect 2501 76347 2559 76353
rect 2501 76313 2513 76347
rect 2547 76344 2559 76347
rect 3234 76344 3240 76356
rect 2547 76316 3240 76344
rect 2547 76313 2559 76316
rect 2501 76307 2559 76313
rect 1397 76279 1455 76285
rect 1397 76245 1409 76279
rect 1443 76276 1455 76279
rect 1670 76276 1676 76288
rect 1443 76248 1676 76276
rect 1443 76245 1455 76248
rect 1397 76239 1455 76245
rect 1670 76236 1676 76248
rect 1728 76236 1734 76288
rect 2424 76276 2452 76307
rect 3234 76304 3240 76316
rect 3292 76304 3298 76356
rect 2590 76276 2596 76288
rect 2424 76248 2596 76276
rect 2590 76236 2596 76248
rect 2648 76236 2654 76288
rect 3786 76276 3792 76288
rect 3747 76248 3792 76276
rect 3786 76236 3792 76248
rect 3844 76236 3850 76288
rect 1104 76186 10856 76208
rect 1104 76134 4214 76186
rect 4266 76134 4278 76186
rect 4330 76134 4342 76186
rect 4394 76134 4406 76186
rect 4458 76134 4470 76186
rect 4522 76134 7478 76186
rect 7530 76134 7542 76186
rect 7594 76134 7606 76186
rect 7658 76134 7670 76186
rect 7722 76134 7734 76186
rect 7786 76134 10856 76186
rect 1104 76112 10856 76134
rect 1397 76075 1455 76081
rect 1397 76041 1409 76075
rect 1443 76072 1455 76075
rect 1762 76072 1768 76084
rect 1443 76044 1768 76072
rect 1443 76041 1455 76044
rect 1397 76035 1455 76041
rect 1762 76032 1768 76044
rect 1820 76032 1826 76084
rect 9953 76075 10011 76081
rect 9953 76072 9965 76075
rect 2746 76044 9965 76072
rect 2746 76004 2774 76044
rect 9953 76041 9965 76044
rect 9999 76041 10011 76075
rect 9953 76035 10011 76041
rect 2424 75976 2774 76004
rect 2978 76007 3036 76013
rect 1578 75936 1584 75948
rect 1539 75908 1584 75936
rect 1578 75896 1584 75908
rect 1636 75896 1642 75948
rect 2424 75945 2452 75976
rect 2978 75973 2990 76007
rect 3024 76004 3036 76007
rect 5258 76004 5264 76016
rect 3024 75976 5264 76004
rect 3024 75973 3036 75976
rect 2978 75967 3036 75973
rect 5258 75964 5264 75976
rect 5316 75964 5322 76016
rect 2409 75939 2467 75945
rect 2409 75905 2421 75939
rect 2455 75905 2467 75939
rect 2590 75936 2596 75948
rect 2503 75908 2596 75936
rect 2409 75899 2467 75905
rect 2590 75896 2596 75908
rect 2648 75896 2654 75948
rect 2685 75939 2743 75945
rect 2685 75905 2697 75939
rect 2731 75905 2743 75939
rect 2685 75899 2743 75905
rect 2038 75828 2044 75880
rect 2096 75868 2102 75880
rect 2608 75868 2636 75896
rect 2096 75840 2636 75868
rect 2700 75868 2728 75899
rect 2774 75896 2780 75948
rect 2832 75945 2838 75948
rect 2832 75936 2840 75945
rect 3142 75936 3148 75948
rect 2832 75908 2877 75936
rect 2976 75908 3148 75936
rect 2832 75899 2840 75908
rect 2832 75896 2838 75899
rect 2976 75868 3004 75908
rect 3142 75896 3148 75908
rect 3200 75896 3206 75948
rect 3694 75936 3700 75948
rect 3655 75908 3700 75936
rect 3694 75896 3700 75908
rect 3752 75896 3758 75948
rect 10134 75936 10140 75948
rect 10095 75908 10140 75936
rect 10134 75896 10140 75908
rect 10192 75896 10198 75948
rect 2700 75840 3004 75868
rect 2096 75828 2102 75840
rect 2314 75760 2320 75812
rect 2372 75800 2378 75812
rect 2774 75800 2780 75812
rect 2372 75772 2780 75800
rect 2372 75760 2378 75772
rect 2774 75760 2780 75772
rect 2832 75760 2838 75812
rect 3510 75732 3516 75744
rect 3471 75704 3516 75732
rect 3510 75692 3516 75704
rect 3568 75692 3574 75744
rect 1104 75642 10856 75664
rect 1104 75590 2582 75642
rect 2634 75590 2646 75642
rect 2698 75590 2710 75642
rect 2762 75590 2774 75642
rect 2826 75590 2838 75642
rect 2890 75590 5846 75642
rect 5898 75590 5910 75642
rect 5962 75590 5974 75642
rect 6026 75590 6038 75642
rect 6090 75590 6102 75642
rect 6154 75590 9110 75642
rect 9162 75590 9174 75642
rect 9226 75590 9238 75642
rect 9290 75590 9302 75642
rect 9354 75590 9366 75642
rect 9418 75590 10856 75642
rect 1104 75568 10856 75590
rect 2498 75460 2504 75472
rect 2459 75432 2504 75460
rect 2498 75420 2504 75432
rect 2556 75420 2562 75472
rect 9953 75463 10011 75469
rect 9953 75460 9965 75463
rect 2746 75432 9965 75460
rect 2746 75392 2774 75432
rect 9953 75429 9965 75432
rect 9999 75429 10011 75463
rect 9953 75423 10011 75429
rect 1964 75364 2774 75392
rect 1964 75333 1992 75364
rect 1949 75327 2007 75333
rect 1949 75293 1961 75327
rect 1995 75293 2007 75327
rect 2314 75324 2320 75336
rect 2372 75333 2378 75336
rect 1949 75287 2007 75293
rect 2056 75296 2320 75324
rect 1854 75216 1860 75268
rect 1912 75256 1918 75268
rect 2056 75256 2084 75296
rect 2314 75284 2320 75296
rect 2372 75287 2380 75333
rect 10134 75324 10140 75336
rect 10095 75296 10140 75324
rect 2372 75284 2378 75287
rect 10134 75284 10140 75296
rect 10192 75284 10198 75336
rect 1912 75228 2084 75256
rect 2133 75259 2191 75265
rect 1912 75216 1918 75228
rect 2133 75225 2145 75259
rect 2179 75225 2191 75259
rect 2133 75219 2191 75225
rect 2225 75259 2283 75265
rect 2225 75225 2237 75259
rect 2271 75256 2283 75259
rect 2958 75256 2964 75268
rect 2271 75228 2964 75256
rect 2271 75225 2283 75228
rect 2225 75219 2283 75225
rect 1486 75148 1492 75200
rect 1544 75188 1550 75200
rect 2038 75188 2044 75200
rect 1544 75160 2044 75188
rect 1544 75148 1550 75160
rect 2038 75148 2044 75160
rect 2096 75188 2102 75200
rect 2148 75188 2176 75219
rect 2958 75216 2964 75228
rect 3016 75216 3022 75268
rect 2096 75160 2176 75188
rect 2096 75148 2102 75160
rect 1104 75098 10856 75120
rect 1104 75046 4214 75098
rect 4266 75046 4278 75098
rect 4330 75046 4342 75098
rect 4394 75046 4406 75098
rect 4458 75046 4470 75098
rect 4522 75046 7478 75098
rect 7530 75046 7542 75098
rect 7594 75046 7606 75098
rect 7658 75046 7670 75098
rect 7722 75046 7734 75098
rect 7786 75046 10856 75098
rect 1104 75024 10856 75046
rect 1673 74919 1731 74925
rect 1673 74885 1685 74919
rect 1719 74916 1731 74919
rect 3878 74916 3884 74928
rect 1719 74888 3884 74916
rect 1719 74885 1731 74888
rect 1673 74879 1731 74885
rect 3878 74876 3884 74888
rect 3936 74876 3942 74928
rect 1397 74851 1455 74857
rect 1397 74817 1409 74851
rect 1443 74817 1455 74851
rect 1397 74811 1455 74817
rect 1412 74780 1440 74811
rect 1486 74808 1492 74860
rect 1544 74848 1550 74860
rect 1854 74857 1860 74860
rect 1581 74851 1639 74857
rect 1581 74848 1593 74851
rect 1544 74820 1593 74848
rect 1544 74808 1550 74820
rect 1581 74817 1593 74820
rect 1627 74817 1639 74851
rect 1581 74811 1639 74817
rect 1817 74851 1860 74857
rect 1817 74817 1829 74851
rect 1817 74811 1860 74817
rect 1854 74808 1860 74811
rect 1912 74808 1918 74860
rect 2685 74851 2743 74857
rect 2685 74817 2697 74851
rect 2731 74848 2743 74851
rect 2958 74848 2964 74860
rect 2731 74820 2964 74848
rect 2731 74817 2743 74820
rect 2685 74811 2743 74817
rect 2958 74808 2964 74820
rect 3016 74808 3022 74860
rect 8294 74780 8300 74792
rect 1412 74752 8300 74780
rect 8294 74740 8300 74752
rect 8352 74740 8358 74792
rect 2038 74672 2044 74724
rect 2096 74712 2102 74724
rect 2501 74715 2559 74721
rect 2501 74712 2513 74715
rect 2096 74684 2513 74712
rect 2096 74672 2102 74684
rect 2501 74681 2513 74684
rect 2547 74681 2559 74715
rect 2501 74675 2559 74681
rect 1949 74647 2007 74653
rect 1949 74613 1961 74647
rect 1995 74644 2007 74647
rect 2314 74644 2320 74656
rect 1995 74616 2320 74644
rect 1995 74613 2007 74616
rect 1949 74607 2007 74613
rect 2314 74604 2320 74616
rect 2372 74604 2378 74656
rect 1104 74554 10856 74576
rect 1104 74502 2582 74554
rect 2634 74502 2646 74554
rect 2698 74502 2710 74554
rect 2762 74502 2774 74554
rect 2826 74502 2838 74554
rect 2890 74502 5846 74554
rect 5898 74502 5910 74554
rect 5962 74502 5974 74554
rect 6026 74502 6038 74554
rect 6090 74502 6102 74554
rect 6154 74502 9110 74554
rect 9162 74502 9174 74554
rect 9226 74502 9238 74554
rect 9290 74502 9302 74554
rect 9354 74502 9366 74554
rect 9418 74502 10856 74554
rect 1104 74480 10856 74502
rect 934 74332 940 74384
rect 992 74372 998 74384
rect 2501 74375 2559 74381
rect 2501 74372 2513 74375
rect 992 74344 2513 74372
rect 992 74332 998 74344
rect 2501 74341 2513 74344
rect 2547 74341 2559 74375
rect 9953 74375 10011 74381
rect 9953 74372 9965 74375
rect 2501 74335 2559 74341
rect 2746 74344 9965 74372
rect 2746 74304 2774 74344
rect 9953 74341 9965 74344
rect 9999 74341 10011 74375
rect 9953 74335 10011 74341
rect 1964 74276 2774 74304
rect 1964 74245 1992 74276
rect 1949 74239 2007 74245
rect 1949 74205 1961 74239
rect 1995 74205 2007 74239
rect 2322 74239 2380 74245
rect 2322 74236 2334 74239
rect 1949 74199 2007 74205
rect 2056 74208 2334 74236
rect 1854 74128 1860 74180
rect 1912 74168 1918 74180
rect 2056 74168 2084 74208
rect 2322 74205 2334 74208
rect 2368 74205 2380 74239
rect 10134 74236 10140 74248
rect 10095 74208 10140 74236
rect 2322 74199 2380 74205
rect 10134 74196 10140 74208
rect 10192 74196 10198 74248
rect 1912 74140 2084 74168
rect 2133 74171 2191 74177
rect 1912 74128 1918 74140
rect 2133 74137 2145 74171
rect 2179 74137 2191 74171
rect 2133 74131 2191 74137
rect 2225 74171 2283 74177
rect 2225 74137 2237 74171
rect 2271 74168 2283 74171
rect 3602 74168 3608 74180
rect 2271 74140 3608 74168
rect 2271 74137 2283 74140
rect 2225 74131 2283 74137
rect 1118 74060 1124 74112
rect 1176 74100 1182 74112
rect 1486 74100 1492 74112
rect 1176 74072 1492 74100
rect 1176 74060 1182 74072
rect 1486 74060 1492 74072
rect 1544 74100 1550 74112
rect 2148 74100 2176 74131
rect 3602 74128 3608 74140
rect 3660 74128 3666 74180
rect 1544 74072 2176 74100
rect 1544 74060 1550 74072
rect 1104 74010 10856 74032
rect 1104 73958 4214 74010
rect 4266 73958 4278 74010
rect 4330 73958 4342 74010
rect 4394 73958 4406 74010
rect 4458 73958 4470 74010
rect 4522 73958 7478 74010
rect 7530 73958 7542 74010
rect 7594 73958 7606 74010
rect 7658 73958 7670 74010
rect 7722 73958 7734 74010
rect 7786 73958 10856 74010
rect 1104 73936 10856 73958
rect 1394 73720 1400 73772
rect 1452 73760 1458 73772
rect 1581 73763 1639 73769
rect 1581 73760 1593 73763
rect 1452 73732 1593 73760
rect 1452 73720 1458 73732
rect 1581 73729 1593 73732
rect 1627 73729 1639 73763
rect 2222 73760 2228 73772
rect 2183 73732 2228 73760
rect 1581 73723 1639 73729
rect 2222 73720 2228 73732
rect 2280 73720 2286 73772
rect 2866 73760 2872 73772
rect 2827 73732 2872 73760
rect 2866 73720 2872 73732
rect 2924 73720 2930 73772
rect 10134 73760 10140 73772
rect 10095 73732 10140 73760
rect 10134 73720 10140 73732
rect 10192 73720 10198 73772
rect 1302 73516 1308 73568
rect 1360 73556 1366 73568
rect 1397 73559 1455 73565
rect 1397 73556 1409 73559
rect 1360 73528 1409 73556
rect 1360 73516 1366 73528
rect 1397 73525 1409 73528
rect 1443 73525 1455 73559
rect 1397 73519 1455 73525
rect 1486 73516 1492 73568
rect 1544 73556 1550 73568
rect 2041 73559 2099 73565
rect 2041 73556 2053 73559
rect 1544 73528 2053 73556
rect 1544 73516 1550 73528
rect 2041 73525 2053 73528
rect 2087 73525 2099 73559
rect 2041 73519 2099 73525
rect 2685 73559 2743 73565
rect 2685 73525 2697 73559
rect 2731 73556 2743 73559
rect 3142 73556 3148 73568
rect 2731 73528 3148 73556
rect 2731 73525 2743 73528
rect 2685 73519 2743 73525
rect 3142 73516 3148 73528
rect 3200 73516 3206 73568
rect 8294 73516 8300 73568
rect 8352 73556 8358 73568
rect 9953 73559 10011 73565
rect 9953 73556 9965 73559
rect 8352 73528 9965 73556
rect 8352 73516 8358 73528
rect 9953 73525 9965 73528
rect 9999 73525 10011 73559
rect 9953 73519 10011 73525
rect 1104 73466 10856 73488
rect 1104 73414 2582 73466
rect 2634 73414 2646 73466
rect 2698 73414 2710 73466
rect 2762 73414 2774 73466
rect 2826 73414 2838 73466
rect 2890 73414 5846 73466
rect 5898 73414 5910 73466
rect 5962 73414 5974 73466
rect 6026 73414 6038 73466
rect 6090 73414 6102 73466
rect 6154 73414 9110 73466
rect 9162 73414 9174 73466
rect 9226 73414 9238 73466
rect 9290 73414 9302 73466
rect 9354 73414 9366 73466
rect 9418 73414 10856 73466
rect 1104 73392 10856 73414
rect 2314 73176 2320 73228
rect 2372 73216 2378 73228
rect 3326 73216 3332 73228
rect 2372 73188 3332 73216
rect 2372 73176 2378 73188
rect 3326 73176 3332 73188
rect 3384 73176 3390 73228
rect 1578 73148 1584 73160
rect 1539 73120 1584 73148
rect 1578 73108 1584 73120
rect 1636 73108 1642 73160
rect 2774 73040 2780 73092
rect 2832 73080 2838 73092
rect 3786 73080 3792 73092
rect 2832 73052 3792 73080
rect 2832 73040 2838 73052
rect 3786 73040 3792 73052
rect 3844 73040 3850 73092
rect 1210 72972 1216 73024
rect 1268 73012 1274 73024
rect 1397 73015 1455 73021
rect 1397 73012 1409 73015
rect 1268 72984 1409 73012
rect 1268 72972 1274 72984
rect 1397 72981 1409 72984
rect 1443 72981 1455 73015
rect 1397 72975 1455 72981
rect 1104 72922 10856 72944
rect 1104 72870 4214 72922
rect 4266 72870 4278 72922
rect 4330 72870 4342 72922
rect 4394 72870 4406 72922
rect 4458 72870 4470 72922
rect 4522 72870 7478 72922
rect 7530 72870 7542 72922
rect 7594 72870 7606 72922
rect 7658 72870 7670 72922
rect 7722 72870 7734 72922
rect 7786 72870 10856 72922
rect 1104 72848 10856 72870
rect 3510 72808 3516 72820
rect 1688 72780 3516 72808
rect 1118 72700 1124 72752
rect 1176 72740 1182 72752
rect 1688 72749 1716 72780
rect 3510 72768 3516 72780
rect 3568 72768 3574 72820
rect 1581 72743 1639 72749
rect 1581 72740 1593 72743
rect 1176 72712 1593 72740
rect 1176 72700 1182 72712
rect 1581 72709 1593 72712
rect 1627 72709 1639 72743
rect 1581 72703 1639 72709
rect 1673 72743 1731 72749
rect 1673 72709 1685 72743
rect 1719 72709 1731 72743
rect 8294 72740 8300 72752
rect 1673 72703 1731 72709
rect 2516 72712 8300 72740
rect 1854 72681 1860 72684
rect 1397 72675 1455 72681
rect 1397 72641 1409 72675
rect 1443 72641 1455 72675
rect 1397 72635 1455 72641
rect 1817 72675 1860 72681
rect 1817 72641 1829 72675
rect 1817 72635 1860 72641
rect 1412 72604 1440 72635
rect 1854 72632 1860 72635
rect 1912 72632 1918 72684
rect 2516 72681 2544 72712
rect 8294 72700 8300 72712
rect 8352 72700 8358 72752
rect 2501 72675 2559 72681
rect 2501 72641 2513 72675
rect 2547 72641 2559 72675
rect 2682 72672 2688 72684
rect 2643 72644 2688 72672
rect 2501 72635 2559 72641
rect 2682 72632 2688 72644
rect 2740 72632 2746 72684
rect 2774 72632 2780 72684
rect 2832 72672 2838 72684
rect 2958 72681 2964 72684
rect 2921 72675 2964 72681
rect 2832 72644 2877 72672
rect 2832 72632 2838 72644
rect 2921 72641 2933 72675
rect 2921 72635 2964 72641
rect 2958 72632 2964 72635
rect 3016 72632 3022 72684
rect 10134 72672 10140 72684
rect 10095 72644 10140 72672
rect 10134 72632 10140 72644
rect 10192 72632 10198 72684
rect 9950 72604 9956 72616
rect 1412 72576 9956 72604
rect 9950 72564 9956 72576
rect 10008 72564 10014 72616
rect 1949 72539 2007 72545
rect 1949 72505 1961 72539
rect 1995 72536 2007 72539
rect 5534 72536 5540 72548
rect 1995 72508 5540 72536
rect 1995 72505 2007 72508
rect 1949 72499 2007 72505
rect 5534 72496 5540 72508
rect 5592 72496 5598 72548
rect 1854 72428 1860 72480
rect 1912 72468 1918 72480
rect 2958 72468 2964 72480
rect 1912 72440 2964 72468
rect 1912 72428 1918 72440
rect 2958 72428 2964 72440
rect 3016 72428 3022 72480
rect 3053 72471 3111 72477
rect 3053 72437 3065 72471
rect 3099 72468 3111 72471
rect 3878 72468 3884 72480
rect 3099 72440 3884 72468
rect 3099 72437 3111 72440
rect 3053 72431 3111 72437
rect 3878 72428 3884 72440
rect 3936 72428 3942 72480
rect 4614 72428 4620 72480
rect 4672 72468 4678 72480
rect 9953 72471 10011 72477
rect 9953 72468 9965 72471
rect 4672 72440 9965 72468
rect 4672 72428 4678 72440
rect 9953 72437 9965 72440
rect 9999 72437 10011 72471
rect 9953 72431 10011 72437
rect 1104 72378 10856 72400
rect 1104 72326 2582 72378
rect 2634 72326 2646 72378
rect 2698 72326 2710 72378
rect 2762 72326 2774 72378
rect 2826 72326 2838 72378
rect 2890 72326 5846 72378
rect 5898 72326 5910 72378
rect 5962 72326 5974 72378
rect 6026 72326 6038 72378
rect 6090 72326 6102 72378
rect 6154 72326 9110 72378
rect 9162 72326 9174 72378
rect 9226 72326 9238 72378
rect 9290 72326 9302 72378
rect 9354 72326 9366 72378
rect 9418 72326 10856 72378
rect 1104 72304 10856 72326
rect 9950 72264 9956 72276
rect 9911 72236 9956 72264
rect 9950 72224 9956 72236
rect 10008 72224 10014 72276
rect 1854 72156 1860 72208
rect 1912 72196 1918 72208
rect 2685 72199 2743 72205
rect 2685 72196 2697 72199
rect 1912 72168 2697 72196
rect 1912 72156 1918 72168
rect 2685 72165 2697 72168
rect 2731 72165 2743 72199
rect 2685 72159 2743 72165
rect 1578 72060 1584 72072
rect 1539 72032 1584 72060
rect 1578 72020 1584 72032
rect 1636 72020 1642 72072
rect 2222 72060 2228 72072
rect 2183 72032 2228 72060
rect 2222 72020 2228 72032
rect 2280 72020 2286 72072
rect 2866 72060 2872 72072
rect 2827 72032 2872 72060
rect 2866 72020 2872 72032
rect 2924 72020 2930 72072
rect 10134 72060 10140 72072
rect 10095 72032 10140 72060
rect 10134 72020 10140 72032
rect 10192 72020 10198 72072
rect 1026 71884 1032 71936
rect 1084 71924 1090 71936
rect 1397 71927 1455 71933
rect 1397 71924 1409 71927
rect 1084 71896 1409 71924
rect 1084 71884 1090 71896
rect 1397 71893 1409 71896
rect 1443 71893 1455 71927
rect 1397 71887 1455 71893
rect 2041 71927 2099 71933
rect 2041 71893 2053 71927
rect 2087 71924 2099 71927
rect 2314 71924 2320 71936
rect 2087 71896 2320 71924
rect 2087 71893 2099 71896
rect 2041 71887 2099 71893
rect 2314 71884 2320 71896
rect 2372 71884 2378 71936
rect 2590 71884 2596 71936
rect 2648 71924 2654 71936
rect 4614 71924 4620 71936
rect 2648 71896 4620 71924
rect 2648 71884 2654 71896
rect 4614 71884 4620 71896
rect 4672 71884 4678 71936
rect 1104 71834 10856 71856
rect 1104 71782 4214 71834
rect 4266 71782 4278 71834
rect 4330 71782 4342 71834
rect 4394 71782 4406 71834
rect 4458 71782 4470 71834
rect 4522 71782 7478 71834
rect 7530 71782 7542 71834
rect 7594 71782 7606 71834
rect 7658 71782 7670 71834
rect 7722 71782 7734 71834
rect 7786 71782 10856 71834
rect 1104 71760 10856 71782
rect 1504 71692 2084 71720
rect 1118 71612 1124 71664
rect 1176 71652 1182 71664
rect 1504 71652 1532 71692
rect 1670 71652 1676 71664
rect 1176 71624 1532 71652
rect 1631 71624 1676 71652
rect 1176 71612 1182 71624
rect 1397 71587 1455 71593
rect 1397 71553 1409 71587
rect 1443 71553 1455 71587
rect 1504 71584 1532 71624
rect 1670 71612 1676 71624
rect 1728 71612 1734 71664
rect 2056 71652 2084 71692
rect 2406 71680 2412 71732
rect 2464 71720 2470 71732
rect 2464 71692 2820 71720
rect 2464 71680 2470 71692
rect 2792 71661 2820 71692
rect 2685 71655 2743 71661
rect 2685 71652 2697 71655
rect 2056 71624 2697 71652
rect 2685 71621 2697 71624
rect 2731 71621 2743 71655
rect 2685 71615 2743 71621
rect 2777 71655 2835 71661
rect 2777 71621 2789 71655
rect 2823 71621 2835 71655
rect 2777 71615 2835 71621
rect 1581 71587 1639 71593
rect 1581 71584 1593 71587
rect 1504 71556 1593 71584
rect 1397 71547 1455 71553
rect 1581 71553 1593 71556
rect 1627 71553 1639 71587
rect 1581 71547 1639 71553
rect 1817 71587 1875 71593
rect 1817 71553 1829 71587
rect 1863 71584 1875 71587
rect 2406 71584 2412 71596
rect 1863 71556 2412 71584
rect 1863 71553 1875 71556
rect 1817 71547 1875 71553
rect 1412 71516 1440 71547
rect 2406 71544 2412 71556
rect 2464 71544 2470 71596
rect 2501 71587 2559 71593
rect 2501 71553 2513 71587
rect 2547 71584 2559 71587
rect 2590 71584 2596 71596
rect 2547 71556 2596 71584
rect 2547 71553 2559 71556
rect 2501 71547 2559 71553
rect 2590 71544 2596 71556
rect 2648 71544 2654 71596
rect 2958 71593 2964 71596
rect 2921 71587 2964 71593
rect 2921 71553 2933 71587
rect 2921 71547 2964 71553
rect 2958 71544 2964 71547
rect 3016 71544 3022 71596
rect 3070 71587 3128 71593
rect 3070 71553 3082 71587
rect 3116 71584 3128 71587
rect 3694 71584 3700 71596
rect 3116 71556 3700 71584
rect 3116 71553 3128 71556
rect 3070 71547 3128 71553
rect 3694 71544 3700 71556
rect 3752 71544 3758 71596
rect 10134 71584 10140 71596
rect 10095 71556 10140 71584
rect 10134 71544 10140 71556
rect 10192 71544 10198 71596
rect 1412 71488 2176 71516
rect 1670 71408 1676 71460
rect 1728 71448 1734 71460
rect 2038 71448 2044 71460
rect 1728 71420 2044 71448
rect 1728 71408 1734 71420
rect 2038 71408 2044 71420
rect 2096 71408 2102 71460
rect 2148 71448 2176 71488
rect 2936 71488 9996 71516
rect 2936 71448 2964 71488
rect 5626 71448 5632 71460
rect 2148 71420 2964 71448
rect 3068 71420 5632 71448
rect 1949 71383 2007 71389
rect 1949 71349 1961 71383
rect 1995 71380 2007 71383
rect 3068 71380 3096 71420
rect 5626 71408 5632 71420
rect 5684 71408 5690 71460
rect 9968 71457 9996 71488
rect 9953 71451 10011 71457
rect 9953 71417 9965 71451
rect 9999 71417 10011 71451
rect 9953 71411 10011 71417
rect 1995 71352 3096 71380
rect 1995 71349 2007 71352
rect 1949 71343 2007 71349
rect 1104 71290 10856 71312
rect 1104 71238 2582 71290
rect 2634 71238 2646 71290
rect 2698 71238 2710 71290
rect 2762 71238 2774 71290
rect 2826 71238 2838 71290
rect 2890 71238 5846 71290
rect 5898 71238 5910 71290
rect 5962 71238 5974 71290
rect 6026 71238 6038 71290
rect 6090 71238 6102 71290
rect 6154 71238 9110 71290
rect 9162 71238 9174 71290
rect 9226 71238 9238 71290
rect 9290 71238 9302 71290
rect 9354 71238 9366 71290
rect 9418 71238 10856 71290
rect 1104 71216 10856 71238
rect 1578 70972 1584 70984
rect 1539 70944 1584 70972
rect 1578 70932 1584 70944
rect 1636 70932 1642 70984
rect 1397 70839 1455 70845
rect 1397 70805 1409 70839
rect 1443 70836 1455 70839
rect 1486 70836 1492 70848
rect 1443 70808 1492 70836
rect 1443 70805 1455 70808
rect 1397 70799 1455 70805
rect 1486 70796 1492 70808
rect 1544 70796 1550 70848
rect 1104 70746 10856 70768
rect 1104 70694 4214 70746
rect 4266 70694 4278 70746
rect 4330 70694 4342 70746
rect 4394 70694 4406 70746
rect 4458 70694 4470 70746
rect 4522 70694 7478 70746
rect 7530 70694 7542 70746
rect 7594 70694 7606 70746
rect 7658 70694 7670 70746
rect 7722 70694 7734 70746
rect 7786 70694 10856 70746
rect 1104 70672 10856 70694
rect 1762 70592 1768 70644
rect 1820 70592 1826 70644
rect 1966 70635 2024 70641
rect 1966 70601 1978 70635
rect 2012 70632 2024 70635
rect 3510 70632 3516 70644
rect 2012 70604 3516 70632
rect 2012 70601 2024 70604
rect 1966 70595 2024 70601
rect 3510 70592 3516 70604
rect 3568 70592 3574 70644
rect 1118 70524 1124 70576
rect 1176 70564 1182 70576
rect 1581 70567 1639 70573
rect 1581 70564 1593 70567
rect 1176 70536 1593 70564
rect 1176 70524 1182 70536
rect 1581 70533 1593 70536
rect 1627 70533 1639 70567
rect 1581 70527 1639 70533
rect 1673 70567 1731 70573
rect 1673 70533 1685 70567
rect 1719 70564 1731 70567
rect 1780 70564 1808 70592
rect 2406 70564 2412 70576
rect 1719 70536 1808 70564
rect 1981 70536 2412 70564
rect 1719 70533 1731 70536
rect 1673 70527 1731 70533
rect 1397 70499 1455 70505
rect 1397 70465 1409 70499
rect 1443 70465 1455 70499
rect 1397 70459 1455 70465
rect 1817 70499 1875 70505
rect 1817 70465 1829 70499
rect 1863 70496 1875 70499
rect 1981 70496 2009 70536
rect 2406 70524 2412 70536
rect 2464 70564 2470 70576
rect 2958 70564 2964 70576
rect 2464 70536 2964 70564
rect 2464 70524 2470 70536
rect 2958 70524 2964 70536
rect 3016 70524 3022 70576
rect 1863 70468 2009 70496
rect 1863 70465 1875 70468
rect 1817 70459 1875 70465
rect 1412 70428 1440 70459
rect 2038 70456 2044 70508
rect 2096 70496 2102 70508
rect 2685 70499 2743 70505
rect 2685 70496 2697 70499
rect 2096 70468 2697 70496
rect 2096 70456 2102 70468
rect 2685 70465 2697 70468
rect 2731 70465 2743 70499
rect 10134 70496 10140 70508
rect 10095 70468 10140 70496
rect 2685 70459 2743 70465
rect 10134 70456 10140 70468
rect 10192 70456 10198 70508
rect 1412 70400 9996 70428
rect 9968 70369 9996 70400
rect 9953 70363 10011 70369
rect 9953 70329 9965 70363
rect 9999 70360 10011 70363
rect 9999 70332 10033 70360
rect 9999 70329 10011 70332
rect 9953 70323 10011 70329
rect 1486 70252 1492 70304
rect 1544 70292 1550 70304
rect 1854 70292 1860 70304
rect 1544 70264 1860 70292
rect 1544 70252 1550 70264
rect 1854 70252 1860 70264
rect 1912 70252 1918 70304
rect 2406 70252 2412 70304
rect 2464 70292 2470 70304
rect 2501 70295 2559 70301
rect 2501 70292 2513 70295
rect 2464 70264 2513 70292
rect 2464 70252 2470 70264
rect 2501 70261 2513 70264
rect 2547 70261 2559 70295
rect 2501 70255 2559 70261
rect 1104 70202 10856 70224
rect 1104 70150 2582 70202
rect 2634 70150 2646 70202
rect 2698 70150 2710 70202
rect 2762 70150 2774 70202
rect 2826 70150 2838 70202
rect 2890 70150 5846 70202
rect 5898 70150 5910 70202
rect 5962 70150 5974 70202
rect 6026 70150 6038 70202
rect 6090 70150 6102 70202
rect 6154 70150 9110 70202
rect 9162 70150 9174 70202
rect 9226 70150 9238 70202
rect 9290 70150 9302 70202
rect 9354 70150 9366 70202
rect 9418 70150 10856 70202
rect 1104 70128 10856 70150
rect 1578 69884 1584 69896
rect 1539 69856 1584 69884
rect 1578 69844 1584 69856
rect 1636 69844 1642 69896
rect 2222 69884 2228 69896
rect 2183 69856 2228 69884
rect 2222 69844 2228 69856
rect 2280 69844 2286 69896
rect 2866 69884 2872 69896
rect 2827 69856 2872 69884
rect 2866 69844 2872 69856
rect 2924 69844 2930 69896
rect 10134 69884 10140 69896
rect 10095 69856 10140 69884
rect 10134 69844 10140 69856
rect 10192 69844 10198 69896
rect 1302 69776 1308 69828
rect 1360 69816 1366 69828
rect 1360 69788 1624 69816
rect 1360 69776 1366 69788
rect 1596 69760 1624 69788
rect 750 69708 756 69760
rect 808 69748 814 69760
rect 1397 69751 1455 69757
rect 1397 69748 1409 69751
rect 808 69720 1409 69748
rect 808 69708 814 69720
rect 1397 69717 1409 69720
rect 1443 69717 1455 69751
rect 1397 69711 1455 69717
rect 1578 69708 1584 69760
rect 1636 69708 1642 69760
rect 2038 69748 2044 69760
rect 1999 69720 2044 69748
rect 2038 69708 2044 69720
rect 2096 69708 2102 69760
rect 2682 69748 2688 69760
rect 2643 69720 2688 69748
rect 2682 69708 2688 69720
rect 2740 69708 2746 69760
rect 3050 69708 3056 69760
rect 3108 69748 3114 69760
rect 3786 69748 3792 69760
rect 3108 69720 3792 69748
rect 3108 69708 3114 69720
rect 3786 69708 3792 69720
rect 3844 69708 3850 69760
rect 9950 69748 9956 69760
rect 9911 69720 9956 69748
rect 9950 69708 9956 69720
rect 10008 69708 10014 69760
rect 1104 69658 10856 69680
rect 1104 69606 4214 69658
rect 4266 69606 4278 69658
rect 4330 69606 4342 69658
rect 4394 69606 4406 69658
rect 4458 69606 4470 69658
rect 4522 69606 7478 69658
rect 7530 69606 7542 69658
rect 7594 69606 7606 69658
rect 7658 69606 7670 69658
rect 7722 69606 7734 69658
rect 7786 69606 10856 69658
rect 1104 69584 10856 69606
rect 1118 69436 1124 69488
rect 1176 69476 1182 69488
rect 1670 69476 1676 69488
rect 1176 69448 1532 69476
rect 1631 69448 1676 69476
rect 1176 69436 1182 69448
rect 1504 69420 1532 69448
rect 1670 69436 1676 69448
rect 1728 69436 1734 69488
rect 3050 69476 3056 69488
rect 1832 69448 3056 69476
rect 1397 69411 1455 69417
rect 1397 69377 1409 69411
rect 1443 69377 1455 69411
rect 1397 69371 1455 69377
rect 1412 69340 1440 69371
rect 1486 69368 1492 69420
rect 1544 69408 1550 69420
rect 1832 69417 1860 69448
rect 3050 69436 3056 69448
rect 3108 69436 3114 69488
rect 1581 69411 1639 69417
rect 1581 69408 1593 69411
rect 1544 69380 1593 69408
rect 1544 69368 1550 69380
rect 1581 69377 1593 69380
rect 1627 69377 1639 69411
rect 1581 69371 1639 69377
rect 1817 69411 1875 69417
rect 1817 69377 1829 69411
rect 1863 69377 1875 69411
rect 1817 69371 1875 69377
rect 2685 69411 2743 69417
rect 2685 69377 2697 69411
rect 2731 69408 2743 69411
rect 2958 69408 2964 69420
rect 2731 69380 2964 69408
rect 2731 69377 2743 69380
rect 2685 69371 2743 69377
rect 2958 69368 2964 69380
rect 3016 69368 3022 69420
rect 9950 69340 9956 69352
rect 1412 69312 9956 69340
rect 9950 69300 9956 69312
rect 10008 69300 10014 69352
rect 1949 69275 2007 69281
rect 1949 69241 1961 69275
rect 1995 69272 2007 69275
rect 5718 69272 5724 69284
rect 1995 69244 5724 69272
rect 1995 69241 2007 69244
rect 1949 69235 2007 69241
rect 5718 69232 5724 69244
rect 5776 69232 5782 69284
rect 1118 69164 1124 69216
rect 1176 69204 1182 69216
rect 2501 69207 2559 69213
rect 2501 69204 2513 69207
rect 1176 69176 2513 69204
rect 1176 69164 1182 69176
rect 2501 69173 2513 69176
rect 2547 69173 2559 69207
rect 2501 69167 2559 69173
rect 1104 69114 10856 69136
rect 1104 69062 2582 69114
rect 2634 69062 2646 69114
rect 2698 69062 2710 69114
rect 2762 69062 2774 69114
rect 2826 69062 2838 69114
rect 2890 69062 5846 69114
rect 5898 69062 5910 69114
rect 5962 69062 5974 69114
rect 6026 69062 6038 69114
rect 6090 69062 6102 69114
rect 6154 69062 9110 69114
rect 9162 69062 9174 69114
rect 9226 69062 9238 69114
rect 9290 69062 9302 69114
rect 9354 69062 9366 69114
rect 9418 69062 10856 69114
rect 1104 69040 10856 69062
rect 9953 69003 10011 69009
rect 9953 69000 9965 69003
rect 2332 68972 9965 69000
rect 1578 68796 1584 68808
rect 1539 68768 1584 68796
rect 1578 68756 1584 68768
rect 1636 68756 1642 68808
rect 2332 68805 2360 68972
rect 9953 68969 9965 68972
rect 9999 68969 10011 69003
rect 9953 68963 10011 68969
rect 2869 68935 2927 68941
rect 2869 68901 2881 68935
rect 2915 68932 2927 68935
rect 4062 68932 4068 68944
rect 2915 68904 4068 68932
rect 2915 68901 2927 68904
rect 2869 68895 2927 68901
rect 4062 68892 4068 68904
rect 4120 68892 4126 68944
rect 2317 68799 2375 68805
rect 2317 68765 2329 68799
rect 2363 68765 2375 68799
rect 2317 68759 2375 68765
rect 2737 68799 2795 68805
rect 2737 68765 2749 68799
rect 2783 68796 2795 68799
rect 2866 68796 2872 68808
rect 2783 68768 2872 68796
rect 2783 68765 2795 68768
rect 2737 68759 2795 68765
rect 2866 68756 2872 68768
rect 2924 68796 2930 68808
rect 3050 68796 3056 68808
rect 2924 68768 3056 68796
rect 2924 68756 2930 68768
rect 3050 68756 3056 68768
rect 3108 68756 3114 68808
rect 10134 68796 10140 68808
rect 10095 68768 10140 68796
rect 10134 68756 10140 68768
rect 10192 68756 10198 68808
rect 1486 68688 1492 68740
rect 1544 68728 1550 68740
rect 2498 68728 2504 68740
rect 1544 68700 2504 68728
rect 1544 68688 1550 68700
rect 2498 68688 2504 68700
rect 2556 68688 2562 68740
rect 2593 68731 2651 68737
rect 2593 68697 2605 68731
rect 2639 68728 2651 68731
rect 3142 68728 3148 68740
rect 2639 68700 3148 68728
rect 2639 68697 2651 68700
rect 2593 68691 2651 68697
rect 3142 68688 3148 68700
rect 3200 68688 3206 68740
rect 1397 68663 1455 68669
rect 1397 68629 1409 68663
rect 1443 68660 1455 68663
rect 2222 68660 2228 68672
rect 1443 68632 2228 68660
rect 1443 68629 1455 68632
rect 1397 68623 1455 68629
rect 2222 68620 2228 68632
rect 2280 68620 2286 68672
rect 1104 68570 10856 68592
rect 1104 68518 4214 68570
rect 4266 68518 4278 68570
rect 4330 68518 4342 68570
rect 4394 68518 4406 68570
rect 4458 68518 4470 68570
rect 4522 68518 7478 68570
rect 7530 68518 7542 68570
rect 7594 68518 7606 68570
rect 7658 68518 7670 68570
rect 7722 68518 7734 68570
rect 7786 68518 10856 68570
rect 1104 68496 10856 68518
rect 658 68280 664 68332
rect 716 68320 722 68332
rect 1673 68323 1731 68329
rect 1673 68320 1685 68323
rect 716 68292 1685 68320
rect 716 68280 722 68292
rect 1673 68289 1685 68292
rect 1719 68289 1731 68323
rect 10134 68320 10140 68332
rect 10095 68292 10140 68320
rect 1673 68283 1731 68289
rect 10134 68280 10140 68292
rect 10192 68280 10198 68332
rect 1302 68212 1308 68264
rect 1360 68252 1366 68264
rect 1397 68255 1455 68261
rect 1397 68252 1409 68255
rect 1360 68224 1409 68252
rect 1360 68212 1366 68224
rect 1397 68221 1409 68224
rect 1443 68221 1455 68255
rect 1397 68215 1455 68221
rect 8294 68076 8300 68128
rect 8352 68116 8358 68128
rect 9953 68119 10011 68125
rect 9953 68116 9965 68119
rect 8352 68088 9965 68116
rect 8352 68076 8358 68088
rect 9953 68085 9965 68088
rect 9999 68085 10011 68119
rect 9953 68079 10011 68085
rect 1104 68026 10856 68048
rect 1104 67974 2582 68026
rect 2634 67974 2646 68026
rect 2698 67974 2710 68026
rect 2762 67974 2774 68026
rect 2826 67974 2838 68026
rect 2890 67974 5846 68026
rect 5898 67974 5910 68026
rect 5962 67974 5974 68026
rect 6026 67974 6038 68026
rect 6090 67974 6102 68026
rect 6154 67974 9110 68026
rect 9162 67974 9174 68026
rect 9226 67974 9238 68026
rect 9290 67974 9302 68026
rect 9354 67974 9366 68026
rect 9418 67974 10856 68026
rect 1104 67952 10856 67974
rect 1394 67708 1400 67720
rect 1355 67680 1400 67708
rect 1394 67668 1400 67680
rect 1452 67668 1458 67720
rect 1670 67708 1676 67720
rect 1631 67680 1676 67708
rect 1670 67668 1676 67680
rect 1728 67668 1734 67720
rect 3510 67600 3516 67652
rect 3568 67640 3574 67652
rect 4798 67640 4804 67652
rect 3568 67612 4804 67640
rect 3568 67600 3574 67612
rect 4798 67600 4804 67612
rect 4856 67600 4862 67652
rect 1104 67482 10856 67504
rect 1104 67430 4214 67482
rect 4266 67430 4278 67482
rect 4330 67430 4342 67482
rect 4394 67430 4406 67482
rect 4458 67430 4470 67482
rect 4522 67430 7478 67482
rect 7530 67430 7542 67482
rect 7594 67430 7606 67482
rect 7658 67430 7670 67482
rect 7722 67430 7734 67482
rect 7786 67430 10856 67482
rect 1104 67408 10856 67430
rect 2222 67260 2228 67312
rect 2280 67300 2286 67312
rect 2406 67300 2412 67312
rect 2280 67272 2412 67300
rect 2280 67260 2286 67272
rect 2406 67260 2412 67272
rect 2464 67260 2470 67312
rect 2869 67235 2927 67241
rect 2869 67201 2881 67235
rect 2915 67232 2927 67235
rect 3050 67232 3056 67244
rect 2915 67204 3056 67232
rect 2915 67201 2927 67204
rect 2869 67195 2927 67201
rect 3050 67192 3056 67204
rect 3108 67192 3114 67244
rect 10134 67232 10140 67244
rect 10095 67204 10140 67232
rect 10134 67192 10140 67204
rect 10192 67192 10198 67244
rect 1394 67164 1400 67176
rect 1355 67136 1400 67164
rect 1394 67124 1400 67136
rect 1452 67124 1458 67176
rect 1673 67167 1731 67173
rect 1673 67133 1685 67167
rect 1719 67164 1731 67167
rect 2406 67164 2412 67176
rect 1719 67136 2412 67164
rect 1719 67133 1731 67136
rect 1673 67127 1731 67133
rect 2406 67124 2412 67136
rect 2464 67124 2470 67176
rect 842 67056 848 67108
rect 900 67096 906 67108
rect 2685 67099 2743 67105
rect 2685 67096 2697 67099
rect 900 67068 2697 67096
rect 900 67056 906 67068
rect 2685 67065 2697 67068
rect 2731 67065 2743 67099
rect 2685 67059 2743 67065
rect 1670 66988 1676 67040
rect 1728 67028 1734 67040
rect 1854 67028 1860 67040
rect 1728 67000 1860 67028
rect 1728 66988 1734 67000
rect 1854 66988 1860 67000
rect 1912 66988 1918 67040
rect 5442 66988 5448 67040
rect 5500 67028 5506 67040
rect 9953 67031 10011 67037
rect 9953 67028 9965 67031
rect 5500 67000 9965 67028
rect 5500 66988 5506 67000
rect 9953 66997 9965 67000
rect 9999 66997 10011 67031
rect 9953 66991 10011 66997
rect 1104 66938 10856 66960
rect 1104 66886 2582 66938
rect 2634 66886 2646 66938
rect 2698 66886 2710 66938
rect 2762 66886 2774 66938
rect 2826 66886 2838 66938
rect 2890 66886 5846 66938
rect 5898 66886 5910 66938
rect 5962 66886 5974 66938
rect 6026 66886 6038 66938
rect 6090 66886 6102 66938
rect 6154 66886 9110 66938
rect 9162 66886 9174 66938
rect 9226 66886 9238 66938
rect 9290 66886 9302 66938
rect 9354 66886 9366 66938
rect 9418 66886 10856 66938
rect 1104 66864 10856 66886
rect 8294 66824 8300 66836
rect 1504 66796 8300 66824
rect 1504 66756 1532 66796
rect 8294 66784 8300 66796
rect 8352 66784 8358 66836
rect 1412 66728 1532 66756
rect 1949 66759 2007 66765
rect 1412 66629 1440 66728
rect 1949 66725 1961 66759
rect 1995 66756 2007 66759
rect 5166 66756 5172 66768
rect 1995 66728 5172 66756
rect 1995 66725 2007 66728
rect 1949 66719 2007 66725
rect 5166 66716 5172 66728
rect 5224 66716 5230 66768
rect 1486 66648 1492 66700
rect 1544 66688 1550 66700
rect 2958 66688 2964 66700
rect 1544 66660 1624 66688
rect 1544 66648 1550 66660
rect 1397 66623 1455 66629
rect 1397 66589 1409 66623
rect 1443 66589 1455 66623
rect 1596 66620 1624 66660
rect 1832 66660 2964 66688
rect 1832 66629 1860 66660
rect 2958 66648 2964 66660
rect 3016 66688 3022 66700
rect 3142 66688 3148 66700
rect 3016 66660 3148 66688
rect 3016 66648 3022 66660
rect 3142 66648 3148 66660
rect 3200 66648 3206 66700
rect 1817 66623 1875 66629
rect 1596 66592 1716 66620
rect 1397 66583 1455 66589
rect 1302 66512 1308 66564
rect 1360 66552 1366 66564
rect 1688 66561 1716 66592
rect 1817 66589 1829 66623
rect 1863 66589 1875 66623
rect 2498 66620 2504 66632
rect 2459 66592 2504 66620
rect 1817 66583 1875 66589
rect 2498 66580 2504 66592
rect 2556 66580 2562 66632
rect 10134 66620 10140 66632
rect 10095 66592 10140 66620
rect 10134 66580 10140 66592
rect 10192 66580 10198 66632
rect 1581 66555 1639 66561
rect 1581 66552 1593 66555
rect 1360 66524 1593 66552
rect 1360 66512 1366 66524
rect 1581 66521 1593 66524
rect 1627 66521 1639 66555
rect 1581 66515 1639 66521
rect 1674 66555 1732 66561
rect 1674 66521 1686 66555
rect 1720 66521 1732 66555
rect 1674 66515 1732 66521
rect 1596 66484 1624 66515
rect 2590 66484 2596 66496
rect 1596 66456 2596 66484
rect 2590 66444 2596 66456
rect 2648 66444 2654 66496
rect 2685 66487 2743 66493
rect 2685 66453 2697 66487
rect 2731 66484 2743 66487
rect 2958 66484 2964 66496
rect 2731 66456 2964 66484
rect 2731 66453 2743 66456
rect 2685 66447 2743 66453
rect 2958 66444 2964 66456
rect 3016 66444 3022 66496
rect 8294 66444 8300 66496
rect 8352 66484 8358 66496
rect 9953 66487 10011 66493
rect 9953 66484 9965 66487
rect 8352 66456 9965 66484
rect 8352 66444 8358 66456
rect 9953 66453 9965 66456
rect 9999 66453 10011 66487
rect 9953 66447 10011 66453
rect 1104 66394 10856 66416
rect 1104 66342 4214 66394
rect 4266 66342 4278 66394
rect 4330 66342 4342 66394
rect 4394 66342 4406 66394
rect 4458 66342 4470 66394
rect 4522 66342 7478 66394
rect 7530 66342 7542 66394
rect 7594 66342 7606 66394
rect 7658 66342 7670 66394
rect 7722 66342 7734 66394
rect 7786 66342 10856 66394
rect 1104 66320 10856 66342
rect 1118 66240 1124 66292
rect 1176 66280 1182 66292
rect 1486 66280 1492 66292
rect 1176 66252 1492 66280
rect 1176 66240 1182 66252
rect 1486 66240 1492 66252
rect 1544 66240 1550 66292
rect 1578 66240 1584 66292
rect 1636 66280 1642 66292
rect 1636 66252 1716 66280
rect 1636 66240 1642 66252
rect 1688 66212 1716 66252
rect 1765 66215 1823 66221
rect 1765 66212 1777 66215
rect 1688 66184 1777 66212
rect 1765 66181 1777 66184
rect 1811 66181 1823 66215
rect 3142 66212 3148 66224
rect 1765 66175 1823 66181
rect 2429 66184 3148 66212
rect 1489 66147 1547 66153
rect 1489 66113 1501 66147
rect 1535 66144 1547 66147
rect 1578 66144 1584 66156
rect 1535 66116 1584 66144
rect 1535 66113 1547 66116
rect 1489 66107 1547 66113
rect 1578 66104 1584 66116
rect 1636 66104 1642 66156
rect 1673 66147 1731 66153
rect 1673 66113 1685 66147
rect 1719 66113 1731 66147
rect 1673 66107 1731 66113
rect 1862 66147 1920 66153
rect 1862 66113 1874 66147
rect 1908 66144 1920 66147
rect 2429 66144 2457 66184
rect 3142 66172 3148 66184
rect 3200 66172 3206 66224
rect 1908 66116 2457 66144
rect 2593 66147 2651 66153
rect 1908 66113 1920 66116
rect 1862 66107 1920 66113
rect 2593 66113 2605 66147
rect 2639 66113 2651 66147
rect 10134 66144 10140 66156
rect 10095 66116 10140 66144
rect 2593 66107 2651 66113
rect 1302 65968 1308 66020
rect 1360 66008 1366 66020
rect 1688 66008 1716 66107
rect 2608 66076 2636 66107
rect 10134 66104 10140 66116
rect 10192 66104 10198 66156
rect 1360 65980 1716 66008
rect 1872 66048 2636 66076
rect 1360 65968 1366 65980
rect 1026 65900 1032 65952
rect 1084 65940 1090 65952
rect 1872 65940 1900 66048
rect 2041 66011 2099 66017
rect 2041 65977 2053 66011
rect 2087 66008 2099 66011
rect 4982 66008 4988 66020
rect 2087 65980 4988 66008
rect 2087 65977 2099 65980
rect 2041 65971 2099 65977
rect 4982 65968 4988 65980
rect 5040 65968 5046 66020
rect 1084 65912 1900 65940
rect 2777 65943 2835 65949
rect 1084 65900 1090 65912
rect 2777 65909 2789 65943
rect 2823 65940 2835 65943
rect 3050 65940 3056 65952
rect 2823 65912 3056 65940
rect 2823 65909 2835 65912
rect 2777 65903 2835 65909
rect 3050 65900 3056 65912
rect 3108 65900 3114 65952
rect 9950 65940 9956 65952
rect 9911 65912 9956 65940
rect 9950 65900 9956 65912
rect 10008 65900 10014 65952
rect 1104 65850 10856 65872
rect 1104 65798 2582 65850
rect 2634 65798 2646 65850
rect 2698 65798 2710 65850
rect 2762 65798 2774 65850
rect 2826 65798 2838 65850
rect 2890 65798 5846 65850
rect 5898 65798 5910 65850
rect 5962 65798 5974 65850
rect 6026 65798 6038 65850
rect 6090 65798 6102 65850
rect 6154 65798 9110 65850
rect 9162 65798 9174 65850
rect 9226 65798 9238 65850
rect 9290 65798 9302 65850
rect 9354 65798 9366 65850
rect 9418 65798 10856 65850
rect 1104 65776 10856 65798
rect 1762 65560 1768 65612
rect 1820 65560 1826 65612
rect 9950 65600 9956 65612
rect 2056 65572 9956 65600
rect 1578 65532 1584 65544
rect 1539 65504 1584 65532
rect 1578 65492 1584 65504
rect 1636 65492 1642 65544
rect 1780 65464 1808 65560
rect 2056 65541 2084 65572
rect 9950 65560 9956 65572
rect 10008 65560 10014 65612
rect 2041 65535 2099 65541
rect 2041 65501 2053 65535
rect 2087 65501 2099 65535
rect 2317 65535 2375 65541
rect 2317 65532 2329 65535
rect 2041 65495 2099 65501
rect 2148 65504 2329 65532
rect 2148 65464 2176 65504
rect 2317 65501 2329 65504
rect 2363 65501 2375 65535
rect 2317 65495 2375 65501
rect 2461 65535 2519 65541
rect 2461 65501 2473 65535
rect 2507 65532 2519 65535
rect 2958 65532 2964 65544
rect 2507 65504 2964 65532
rect 2507 65501 2519 65504
rect 2461 65495 2519 65501
rect 2958 65492 2964 65504
rect 3016 65492 3022 65544
rect 3602 65492 3608 65544
rect 3660 65532 3666 65544
rect 3789 65535 3847 65541
rect 3789 65532 3801 65535
rect 3660 65504 3801 65532
rect 3660 65492 3666 65504
rect 3789 65501 3801 65504
rect 3835 65501 3847 65535
rect 3789 65495 3847 65501
rect 1780 65436 2176 65464
rect 2225 65467 2283 65473
rect 2225 65433 2237 65467
rect 2271 65433 2283 65467
rect 2225 65427 2283 65433
rect 382 65356 388 65408
rect 440 65396 446 65408
rect 1397 65399 1455 65405
rect 1397 65396 1409 65399
rect 440 65368 1409 65396
rect 440 65356 446 65368
rect 1397 65365 1409 65368
rect 1443 65365 1455 65399
rect 1397 65359 1455 65365
rect 1854 65356 1860 65408
rect 1912 65396 1918 65408
rect 2240 65396 2268 65427
rect 2774 65424 2780 65476
rect 2832 65464 2838 65476
rect 7834 65464 7840 65476
rect 2832 65436 7840 65464
rect 2832 65424 2838 65436
rect 7834 65424 7840 65436
rect 7892 65424 7898 65476
rect 1912 65368 2268 65396
rect 2610 65399 2668 65405
rect 1912 65356 1918 65368
rect 2610 65365 2622 65399
rect 2656 65396 2668 65399
rect 3694 65396 3700 65408
rect 2656 65368 3700 65396
rect 2656 65365 2668 65368
rect 2610 65359 2668 65365
rect 3694 65356 3700 65368
rect 3752 65356 3758 65408
rect 3970 65396 3976 65408
rect 3931 65368 3976 65396
rect 3970 65356 3976 65368
rect 4028 65356 4034 65408
rect 1104 65306 10856 65328
rect 1104 65254 4214 65306
rect 4266 65254 4278 65306
rect 4330 65254 4342 65306
rect 4394 65254 4406 65306
rect 4458 65254 4470 65306
rect 4522 65254 7478 65306
rect 7530 65254 7542 65306
rect 7594 65254 7606 65306
rect 7658 65254 7670 65306
rect 7722 65254 7734 65306
rect 7786 65254 10856 65306
rect 1104 65232 10856 65254
rect 8294 65192 8300 65204
rect 1412 65164 8300 65192
rect 1412 65065 1440 65164
rect 8294 65152 8300 65164
rect 8352 65152 8358 65204
rect 1486 65084 1492 65136
rect 1544 65124 1550 65136
rect 1966 65127 2024 65133
rect 1966 65124 1978 65127
rect 1544 65096 1978 65124
rect 1544 65084 1550 65096
rect 1966 65093 1978 65096
rect 2012 65093 2024 65127
rect 2685 65127 2743 65133
rect 2685 65124 2697 65127
rect 1966 65087 2024 65093
rect 2148 65096 2697 65124
rect 1397 65059 1455 65065
rect 1397 65025 1409 65059
rect 1443 65025 1455 65059
rect 1397 65019 1455 65025
rect 1581 65059 1639 65065
rect 1581 65025 1593 65059
rect 1627 65025 1639 65059
rect 1581 65019 1639 65025
rect 1673 65059 1731 65065
rect 1673 65025 1685 65059
rect 1719 65025 1731 65059
rect 1673 65019 1731 65025
rect 1770 65059 1828 65065
rect 1770 65025 1782 65059
rect 1816 65025 1828 65059
rect 2148 65056 2176 65096
rect 2685 65093 2697 65096
rect 2731 65093 2743 65127
rect 2685 65087 2743 65093
rect 2777 65127 2835 65133
rect 2777 65093 2789 65127
rect 2823 65124 2835 65127
rect 3234 65124 3240 65136
rect 2823 65096 3240 65124
rect 2823 65093 2835 65096
rect 2777 65087 2835 65093
rect 3234 65084 3240 65096
rect 3292 65084 3298 65136
rect 3694 65084 3700 65136
rect 3752 65124 3758 65136
rect 4890 65124 4896 65136
rect 3752 65096 4896 65124
rect 3752 65084 3758 65096
rect 4890 65084 4896 65096
rect 4948 65084 4954 65136
rect 1770 65019 1828 65025
rect 1872 65028 2176 65056
rect 2501 65059 2559 65065
rect 1302 64948 1308 65000
rect 1360 64988 1366 65000
rect 1596 64988 1624 65019
rect 1360 64960 1624 64988
rect 1360 64948 1366 64960
rect 1394 64880 1400 64932
rect 1452 64920 1458 64932
rect 1688 64920 1716 65019
rect 1452 64892 1716 64920
rect 1452 64880 1458 64892
rect 1780 64852 1808 65019
rect 1872 65000 1900 65028
rect 2501 65025 2513 65059
rect 2547 65025 2559 65059
rect 2501 65019 2559 65025
rect 2869 65059 2927 65065
rect 2869 65025 2881 65059
rect 2915 65056 2927 65059
rect 2958 65056 2964 65068
rect 2915 65028 2964 65056
rect 2915 65025 2927 65028
rect 2869 65019 2927 65025
rect 1854 64948 1860 65000
rect 1912 64948 1918 65000
rect 2516 64988 2544 65019
rect 2958 65016 2964 65028
rect 3016 65016 3022 65068
rect 3142 65016 3148 65068
rect 3200 65056 3206 65068
rect 3510 65056 3516 65068
rect 3200 65028 3372 65056
rect 3471 65028 3516 65056
rect 3200 65016 3206 65028
rect 2774 64988 2780 65000
rect 2516 64960 2780 64988
rect 2774 64948 2780 64960
rect 2832 64948 2838 65000
rect 3344 64988 3372 65028
rect 3510 65016 3516 65028
rect 3568 65016 3574 65068
rect 10134 65056 10140 65068
rect 10095 65028 10140 65056
rect 10134 65016 10140 65028
rect 10192 65016 10198 65068
rect 3697 64991 3755 64997
rect 3697 64988 3709 64991
rect 2884 64960 3709 64988
rect 2884 64852 2912 64960
rect 3697 64957 3709 64960
rect 3743 64957 3755 64991
rect 3697 64951 3755 64957
rect 3053 64923 3111 64929
rect 3053 64889 3065 64923
rect 3099 64920 3111 64923
rect 3142 64920 3148 64932
rect 3099 64892 3148 64920
rect 3099 64889 3111 64892
rect 3053 64883 3111 64889
rect 3142 64880 3148 64892
rect 3200 64880 3206 64932
rect 8294 64880 8300 64932
rect 8352 64920 8358 64932
rect 9953 64923 10011 64929
rect 9953 64920 9965 64923
rect 8352 64892 9965 64920
rect 8352 64880 8358 64892
rect 9953 64889 9965 64892
rect 9999 64889 10011 64923
rect 9953 64883 10011 64889
rect 1780 64824 2912 64852
rect 3234 64812 3240 64864
rect 3292 64852 3298 64864
rect 3510 64852 3516 64864
rect 3292 64824 3516 64852
rect 3292 64812 3298 64824
rect 3510 64812 3516 64824
rect 3568 64812 3574 64864
rect 1104 64762 10856 64784
rect 1104 64710 2582 64762
rect 2634 64710 2646 64762
rect 2698 64710 2710 64762
rect 2762 64710 2774 64762
rect 2826 64710 2838 64762
rect 2890 64710 5846 64762
rect 5898 64710 5910 64762
rect 5962 64710 5974 64762
rect 6026 64710 6038 64762
rect 6090 64710 6102 64762
rect 6154 64710 9110 64762
rect 9162 64710 9174 64762
rect 9226 64710 9238 64762
rect 9290 64710 9302 64762
rect 9354 64710 9366 64762
rect 9418 64710 10856 64762
rect 1104 64688 10856 64710
rect 1762 64540 1768 64592
rect 1820 64580 1826 64592
rect 2222 64580 2228 64592
rect 1820 64552 2228 64580
rect 1820 64540 1826 64552
rect 2222 64540 2228 64552
rect 2280 64540 2286 64592
rect 2501 64583 2559 64589
rect 2501 64549 2513 64583
rect 2547 64580 2559 64583
rect 3510 64580 3516 64592
rect 2547 64552 3516 64580
rect 2547 64549 2559 64552
rect 2501 64543 2559 64549
rect 3510 64540 3516 64552
rect 3568 64540 3574 64592
rect 8294 64512 8300 64524
rect 1964 64484 8300 64512
rect 1964 64453 1992 64484
rect 8294 64472 8300 64484
rect 8352 64472 8358 64524
rect 1949 64447 2007 64453
rect 1949 64413 1961 64447
rect 1995 64413 2007 64447
rect 2222 64444 2228 64456
rect 2183 64416 2228 64444
rect 1949 64407 2007 64413
rect 2222 64404 2228 64416
rect 2280 64404 2286 64456
rect 2369 64447 2427 64453
rect 2369 64413 2381 64447
rect 2415 64444 2427 64447
rect 2958 64444 2964 64456
rect 2415 64416 2964 64444
rect 2415 64413 2427 64416
rect 2369 64407 2427 64413
rect 2958 64404 2964 64416
rect 3016 64404 3022 64456
rect 3789 64447 3847 64453
rect 3789 64413 3801 64447
rect 3835 64444 3847 64447
rect 4062 64444 4068 64456
rect 3835 64416 4068 64444
rect 3835 64413 3847 64416
rect 3789 64407 3847 64413
rect 4062 64404 4068 64416
rect 4120 64404 4126 64456
rect 10134 64444 10140 64456
rect 10095 64416 10140 64444
rect 10134 64404 10140 64416
rect 10192 64404 10198 64456
rect 1854 64336 1860 64388
rect 1912 64376 1918 64388
rect 2133 64379 2191 64385
rect 2133 64376 2145 64379
rect 1912 64348 2145 64376
rect 1912 64336 1918 64348
rect 2133 64345 2145 64348
rect 2179 64345 2191 64379
rect 2133 64339 2191 64345
rect 3050 64268 3056 64320
rect 3108 64308 3114 64320
rect 3973 64311 4031 64317
rect 3973 64308 3985 64311
rect 3108 64280 3985 64308
rect 3108 64268 3114 64280
rect 3973 64277 3985 64280
rect 4019 64277 4031 64311
rect 3973 64271 4031 64277
rect 8294 64268 8300 64320
rect 8352 64308 8358 64320
rect 9953 64311 10011 64317
rect 9953 64308 9965 64311
rect 8352 64280 9965 64308
rect 8352 64268 8358 64280
rect 9953 64277 9965 64280
rect 9999 64277 10011 64311
rect 9953 64271 10011 64277
rect 1104 64218 10856 64240
rect 1104 64166 4214 64218
rect 4266 64166 4278 64218
rect 4330 64166 4342 64218
rect 4394 64166 4406 64218
rect 4458 64166 4470 64218
rect 4522 64166 7478 64218
rect 7530 64166 7542 64218
rect 7594 64166 7606 64218
rect 7658 64166 7670 64218
rect 7722 64166 7734 64218
rect 7786 64166 10856 64218
rect 1104 64144 10856 64166
rect 1302 63996 1308 64048
rect 1360 64036 1366 64048
rect 3789 64039 3847 64045
rect 3789 64036 3801 64039
rect 1360 64008 3801 64036
rect 1360 63996 1366 64008
rect 3789 64005 3801 64008
rect 3835 64005 3847 64039
rect 3789 63999 3847 64005
rect 290 63928 296 63980
rect 348 63968 354 63980
rect 1397 63971 1455 63977
rect 1397 63968 1409 63971
rect 348 63940 1409 63968
rect 348 63928 354 63940
rect 1397 63937 1409 63940
rect 1443 63937 1455 63971
rect 1397 63931 1455 63937
rect 2593 63971 2651 63977
rect 2593 63937 2605 63971
rect 2639 63968 2651 63971
rect 3234 63968 3240 63980
rect 2639 63940 3240 63968
rect 2639 63937 2651 63940
rect 2593 63931 2651 63937
rect 3234 63928 3240 63940
rect 3292 63928 3298 63980
rect 3513 63971 3571 63977
rect 3513 63937 3525 63971
rect 3559 63968 3571 63971
rect 3694 63968 3700 63980
rect 3559 63940 3700 63968
rect 3559 63937 3571 63940
rect 3513 63931 3571 63937
rect 3694 63928 3700 63940
rect 3752 63928 3758 63980
rect 2869 63903 2927 63909
rect 2869 63869 2881 63903
rect 2915 63900 2927 63903
rect 2958 63900 2964 63912
rect 2915 63872 2964 63900
rect 2915 63869 2927 63872
rect 2869 63863 2927 63869
rect 2958 63860 2964 63872
rect 3016 63860 3022 63912
rect 1578 63764 1584 63776
rect 1539 63736 1584 63764
rect 1578 63724 1584 63736
rect 1636 63724 1642 63776
rect 1104 63674 10856 63696
rect 1104 63622 2582 63674
rect 2634 63622 2646 63674
rect 2698 63622 2710 63674
rect 2762 63622 2774 63674
rect 2826 63622 2838 63674
rect 2890 63622 5846 63674
rect 5898 63622 5910 63674
rect 5962 63622 5974 63674
rect 6026 63622 6038 63674
rect 6090 63622 6102 63674
rect 6154 63622 9110 63674
rect 9162 63622 9174 63674
rect 9226 63622 9238 63674
rect 9290 63622 9302 63674
rect 9354 63622 9366 63674
rect 9418 63622 10856 63674
rect 1104 63600 10856 63622
rect 1670 63452 1676 63504
rect 1728 63492 1734 63504
rect 2317 63495 2375 63501
rect 2317 63492 2329 63495
rect 1728 63464 2329 63492
rect 1728 63452 1734 63464
rect 2317 63461 2329 63464
rect 2363 63461 2375 63495
rect 3050 63492 3056 63504
rect 3011 63464 3056 63492
rect 2317 63455 2375 63461
rect 3050 63452 3056 63464
rect 3108 63452 3114 63504
rect 1397 63359 1455 63365
rect 1397 63325 1409 63359
rect 1443 63325 1455 63359
rect 1397 63319 1455 63325
rect 1412 63288 1440 63319
rect 1670 63316 1676 63368
rect 1728 63356 1734 63368
rect 2133 63359 2191 63365
rect 2133 63356 2145 63359
rect 1728 63328 2145 63356
rect 1728 63316 1734 63328
rect 2133 63325 2145 63328
rect 2179 63325 2191 63359
rect 2866 63356 2872 63368
rect 2827 63328 2872 63356
rect 2133 63319 2191 63325
rect 2866 63316 2872 63328
rect 2924 63316 2930 63368
rect 10134 63356 10140 63368
rect 10095 63328 10140 63356
rect 10134 63316 10140 63328
rect 10192 63316 10198 63368
rect 3234 63288 3240 63300
rect 1412 63260 3240 63288
rect 3234 63248 3240 63260
rect 3292 63248 3298 63300
rect 1394 63180 1400 63232
rect 1452 63220 1458 63232
rect 1581 63223 1639 63229
rect 1581 63220 1593 63223
rect 1452 63192 1593 63220
rect 1452 63180 1458 63192
rect 1581 63189 1593 63192
rect 1627 63189 1639 63223
rect 1581 63183 1639 63189
rect 8478 63180 8484 63232
rect 8536 63220 8542 63232
rect 9953 63223 10011 63229
rect 9953 63220 9965 63223
rect 8536 63192 9965 63220
rect 8536 63180 8542 63192
rect 9953 63189 9965 63192
rect 9999 63189 10011 63223
rect 9953 63183 10011 63189
rect 566 63112 572 63164
rect 624 63152 630 63164
rect 934 63152 940 63164
rect 624 63124 940 63152
rect 624 63112 630 63124
rect 934 63112 940 63124
rect 992 63112 998 63164
rect 1104 63130 10856 63152
rect 1104 63078 4214 63130
rect 4266 63078 4278 63130
rect 4330 63078 4342 63130
rect 4394 63078 4406 63130
rect 4458 63078 4470 63130
rect 4522 63078 7478 63130
rect 7530 63078 7542 63130
rect 7594 63078 7606 63130
rect 7658 63078 7670 63130
rect 7722 63078 7734 63130
rect 7786 63078 10856 63130
rect 1104 63056 10856 63078
rect 1026 62840 1032 62892
rect 1084 62880 1090 62892
rect 1397 62883 1455 62889
rect 1397 62880 1409 62883
rect 1084 62852 1409 62880
rect 1084 62840 1090 62852
rect 1397 62849 1409 62852
rect 1443 62849 1455 62883
rect 1397 62843 1455 62849
rect 2133 62883 2191 62889
rect 2133 62849 2145 62883
rect 2179 62880 2191 62883
rect 3050 62880 3056 62892
rect 2179 62852 3056 62880
rect 2179 62849 2191 62852
rect 2133 62843 2191 62849
rect 3050 62840 3056 62852
rect 3108 62840 3114 62892
rect 10134 62880 10140 62892
rect 10095 62852 10140 62880
rect 10134 62840 10140 62852
rect 10192 62840 10198 62892
rect 1578 62676 1584 62688
rect 1539 62648 1584 62676
rect 1578 62636 1584 62648
rect 1636 62636 1642 62688
rect 2314 62676 2320 62688
rect 2275 62648 2320 62676
rect 2314 62636 2320 62648
rect 2372 62636 2378 62688
rect 6178 62636 6184 62688
rect 6236 62676 6242 62688
rect 9953 62679 10011 62685
rect 9953 62676 9965 62679
rect 6236 62648 9965 62676
rect 6236 62636 6242 62648
rect 9953 62645 9965 62648
rect 9999 62645 10011 62679
rect 9953 62639 10011 62645
rect 1104 62586 10856 62608
rect 1104 62534 2582 62586
rect 2634 62534 2646 62586
rect 2698 62534 2710 62586
rect 2762 62534 2774 62586
rect 2826 62534 2838 62586
rect 2890 62534 5846 62586
rect 5898 62534 5910 62586
rect 5962 62534 5974 62586
rect 6026 62534 6038 62586
rect 6090 62534 6102 62586
rect 6154 62534 9110 62586
rect 9162 62534 9174 62586
rect 9226 62534 9238 62586
rect 9290 62534 9302 62586
rect 9354 62534 9366 62586
rect 9418 62534 10856 62586
rect 1104 62512 10856 62534
rect 2501 62407 2559 62413
rect 2501 62373 2513 62407
rect 2547 62404 2559 62407
rect 5350 62404 5356 62416
rect 2547 62376 5356 62404
rect 2547 62373 2559 62376
rect 2501 62367 2559 62373
rect 5350 62364 5356 62376
rect 5408 62364 5414 62416
rect 8294 62336 8300 62348
rect 1964 62308 8300 62336
rect 1964 62277 1992 62308
rect 8294 62296 8300 62308
rect 8352 62296 8358 62348
rect 2406 62277 2412 62280
rect 1949 62271 2007 62277
rect 1949 62237 1961 62271
rect 1995 62237 2007 62271
rect 2225 62271 2283 62277
rect 2225 62268 2237 62271
rect 1949 62231 2007 62237
rect 2056 62240 2237 62268
rect 1118 62160 1124 62212
rect 1176 62200 1182 62212
rect 2056 62200 2084 62240
rect 2225 62237 2237 62240
rect 2271 62237 2283 62271
rect 2225 62231 2283 62237
rect 2369 62271 2412 62277
rect 2369 62237 2381 62271
rect 2464 62268 2470 62280
rect 2958 62268 2964 62280
rect 2464 62240 2964 62268
rect 2369 62231 2412 62237
rect 2406 62228 2412 62231
rect 2464 62228 2470 62240
rect 2958 62228 2964 62240
rect 3016 62228 3022 62280
rect 10134 62268 10140 62280
rect 10095 62240 10140 62268
rect 10134 62228 10140 62240
rect 10192 62228 10198 62280
rect 1176 62172 2084 62200
rect 2133 62203 2191 62209
rect 1176 62160 1182 62172
rect 2133 62169 2145 62203
rect 2179 62200 2191 62203
rect 2590 62200 2596 62212
rect 2179 62172 2596 62200
rect 2179 62169 2191 62172
rect 2133 62163 2191 62169
rect 1854 62092 1860 62144
rect 1912 62132 1918 62144
rect 2148 62132 2176 62163
rect 2590 62160 2596 62172
rect 2648 62160 2654 62212
rect 1912 62104 2176 62132
rect 1912 62092 1918 62104
rect 2958 62092 2964 62144
rect 3016 62132 3022 62144
rect 3510 62132 3516 62144
rect 3016 62104 3516 62132
rect 3016 62092 3022 62104
rect 3510 62092 3516 62104
rect 3568 62092 3574 62144
rect 8294 62092 8300 62144
rect 8352 62132 8358 62144
rect 9953 62135 10011 62141
rect 9953 62132 9965 62135
rect 8352 62104 9965 62132
rect 8352 62092 8358 62104
rect 9953 62101 9965 62104
rect 9999 62101 10011 62135
rect 9953 62095 10011 62101
rect 1104 62042 10856 62064
rect 1104 61990 4214 62042
rect 4266 61990 4278 62042
rect 4330 61990 4342 62042
rect 4394 61990 4406 62042
rect 4458 61990 4470 62042
rect 4522 61990 7478 62042
rect 7530 61990 7542 62042
rect 7594 61990 7606 62042
rect 7658 61990 7670 62042
rect 7722 61990 7734 62042
rect 7786 61990 10856 62042
rect 1104 61968 10856 61990
rect 9950 61860 9956 61872
rect 1412 61832 9956 61860
rect 1412 61801 1440 61832
rect 9950 61820 9956 61832
rect 10008 61820 10014 61872
rect 1397 61795 1455 61801
rect 1397 61761 1409 61795
rect 1443 61761 1455 61795
rect 1397 61755 1455 61761
rect 1486 61752 1492 61804
rect 1544 61792 1550 61804
rect 1581 61795 1639 61801
rect 1581 61792 1593 61795
rect 1544 61764 1593 61792
rect 1544 61752 1550 61764
rect 1581 61761 1593 61764
rect 1627 61761 1639 61795
rect 1581 61755 1639 61761
rect 1673 61795 1731 61801
rect 1673 61761 1685 61795
rect 1719 61761 1731 61795
rect 1673 61755 1731 61761
rect 1596 61656 1624 61755
rect 1688 61724 1716 61755
rect 1762 61752 1768 61804
rect 1820 61801 1826 61804
rect 1820 61792 1828 61801
rect 2406 61792 2412 61804
rect 1820 61764 2412 61792
rect 1820 61755 1828 61764
rect 1820 61752 1826 61755
rect 2406 61752 2412 61764
rect 2464 61752 2470 61804
rect 2593 61795 2651 61801
rect 2593 61761 2605 61795
rect 2639 61792 2651 61795
rect 2682 61792 2688 61804
rect 2639 61764 2688 61792
rect 2639 61761 2651 61764
rect 2593 61755 2651 61761
rect 2682 61752 2688 61764
rect 2740 61752 2746 61804
rect 3510 61792 3516 61804
rect 3471 61764 3516 61792
rect 3510 61752 3516 61764
rect 3568 61752 3574 61804
rect 2222 61724 2228 61736
rect 1688 61696 2228 61724
rect 2222 61684 2228 61696
rect 2280 61684 2286 61736
rect 2777 61727 2835 61733
rect 2777 61693 2789 61727
rect 2823 61693 2835 61727
rect 2777 61687 2835 61693
rect 2590 61656 2596 61668
rect 1596 61628 2596 61656
rect 2590 61616 2596 61628
rect 2648 61656 2654 61668
rect 2792 61656 2820 61687
rect 3694 61656 3700 61668
rect 2648 61628 2820 61656
rect 3655 61628 3700 61656
rect 2648 61616 2654 61628
rect 3694 61616 3700 61628
rect 3752 61616 3758 61668
rect 1854 61548 1860 61600
rect 1912 61588 1918 61600
rect 1949 61591 2007 61597
rect 1949 61588 1961 61591
rect 1912 61560 1961 61588
rect 1912 61548 1918 61560
rect 1949 61557 1961 61560
rect 1995 61557 2007 61591
rect 1949 61551 2007 61557
rect 2130 61548 2136 61600
rect 2188 61588 2194 61600
rect 2406 61588 2412 61600
rect 2188 61560 2412 61588
rect 2188 61548 2194 61560
rect 2406 61548 2412 61560
rect 2464 61548 2470 61600
rect 1104 61498 10856 61520
rect 1104 61446 2582 61498
rect 2634 61446 2646 61498
rect 2698 61446 2710 61498
rect 2762 61446 2774 61498
rect 2826 61446 2838 61498
rect 2890 61446 5846 61498
rect 5898 61446 5910 61498
rect 5962 61446 5974 61498
rect 6026 61446 6038 61498
rect 6090 61446 6102 61498
rect 6154 61446 9110 61498
rect 9162 61446 9174 61498
rect 9226 61446 9238 61498
rect 9290 61446 9302 61498
rect 9354 61446 9366 61498
rect 9418 61446 10856 61498
rect 1104 61424 10856 61446
rect 9950 61384 9956 61396
rect 9911 61356 9956 61384
rect 9950 61344 9956 61356
rect 10008 61344 10014 61396
rect 1949 61319 2007 61325
rect 1949 61285 1961 61319
rect 1995 61316 2007 61319
rect 2222 61316 2228 61328
rect 1995 61288 2228 61316
rect 1995 61285 2007 61288
rect 1949 61279 2007 61285
rect 2222 61276 2228 61288
rect 2280 61276 2286 61328
rect 8294 61248 8300 61260
rect 1412 61220 8300 61248
rect 1412 61189 1440 61220
rect 8294 61208 8300 61220
rect 8352 61208 8358 61260
rect 1397 61183 1455 61189
rect 1397 61149 1409 61183
rect 1443 61149 1455 61183
rect 1397 61143 1455 61149
rect 1762 61140 1768 61192
rect 1820 61189 1826 61192
rect 1820 61180 1828 61189
rect 2501 61183 2559 61189
rect 1820 61152 1865 61180
rect 1820 61143 1828 61152
rect 2501 61149 2513 61183
rect 2547 61149 2559 61183
rect 10134 61180 10140 61192
rect 10095 61152 10140 61180
rect 2501 61143 2559 61149
rect 1820 61140 1826 61143
rect 1118 61072 1124 61124
rect 1176 61112 1182 61124
rect 1486 61112 1492 61124
rect 1176 61084 1492 61112
rect 1176 61072 1182 61084
rect 1486 61072 1492 61084
rect 1544 61112 1550 61124
rect 1581 61115 1639 61121
rect 1581 61112 1593 61115
rect 1544 61084 1593 61112
rect 1544 61072 1550 61084
rect 1581 61081 1593 61084
rect 1627 61081 1639 61115
rect 1581 61075 1639 61081
rect 1670 61072 1676 61124
rect 1728 61112 1734 61124
rect 1728 61084 1773 61112
rect 1728 61072 1734 61084
rect 14 61004 20 61056
rect 72 61044 78 61056
rect 2516 61044 2544 61143
rect 10134 61140 10140 61152
rect 10192 61140 10198 61192
rect 72 61016 2544 61044
rect 2685 61047 2743 61053
rect 72 61004 78 61016
rect 2685 61013 2697 61047
rect 2731 61044 2743 61047
rect 2774 61044 2780 61056
rect 2731 61016 2780 61044
rect 2731 61013 2743 61016
rect 2685 61007 2743 61013
rect 2774 61004 2780 61016
rect 2832 61004 2838 61056
rect 1104 60954 10856 60976
rect 1104 60902 4214 60954
rect 4266 60902 4278 60954
rect 4330 60902 4342 60954
rect 4394 60902 4406 60954
rect 4458 60902 4470 60954
rect 4522 60902 7478 60954
rect 7530 60902 7542 60954
rect 7594 60902 7606 60954
rect 7658 60902 7670 60954
rect 7722 60902 7734 60954
rect 7786 60902 10856 60954
rect 1104 60880 10856 60902
rect 842 60800 848 60852
rect 900 60800 906 60852
rect 1210 60800 1216 60852
rect 1268 60840 1274 60852
rect 1670 60840 1676 60852
rect 1268 60812 1676 60840
rect 1268 60800 1274 60812
rect 1670 60800 1676 60812
rect 1728 60800 1734 60852
rect 1946 60800 1952 60852
rect 2004 60840 2010 60852
rect 2682 60840 2688 60852
rect 2004 60812 2688 60840
rect 2004 60800 2010 60812
rect 2682 60800 2688 60812
rect 2740 60800 2746 60852
rect 860 60772 888 60800
rect 1486 60772 1492 60784
rect 860 60744 1492 60772
rect 1486 60732 1492 60744
rect 1544 60732 1550 60784
rect 1397 60707 1455 60713
rect 1397 60673 1409 60707
rect 1443 60704 1455 60707
rect 1443 60676 1716 60704
rect 1443 60673 1455 60676
rect 1397 60667 1455 60673
rect 1688 60568 1716 60676
rect 1762 60664 1768 60716
rect 1820 60704 1826 60716
rect 2133 60707 2191 60713
rect 2133 60704 2145 60707
rect 1820 60676 2145 60704
rect 1820 60664 1826 60676
rect 2133 60673 2145 60676
rect 2179 60673 2191 60707
rect 2133 60667 2191 60673
rect 2869 60707 2927 60713
rect 2869 60673 2881 60707
rect 2915 60673 2927 60707
rect 2869 60667 2927 60673
rect 2884 60636 2912 60667
rect 3234 60664 3240 60716
rect 3292 60704 3298 60716
rect 3418 60704 3424 60716
rect 3292 60676 3424 60704
rect 3292 60664 3298 60676
rect 3418 60664 3424 60676
rect 3476 60664 3482 60716
rect 10134 60704 10140 60716
rect 10095 60676 10140 60704
rect 10134 60664 10140 60676
rect 10192 60664 10198 60716
rect 3970 60636 3976 60648
rect 2884 60608 3976 60636
rect 3970 60596 3976 60608
rect 4028 60596 4034 60648
rect 1412 60540 1716 60568
rect 1210 60460 1216 60512
rect 1268 60500 1274 60512
rect 1412 60500 1440 60540
rect 2958 60528 2964 60580
rect 3016 60568 3022 60580
rect 3053 60571 3111 60577
rect 3053 60568 3065 60571
rect 3016 60540 3065 60568
rect 3016 60528 3022 60540
rect 3053 60537 3065 60540
rect 3099 60537 3111 60571
rect 3053 60531 3111 60537
rect 1578 60500 1584 60512
rect 1268 60472 1440 60500
rect 1539 60472 1584 60500
rect 1268 60460 1274 60472
rect 1578 60460 1584 60472
rect 1636 60460 1642 60512
rect 2314 60500 2320 60512
rect 2275 60472 2320 60500
rect 2314 60460 2320 60472
rect 2372 60460 2378 60512
rect 9950 60500 9956 60512
rect 9911 60472 9956 60500
rect 9950 60460 9956 60472
rect 10008 60460 10014 60512
rect 1104 60410 10856 60432
rect 1104 60358 2582 60410
rect 2634 60358 2646 60410
rect 2698 60358 2710 60410
rect 2762 60358 2774 60410
rect 2826 60358 2838 60410
rect 2890 60358 5846 60410
rect 5898 60358 5910 60410
rect 5962 60358 5974 60410
rect 6026 60358 6038 60410
rect 6090 60358 6102 60410
rect 6154 60358 9110 60410
rect 9162 60358 9174 60410
rect 9226 60358 9238 60410
rect 9290 60358 9302 60410
rect 9354 60358 9366 60410
rect 9418 60358 10856 60410
rect 1104 60336 10856 60358
rect 106 60256 112 60308
rect 164 60296 170 60308
rect 1762 60296 1768 60308
rect 164 60268 1768 60296
rect 164 60256 170 60268
rect 1762 60256 1768 60268
rect 1820 60256 1826 60308
rect 566 60188 572 60240
rect 624 60228 630 60240
rect 1302 60228 1308 60240
rect 624 60200 1308 60228
rect 624 60188 630 60200
rect 1302 60188 1308 60200
rect 1360 60188 1366 60240
rect 2222 60188 2228 60240
rect 2280 60228 2286 60240
rect 2682 60228 2688 60240
rect 2280 60200 2688 60228
rect 2280 60188 2286 60200
rect 2682 60188 2688 60200
rect 2740 60188 2746 60240
rect 750 60120 756 60172
rect 808 60160 814 60172
rect 2590 60160 2596 60172
rect 808 60132 2596 60160
rect 808 60120 814 60132
rect 2590 60120 2596 60132
rect 2648 60120 2654 60172
rect 474 60052 480 60104
rect 532 60092 538 60104
rect 2225 60095 2283 60101
rect 2225 60092 2237 60095
rect 532 60064 2237 60092
rect 532 60052 538 60064
rect 2225 60061 2237 60064
rect 2271 60092 2283 60095
rect 2777 60095 2835 60101
rect 2777 60092 2789 60095
rect 2271 60064 2789 60092
rect 2271 60061 2283 60064
rect 2225 60055 2283 60061
rect 2777 60061 2789 60064
rect 2823 60061 2835 60095
rect 2777 60055 2835 60061
rect 1762 59984 1768 60036
rect 1820 60024 1826 60036
rect 2498 60024 2504 60036
rect 1820 59996 2504 60024
rect 1820 59984 1826 59996
rect 2498 59984 2504 59996
rect 2556 59984 2562 60036
rect 2038 59956 2044 59968
rect 1044 59928 2044 59956
rect 1044 59684 1072 59928
rect 2038 59916 2044 59928
rect 2096 59916 2102 59968
rect 2593 59959 2651 59965
rect 2593 59925 2605 59959
rect 2639 59956 2651 59959
rect 2774 59956 2780 59968
rect 2639 59928 2780 59956
rect 2639 59925 2651 59928
rect 2593 59919 2651 59925
rect 2774 59916 2780 59928
rect 2832 59916 2838 59968
rect 1104 59866 10856 59888
rect 1104 59814 4214 59866
rect 4266 59814 4278 59866
rect 4330 59814 4342 59866
rect 4394 59814 4406 59866
rect 4458 59814 4470 59866
rect 4522 59814 7478 59866
rect 7530 59814 7542 59866
rect 7594 59814 7606 59866
rect 7658 59814 7670 59866
rect 7722 59814 7734 59866
rect 7786 59814 10856 59866
rect 1104 59792 10856 59814
rect 1118 59712 1124 59764
rect 1176 59752 1182 59764
rect 2038 59752 2044 59764
rect 1176 59724 2044 59752
rect 1176 59712 1182 59724
rect 1596 59693 1624 59724
rect 2038 59712 2044 59724
rect 2096 59712 2102 59764
rect 2590 59752 2596 59764
rect 2424 59724 2596 59752
rect 2424 59693 2452 59724
rect 2590 59712 2596 59724
rect 2648 59712 2654 59764
rect 1581 59687 1639 59693
rect 1044 59656 1532 59684
rect 1118 59576 1124 59628
rect 1176 59616 1182 59628
rect 1397 59619 1455 59625
rect 1397 59616 1409 59619
rect 1176 59588 1409 59616
rect 1176 59576 1182 59588
rect 1397 59585 1409 59588
rect 1443 59585 1455 59619
rect 1504 59616 1532 59656
rect 1581 59653 1593 59687
rect 1627 59653 1639 59687
rect 1581 59647 1639 59653
rect 1673 59687 1731 59693
rect 1673 59653 1685 59687
rect 1719 59653 1731 59687
rect 2317 59687 2375 59693
rect 1673 59647 1731 59653
rect 1785 59656 2009 59684
rect 1688 59616 1716 59647
rect 1785 59625 1813 59656
rect 1504 59588 1716 59616
rect 1770 59619 1828 59625
rect 1397 59579 1455 59585
rect 1770 59585 1782 59619
rect 1816 59585 1828 59619
rect 1770 59579 1828 59585
rect 1981 59548 2009 59656
rect 2317 59653 2329 59687
rect 2363 59653 2375 59687
rect 2317 59647 2375 59653
rect 2409 59687 2467 59693
rect 2409 59653 2421 59687
rect 2455 59653 2467 59687
rect 2409 59647 2467 59653
rect 2130 59576 2136 59628
rect 2188 59616 2194 59628
rect 2188 59588 2233 59616
rect 2188 59576 2194 59588
rect 1981 59520 2084 59548
rect 750 59372 756 59424
rect 808 59412 814 59424
rect 1949 59415 2007 59421
rect 1949 59412 1961 59415
rect 808 59384 1961 59412
rect 808 59372 814 59384
rect 1949 59381 1961 59384
rect 1995 59381 2007 59415
rect 2056 59412 2084 59520
rect 2332 59492 2360 59647
rect 2590 59625 2596 59628
rect 2553 59619 2596 59625
rect 2553 59585 2565 59619
rect 2553 59579 2596 59585
rect 2590 59576 2596 59579
rect 2648 59576 2654 59628
rect 10134 59616 10140 59628
rect 10095 59588 10140 59616
rect 10134 59576 10140 59588
rect 10192 59576 10198 59628
rect 2682 59548 2688 59560
rect 2424 59520 2688 59548
rect 2424 59492 2452 59520
rect 2682 59508 2688 59520
rect 2740 59508 2746 59560
rect 5074 59508 5080 59560
rect 5132 59548 5138 59560
rect 9950 59548 9956 59560
rect 5132 59520 9956 59548
rect 5132 59508 5138 59520
rect 9950 59508 9956 59520
rect 10008 59508 10014 59560
rect 2314 59440 2320 59492
rect 2372 59440 2378 59492
rect 2406 59440 2412 59492
rect 2464 59440 2470 59492
rect 2130 59412 2136 59424
rect 2056 59384 2136 59412
rect 1949 59375 2007 59381
rect 2130 59372 2136 59384
rect 2188 59372 2194 59424
rect 2222 59372 2228 59424
rect 2280 59412 2286 59424
rect 2685 59415 2743 59421
rect 2685 59412 2697 59415
rect 2280 59384 2697 59412
rect 2280 59372 2286 59384
rect 2685 59381 2697 59384
rect 2731 59381 2743 59415
rect 2685 59375 2743 59381
rect 3234 59372 3240 59424
rect 3292 59412 3298 59424
rect 3694 59412 3700 59424
rect 3292 59384 3700 59412
rect 3292 59372 3298 59384
rect 3694 59372 3700 59384
rect 3752 59372 3758 59424
rect 3970 59372 3976 59424
rect 4028 59412 4034 59424
rect 4614 59412 4620 59424
rect 4028 59384 4620 59412
rect 4028 59372 4034 59384
rect 4614 59372 4620 59384
rect 4672 59372 4678 59424
rect 8294 59372 8300 59424
rect 8352 59412 8358 59424
rect 9953 59415 10011 59421
rect 9953 59412 9965 59415
rect 8352 59384 9965 59412
rect 8352 59372 8358 59384
rect 9953 59381 9965 59384
rect 9999 59381 10011 59415
rect 9953 59375 10011 59381
rect 1104 59322 10856 59344
rect 1104 59270 2582 59322
rect 2634 59270 2646 59322
rect 2698 59270 2710 59322
rect 2762 59270 2774 59322
rect 2826 59270 2838 59322
rect 2890 59270 5846 59322
rect 5898 59270 5910 59322
rect 5962 59270 5974 59322
rect 6026 59270 6038 59322
rect 6090 59270 6102 59322
rect 6154 59270 9110 59322
rect 9162 59270 9174 59322
rect 9226 59270 9238 59322
rect 9290 59270 9302 59322
rect 9354 59270 9366 59322
rect 9418 59270 10856 59322
rect 1104 59248 10856 59270
rect 1397 59211 1455 59217
rect 1397 59177 1409 59211
rect 1443 59208 1455 59211
rect 1946 59208 1952 59220
rect 1443 59180 1952 59208
rect 1443 59177 1455 59180
rect 1397 59171 1455 59177
rect 1946 59168 1952 59180
rect 2004 59168 2010 59220
rect 2038 59168 2044 59220
rect 2096 59208 2102 59220
rect 2314 59208 2320 59220
rect 2096 59180 2320 59208
rect 2096 59168 2102 59180
rect 2314 59168 2320 59180
rect 2372 59168 2378 59220
rect 566 59100 572 59152
rect 624 59140 630 59152
rect 2593 59143 2651 59149
rect 2593 59140 2605 59143
rect 624 59112 2605 59140
rect 624 59100 630 59112
rect 2593 59109 2605 59112
rect 2639 59109 2651 59143
rect 2593 59103 2651 59109
rect 8478 59072 8484 59084
rect 2056 59044 8484 59072
rect 1578 59004 1584 59016
rect 1539 58976 1584 59004
rect 1578 58964 1584 58976
rect 1636 58964 1642 59016
rect 2056 59013 2084 59044
rect 8478 59032 8484 59044
rect 8536 59032 8542 59084
rect 2041 59007 2099 59013
rect 2041 58973 2053 59007
rect 2087 58973 2099 59007
rect 2317 59007 2375 59013
rect 2317 59004 2329 59007
rect 2041 58967 2099 58973
rect 2148 58976 2329 59004
rect 1394 58896 1400 58948
rect 1452 58936 1458 58948
rect 2148 58936 2176 58976
rect 2317 58973 2329 58976
rect 2363 58973 2375 59007
rect 2317 58967 2375 58973
rect 2461 59007 2519 59013
rect 2461 58973 2473 59007
rect 2507 59004 2519 59007
rect 3789 59007 3847 59013
rect 2507 58976 2728 59004
rect 2507 58973 2519 58976
rect 2461 58967 2519 58973
rect 1452 58908 2176 58936
rect 2225 58939 2283 58945
rect 1452 58896 1458 58908
rect 2225 58905 2237 58939
rect 2271 58936 2283 58939
rect 2590 58936 2596 58948
rect 2271 58908 2596 58936
rect 2271 58905 2283 58908
rect 2225 58899 2283 58905
rect 2590 58896 2596 58908
rect 2648 58896 2654 58948
rect 382 58828 388 58880
rect 440 58868 446 58880
rect 2038 58868 2044 58880
rect 440 58840 2044 58868
rect 440 58828 446 58840
rect 2038 58828 2044 58840
rect 2096 58828 2102 58880
rect 2130 58828 2136 58880
rect 2188 58868 2194 58880
rect 2700 58868 2728 58976
rect 3789 58973 3801 59007
rect 3835 59004 3847 59007
rect 4706 59004 4712 59016
rect 3835 58976 4712 59004
rect 3835 58973 3847 58976
rect 3789 58967 3847 58973
rect 4706 58964 4712 58976
rect 4764 58964 4770 59016
rect 10134 59004 10140 59016
rect 10095 58976 10140 59004
rect 10134 58964 10140 58976
rect 10192 58964 10198 59016
rect 3970 58868 3976 58880
rect 2188 58840 2728 58868
rect 3931 58840 3976 58868
rect 2188 58828 2194 58840
rect 3970 58828 3976 58840
rect 4028 58828 4034 58880
rect 9950 58868 9956 58880
rect 9911 58840 9956 58868
rect 9950 58828 9956 58840
rect 10008 58828 10014 58880
rect 1104 58778 10856 58800
rect 1104 58726 4214 58778
rect 4266 58726 4278 58778
rect 4330 58726 4342 58778
rect 4394 58726 4406 58778
rect 4458 58726 4470 58778
rect 4522 58726 7478 58778
rect 7530 58726 7542 58778
rect 7594 58726 7606 58778
rect 7658 58726 7670 58778
rect 7722 58726 7734 58778
rect 7786 58726 10856 58778
rect 1104 58704 10856 58726
rect 1578 58624 1584 58676
rect 1636 58664 1642 58676
rect 2869 58667 2927 58673
rect 2869 58664 2881 58667
rect 1636 58636 2881 58664
rect 1636 58624 1642 58636
rect 2869 58633 2881 58636
rect 2915 58633 2927 58667
rect 2869 58627 2927 58633
rect 750 58556 756 58608
rect 808 58596 814 58608
rect 2222 58596 2228 58608
rect 808 58568 2228 58596
rect 808 58556 814 58568
rect 2222 58556 2228 58568
rect 2280 58556 2286 58608
rect 2314 58556 2320 58608
rect 2372 58596 2378 58608
rect 2590 58596 2596 58608
rect 2372 58568 2596 58596
rect 2372 58556 2378 58568
rect 2590 58556 2596 58568
rect 2648 58556 2654 58608
rect 3510 58556 3516 58608
rect 3568 58596 3574 58608
rect 3970 58596 3976 58608
rect 3568 58568 3976 58596
rect 3568 58556 3574 58568
rect 3970 58556 3976 58568
rect 4028 58556 4034 58608
rect 198 58488 204 58540
rect 256 58528 262 58540
rect 1397 58531 1455 58537
rect 1397 58528 1409 58531
rect 256 58500 1409 58528
rect 256 58488 262 58500
rect 1397 58497 1409 58500
rect 1443 58497 1455 58531
rect 1397 58491 1455 58497
rect 1946 58488 1952 58540
rect 2004 58528 2010 58540
rect 2682 58528 2688 58540
rect 2004 58500 2688 58528
rect 2004 58488 2010 58500
rect 2682 58488 2688 58500
rect 2740 58488 2746 58540
rect 3329 58531 3387 58537
rect 3329 58497 3341 58531
rect 3375 58528 3387 58531
rect 3694 58528 3700 58540
rect 3375 58500 3700 58528
rect 3375 58497 3387 58500
rect 3329 58491 3387 58497
rect 3694 58488 3700 58500
rect 3752 58488 3758 58540
rect 5074 58488 5080 58540
rect 5132 58528 5138 58540
rect 9585 58531 9643 58537
rect 9585 58528 9597 58531
rect 5132 58500 9597 58528
rect 5132 58488 5138 58500
rect 9585 58497 9597 58500
rect 9631 58497 9643 58531
rect 9585 58491 9643 58497
rect 2501 58463 2559 58469
rect 2501 58429 2513 58463
rect 2547 58460 2559 58463
rect 4154 58460 4160 58472
rect 2547 58432 4160 58460
rect 2547 58429 2559 58432
rect 2501 58423 2559 58429
rect 4154 58420 4160 58432
rect 4212 58420 4218 58472
rect 9309 58463 9367 58469
rect 9309 58429 9321 58463
rect 9355 58460 9367 58463
rect 9490 58460 9496 58472
rect 9355 58432 9496 58460
rect 9355 58429 9367 58432
rect 9309 58423 9367 58429
rect 9490 58420 9496 58432
rect 9548 58420 9554 58472
rect 3510 58392 3516 58404
rect 3471 58364 3516 58392
rect 3510 58352 3516 58364
rect 3568 58352 3574 58404
rect 1394 58284 1400 58336
rect 1452 58324 1458 58336
rect 1581 58327 1639 58333
rect 1581 58324 1593 58327
rect 1452 58296 1593 58324
rect 1452 58284 1458 58296
rect 1581 58293 1593 58296
rect 1627 58293 1639 58327
rect 1581 58287 1639 58293
rect 1104 58234 10856 58256
rect 1104 58182 2582 58234
rect 2634 58182 2646 58234
rect 2698 58182 2710 58234
rect 2762 58182 2774 58234
rect 2826 58182 2838 58234
rect 2890 58182 5846 58234
rect 5898 58182 5910 58234
rect 5962 58182 5974 58234
rect 6026 58182 6038 58234
rect 6090 58182 6102 58234
rect 6154 58182 9110 58234
rect 9162 58182 9174 58234
rect 9226 58182 9238 58234
rect 9290 58182 9302 58234
rect 9354 58182 9366 58234
rect 9418 58182 10856 58234
rect 1104 58160 10856 58182
rect 3510 58080 3516 58132
rect 3568 58120 3574 58132
rect 4154 58120 4160 58132
rect 3568 58092 4160 58120
rect 3568 58080 3574 58092
rect 4154 58080 4160 58092
rect 4212 58080 4218 58132
rect 2774 58012 2780 58064
rect 2832 58052 2838 58064
rect 3234 58052 3240 58064
rect 2832 58024 3240 58052
rect 2832 58012 2838 58024
rect 3234 58012 3240 58024
rect 3292 58012 3298 58064
rect 750 57876 756 57928
rect 808 57916 814 57928
rect 1397 57919 1455 57925
rect 1397 57916 1409 57919
rect 808 57888 1409 57916
rect 808 57876 814 57888
rect 1397 57885 1409 57888
rect 1443 57885 1455 57919
rect 1397 57879 1455 57885
rect 2133 57919 2191 57925
rect 2133 57885 2145 57919
rect 2179 57885 2191 57919
rect 2133 57879 2191 57885
rect 382 57808 388 57860
rect 440 57848 446 57860
rect 2148 57848 2176 57879
rect 440 57820 2176 57848
rect 440 57808 446 57820
rect 1578 57780 1584 57792
rect 1539 57752 1584 57780
rect 1578 57740 1584 57752
rect 1636 57740 1642 57792
rect 2317 57783 2375 57789
rect 2317 57749 2329 57783
rect 2363 57780 2375 57783
rect 2590 57780 2596 57792
rect 2363 57752 2596 57780
rect 2363 57749 2375 57752
rect 2317 57743 2375 57749
rect 2590 57740 2596 57752
rect 2648 57740 2654 57792
rect 1104 57690 10856 57712
rect 1104 57638 4214 57690
rect 4266 57638 4278 57690
rect 4330 57638 4342 57690
rect 4394 57638 4406 57690
rect 4458 57638 4470 57690
rect 4522 57638 7478 57690
rect 7530 57638 7542 57690
rect 7594 57638 7606 57690
rect 7658 57638 7670 57690
rect 7722 57638 7734 57690
rect 7786 57638 10856 57690
rect 1104 57616 10856 57638
rect 1762 57576 1768 57588
rect 1688 57548 1768 57576
rect 1688 57517 1716 57548
rect 1762 57536 1768 57548
rect 1820 57536 1826 57588
rect 1673 57511 1731 57517
rect 1673 57477 1685 57511
rect 1719 57477 1731 57511
rect 1673 57471 1731 57477
rect 1397 57443 1455 57449
rect 1397 57409 1409 57443
rect 1443 57409 1455 57443
rect 1397 57403 1455 57409
rect 1581 57443 1639 57449
rect 1581 57409 1593 57443
rect 1627 57409 1639 57443
rect 1581 57403 1639 57409
rect 1412 57372 1440 57403
rect 1320 57344 1440 57372
rect 1596 57372 1624 57403
rect 1762 57400 1768 57452
rect 1820 57449 1826 57452
rect 1820 57443 1875 57449
rect 1820 57409 1829 57443
rect 1863 57440 1875 57443
rect 2130 57440 2136 57452
rect 1863 57412 2136 57440
rect 1863 57409 1875 57412
rect 1820 57403 1875 57409
rect 1820 57400 1826 57403
rect 2130 57400 2136 57412
rect 2188 57400 2194 57452
rect 6546 57400 6552 57452
rect 6604 57440 6610 57452
rect 9585 57443 9643 57449
rect 9585 57440 9597 57443
rect 6604 57412 9597 57440
rect 6604 57400 6610 57412
rect 9585 57409 9597 57412
rect 9631 57409 9643 57443
rect 9585 57403 9643 57409
rect 2314 57372 2320 57384
rect 1596 57344 2320 57372
rect 1320 57236 1348 57344
rect 2314 57332 2320 57344
rect 2372 57332 2378 57384
rect 3050 57332 3056 57384
rect 3108 57372 3114 57384
rect 3234 57372 3240 57384
rect 3108 57344 3240 57372
rect 3108 57332 3114 57344
rect 3234 57332 3240 57344
rect 3292 57332 3298 57384
rect 9309 57375 9367 57381
rect 9309 57341 9321 57375
rect 9355 57372 9367 57375
rect 9490 57372 9496 57384
rect 9355 57344 9496 57372
rect 9355 57341 9367 57344
rect 9309 57335 9367 57341
rect 9490 57332 9496 57344
rect 9548 57332 9554 57384
rect 9950 57304 9956 57316
rect 1688 57276 9956 57304
rect 1688 57236 1716 57276
rect 9950 57264 9956 57276
rect 10008 57264 10014 57316
rect 1320 57208 1716 57236
rect 1949 57239 2007 57245
rect 1949 57205 1961 57239
rect 1995 57236 2007 57239
rect 2130 57236 2136 57248
rect 1995 57208 2136 57236
rect 1995 57205 2007 57208
rect 1949 57199 2007 57205
rect 2130 57196 2136 57208
rect 2188 57196 2194 57248
rect 1104 57146 10856 57168
rect 1104 57094 2582 57146
rect 2634 57094 2646 57146
rect 2698 57094 2710 57146
rect 2762 57094 2774 57146
rect 2826 57094 2838 57146
rect 2890 57094 5846 57146
rect 5898 57094 5910 57146
rect 5962 57094 5974 57146
rect 6026 57094 6038 57146
rect 6090 57094 6102 57146
rect 6154 57094 9110 57146
rect 9162 57094 9174 57146
rect 9226 57094 9238 57146
rect 9290 57094 9302 57146
rect 9354 57094 9366 57146
rect 9418 57094 10856 57146
rect 1104 57072 10856 57094
rect 842 56992 848 57044
rect 900 57032 906 57044
rect 2501 57035 2559 57041
rect 2501 57032 2513 57035
rect 900 57004 2513 57032
rect 900 56992 906 57004
rect 2501 57001 2513 57004
rect 2547 57001 2559 57035
rect 2501 56995 2559 57001
rect 1946 56964 1952 56976
rect 1907 56936 1952 56964
rect 1946 56924 1952 56936
rect 2004 56924 2010 56976
rect 8294 56896 8300 56908
rect 1412 56868 8300 56896
rect 1412 56837 1440 56868
rect 8294 56856 8300 56868
rect 8352 56856 8358 56908
rect 8478 56856 8484 56908
rect 8536 56896 8542 56908
rect 9585 56899 9643 56905
rect 9585 56896 9597 56899
rect 8536 56868 9597 56896
rect 8536 56856 8542 56868
rect 9585 56865 9597 56868
rect 9631 56865 9643 56899
rect 9585 56859 9643 56865
rect 1397 56831 1455 56837
rect 1397 56797 1409 56831
rect 1443 56797 1455 56831
rect 1670 56828 1676 56840
rect 1631 56800 1676 56828
rect 1397 56791 1455 56797
rect 1670 56788 1676 56800
rect 1728 56788 1734 56840
rect 1762 56788 1768 56840
rect 1820 56837 1826 56840
rect 1820 56828 1828 56837
rect 2314 56828 2320 56840
rect 1820 56800 2320 56828
rect 1820 56791 1828 56800
rect 1820 56788 1826 56791
rect 2314 56788 2320 56800
rect 2372 56788 2378 56840
rect 2685 56831 2743 56837
rect 2685 56797 2697 56831
rect 2731 56828 2743 56831
rect 3050 56828 3056 56840
rect 2731 56800 3056 56828
rect 2731 56797 2743 56800
rect 2685 56791 2743 56797
rect 3050 56788 3056 56800
rect 3108 56788 3114 56840
rect 9306 56828 9312 56840
rect 9267 56800 9312 56828
rect 9306 56788 9312 56800
rect 9364 56788 9370 56840
rect 1578 56760 1584 56772
rect 1491 56732 1584 56760
rect 1578 56720 1584 56732
rect 1636 56760 1642 56772
rect 2406 56760 2412 56772
rect 1636 56732 2412 56760
rect 1636 56720 1642 56732
rect 2406 56720 2412 56732
rect 2464 56720 2470 56772
rect 1104 56602 10856 56624
rect 1104 56550 4214 56602
rect 4266 56550 4278 56602
rect 4330 56550 4342 56602
rect 4394 56550 4406 56602
rect 4458 56550 4470 56602
rect 4522 56550 7478 56602
rect 7530 56550 7542 56602
rect 7594 56550 7606 56602
rect 7658 56550 7670 56602
rect 7722 56550 7734 56602
rect 7786 56550 10856 56602
rect 1104 56528 10856 56550
rect 1581 56491 1639 56497
rect 1581 56457 1593 56491
rect 1627 56488 1639 56491
rect 1670 56488 1676 56500
rect 1627 56460 1676 56488
rect 1627 56457 1639 56460
rect 1581 56451 1639 56457
rect 1670 56448 1676 56460
rect 1728 56448 1734 56500
rect 3602 56488 3608 56500
rect 3563 56460 3608 56488
rect 3602 56448 3608 56460
rect 3660 56448 3666 56500
rect 1762 56420 1768 56432
rect 1412 56392 1768 56420
rect 1412 56361 1440 56392
rect 1762 56380 1768 56392
rect 1820 56380 1826 56432
rect 1397 56355 1455 56361
rect 1397 56321 1409 56355
rect 1443 56321 1455 56355
rect 1397 56315 1455 56321
rect 1486 56312 1492 56364
rect 1544 56352 1550 56364
rect 1670 56352 1676 56364
rect 1544 56324 1676 56352
rect 1544 56312 1550 56324
rect 1670 56312 1676 56324
rect 1728 56312 1734 56364
rect 2133 56355 2191 56361
rect 2133 56321 2145 56355
rect 2179 56321 2191 56355
rect 2133 56315 2191 56321
rect 2869 56355 2927 56361
rect 2869 56321 2881 56355
rect 2915 56321 2927 56355
rect 2869 56315 2927 56321
rect 1210 56244 1216 56296
rect 1268 56284 1274 56296
rect 2148 56284 2176 56315
rect 1268 56256 2176 56284
rect 2884 56284 2912 56315
rect 3602 56312 3608 56364
rect 3660 56352 3666 56364
rect 3789 56355 3847 56361
rect 3789 56352 3801 56355
rect 3660 56324 3801 56352
rect 3660 56312 3666 56324
rect 3789 56321 3801 56324
rect 3835 56321 3847 56355
rect 10134 56352 10140 56364
rect 10095 56324 10140 56352
rect 3789 56315 3847 56321
rect 10134 56312 10140 56324
rect 10192 56312 10198 56364
rect 6362 56284 6368 56296
rect 2884 56256 6368 56284
rect 1268 56244 1274 56256
rect 6362 56244 6368 56256
rect 6420 56244 6426 56296
rect 2682 56176 2688 56228
rect 2740 56216 2746 56228
rect 3053 56219 3111 56225
rect 3053 56216 3065 56219
rect 2740 56188 3065 56216
rect 2740 56176 2746 56188
rect 3053 56185 3065 56188
rect 3099 56185 3111 56219
rect 3053 56179 3111 56185
rect 2314 56148 2320 56160
rect 2275 56120 2320 56148
rect 2314 56108 2320 56120
rect 2372 56108 2378 56160
rect 4982 56108 4988 56160
rect 5040 56148 5046 56160
rect 5442 56148 5448 56160
rect 5040 56120 5448 56148
rect 5040 56108 5046 56120
rect 5442 56108 5448 56120
rect 5500 56108 5506 56160
rect 6178 56108 6184 56160
rect 6236 56148 6242 56160
rect 9953 56151 10011 56157
rect 9953 56148 9965 56151
rect 6236 56120 9965 56148
rect 6236 56108 6242 56120
rect 9953 56117 9965 56120
rect 9999 56117 10011 56151
rect 9953 56111 10011 56117
rect 1104 56058 10856 56080
rect 1104 56006 2582 56058
rect 2634 56006 2646 56058
rect 2698 56006 2710 56058
rect 2762 56006 2774 56058
rect 2826 56006 2838 56058
rect 2890 56006 5846 56058
rect 5898 56006 5910 56058
rect 5962 56006 5974 56058
rect 6026 56006 6038 56058
rect 6090 56006 6102 56058
rect 6154 56006 9110 56058
rect 9162 56006 9174 56058
rect 9226 56006 9238 56058
rect 9290 56006 9302 56058
rect 9354 56006 9366 56058
rect 9418 56006 10856 56058
rect 1104 55984 10856 56006
rect 4982 55836 4988 55888
rect 5040 55876 5046 55888
rect 5350 55876 5356 55888
rect 5040 55848 5356 55876
rect 5040 55836 5046 55848
rect 5350 55836 5356 55848
rect 5408 55836 5414 55888
rect 3234 55808 3240 55820
rect 3068 55780 3240 55808
rect 842 55700 848 55752
rect 900 55740 906 55752
rect 1397 55743 1455 55749
rect 1397 55740 1409 55743
rect 900 55712 1409 55740
rect 900 55700 906 55712
rect 1397 55709 1409 55712
rect 1443 55709 1455 55743
rect 1397 55703 1455 55709
rect 2133 55743 2191 55749
rect 2133 55709 2145 55743
rect 2179 55740 2191 55743
rect 2179 55712 2774 55740
rect 2179 55709 2191 55712
rect 2133 55703 2191 55709
rect 2746 55672 2774 55712
rect 2866 55700 2872 55752
rect 2924 55740 2930 55752
rect 3068 55749 3096 55780
rect 3234 55768 3240 55780
rect 3292 55808 3298 55820
rect 3292 55780 4016 55808
rect 3292 55768 3298 55780
rect 3053 55743 3111 55749
rect 2924 55712 2969 55740
rect 2924 55700 2930 55712
rect 3053 55709 3065 55743
rect 3099 55709 3111 55743
rect 3053 55703 3111 55709
rect 3510 55700 3516 55752
rect 3568 55740 3574 55752
rect 3988 55749 4016 55780
rect 3789 55743 3847 55749
rect 3789 55740 3801 55743
rect 3568 55712 3801 55740
rect 3568 55700 3574 55712
rect 3789 55709 3801 55712
rect 3835 55709 3847 55743
rect 3789 55703 3847 55709
rect 3973 55743 4031 55749
rect 3973 55709 3985 55743
rect 4019 55740 4031 55743
rect 4154 55740 4160 55752
rect 4019 55712 4160 55740
rect 4019 55709 4031 55712
rect 3973 55703 4031 55709
rect 4154 55700 4160 55712
rect 4212 55700 4218 55752
rect 9582 55700 9588 55752
rect 9640 55740 9646 55752
rect 10137 55743 10195 55749
rect 10137 55740 10149 55743
rect 9640 55712 10149 55740
rect 9640 55700 9646 55712
rect 10137 55709 10149 55712
rect 10183 55709 10195 55743
rect 10137 55703 10195 55709
rect 6454 55672 6460 55684
rect 2746 55644 6460 55672
rect 6454 55632 6460 55644
rect 6512 55632 6518 55684
rect 1578 55604 1584 55616
rect 1539 55576 1584 55604
rect 1578 55564 1584 55576
rect 1636 55564 1642 55616
rect 2314 55604 2320 55616
rect 2275 55576 2320 55604
rect 2314 55564 2320 55576
rect 2372 55564 2378 55616
rect 3234 55604 3240 55616
rect 3195 55576 3240 55604
rect 3234 55564 3240 55576
rect 3292 55564 3298 55616
rect 4157 55607 4215 55613
rect 4157 55573 4169 55607
rect 4203 55604 4215 55607
rect 6822 55604 6828 55616
rect 4203 55576 6828 55604
rect 4203 55573 4215 55576
rect 4157 55567 4215 55573
rect 6822 55564 6828 55576
rect 6880 55564 6886 55616
rect 8294 55564 8300 55616
rect 8352 55604 8358 55616
rect 9953 55607 10011 55613
rect 9953 55604 9965 55607
rect 8352 55576 9965 55604
rect 8352 55564 8358 55576
rect 9953 55573 9965 55576
rect 9999 55573 10011 55607
rect 9953 55567 10011 55573
rect 566 55536 572 55548
rect 400 55508 572 55536
rect 400 52816 428 55508
rect 566 55496 572 55508
rect 624 55496 630 55548
rect 1104 55514 10856 55536
rect 1104 55462 4214 55514
rect 4266 55462 4278 55514
rect 4330 55462 4342 55514
rect 4394 55462 4406 55514
rect 4458 55462 4470 55514
rect 4522 55462 7478 55514
rect 7530 55462 7542 55514
rect 7594 55462 7606 55514
rect 7658 55462 7670 55514
rect 7722 55462 7734 55514
rect 7786 55462 10856 55514
rect 1104 55440 10856 55462
rect 2777 55403 2835 55409
rect 2777 55369 2789 55403
rect 2823 55400 2835 55403
rect 3050 55400 3056 55412
rect 2823 55372 3056 55400
rect 2823 55369 2835 55372
rect 2777 55363 2835 55369
rect 3050 55360 3056 55372
rect 3108 55360 3114 55412
rect 3234 55360 3240 55412
rect 3292 55360 3298 55412
rect 3602 55400 3608 55412
rect 3563 55372 3608 55400
rect 3602 55360 3608 55372
rect 3660 55360 3666 55412
rect 4433 55403 4491 55409
rect 4433 55369 4445 55403
rect 4479 55400 4491 55403
rect 10134 55400 10140 55412
rect 4479 55372 10140 55400
rect 4479 55369 4491 55372
rect 4433 55363 4491 55369
rect 10134 55360 10140 55372
rect 10192 55360 10198 55412
rect 1302 55292 1308 55344
rect 1360 55332 1366 55344
rect 3252 55332 3280 55360
rect 1360 55304 2544 55332
rect 3252 55304 10180 55332
rect 1360 55292 1366 55304
rect 1397 55267 1455 55273
rect 1397 55233 1409 55267
rect 1443 55264 1455 55267
rect 1762 55264 1768 55276
rect 1443 55236 1768 55264
rect 1443 55233 1455 55236
rect 1397 55227 1455 55233
rect 1762 55224 1768 55236
rect 1820 55224 1826 55276
rect 2409 55199 2467 55205
rect 2409 55165 2421 55199
rect 2455 55165 2467 55199
rect 2516 55196 2544 55304
rect 2593 55267 2651 55273
rect 2593 55233 2605 55267
rect 2639 55264 2651 55267
rect 3421 55267 3479 55273
rect 3421 55264 3433 55267
rect 2639 55262 3096 55264
rect 3160 55262 3433 55264
rect 2639 55236 3433 55262
rect 2639 55233 2651 55236
rect 3068 55234 3188 55236
rect 2593 55227 2651 55233
rect 3421 55233 3433 55236
rect 3467 55264 3479 55267
rect 3602 55264 3608 55276
rect 3467 55236 3608 55264
rect 3467 55233 3479 55236
rect 3421 55227 3479 55233
rect 3602 55224 3608 55236
rect 3660 55224 3666 55276
rect 10152 55273 10180 55304
rect 4249 55267 4307 55273
rect 4249 55233 4261 55267
rect 4295 55264 4307 55267
rect 10137 55267 10195 55273
rect 4295 55236 4384 55264
rect 4295 55233 4307 55236
rect 4249 55227 4307 55233
rect 4356 55208 4384 55236
rect 10137 55233 10149 55267
rect 10183 55233 10195 55267
rect 10137 55227 10195 55233
rect 3237 55199 3295 55205
rect 2516 55168 3188 55196
rect 2409 55159 2467 55165
rect 1302 55088 1308 55140
rect 1360 55128 1366 55140
rect 1360 55100 1900 55128
rect 1360 55088 1366 55100
rect 658 55020 664 55072
rect 716 55060 722 55072
rect 1118 55060 1124 55072
rect 716 55032 1124 55060
rect 716 55020 722 55032
rect 1118 55020 1124 55032
rect 1176 55020 1182 55072
rect 1486 55020 1492 55072
rect 1544 55060 1550 55072
rect 1581 55063 1639 55069
rect 1581 55060 1593 55063
rect 1544 55032 1593 55060
rect 1544 55020 1550 55032
rect 1581 55029 1593 55032
rect 1627 55029 1639 55063
rect 1872 55060 1900 55100
rect 2424 55060 2452 55159
rect 3160 55140 3188 55168
rect 3237 55165 3249 55199
rect 3283 55196 3295 55199
rect 3510 55196 3516 55208
rect 3283 55168 3516 55196
rect 3283 55165 3295 55168
rect 3237 55159 3295 55165
rect 3510 55156 3516 55168
rect 3568 55156 3574 55208
rect 4065 55199 4123 55205
rect 4065 55165 4077 55199
rect 4111 55165 4123 55199
rect 4065 55159 4123 55165
rect 3142 55088 3148 55140
rect 3200 55088 3206 55140
rect 4080 55060 4108 55159
rect 4338 55156 4344 55208
rect 4396 55156 4402 55208
rect 1872 55032 4108 55060
rect 1581 55023 1639 55029
rect 9858 55020 9864 55072
rect 9916 55060 9922 55072
rect 9953 55063 10011 55069
rect 9953 55060 9965 55063
rect 9916 55032 9965 55060
rect 9916 55020 9922 55032
rect 9953 55029 9965 55032
rect 9999 55029 10011 55063
rect 9953 55023 10011 55029
rect 1104 54970 10856 54992
rect 1104 54918 2582 54970
rect 2634 54918 2646 54970
rect 2698 54918 2710 54970
rect 2762 54918 2774 54970
rect 2826 54918 2838 54970
rect 2890 54918 5846 54970
rect 5898 54918 5910 54970
rect 5962 54918 5974 54970
rect 6026 54918 6038 54970
rect 6090 54918 6102 54970
rect 6154 54918 9110 54970
rect 9162 54918 9174 54970
rect 9226 54918 9238 54970
rect 9290 54918 9302 54970
rect 9354 54918 9366 54970
rect 9418 54918 10856 54970
rect 1104 54896 10856 54918
rect 3510 54816 3516 54868
rect 3568 54856 3574 54868
rect 4062 54856 4068 54868
rect 3568 54828 4068 54856
rect 3568 54816 3574 54828
rect 4062 54816 4068 54828
rect 4120 54816 4126 54868
rect 1670 54788 1676 54800
rect 1596 54760 1676 54788
rect 1397 54655 1455 54661
rect 1397 54621 1409 54655
rect 1443 54621 1455 54655
rect 1596 54652 1624 54760
rect 1670 54748 1676 54760
rect 1728 54748 1734 54800
rect 1949 54791 2007 54797
rect 1949 54757 1961 54791
rect 1995 54788 2007 54791
rect 2406 54788 2412 54800
rect 1995 54760 2412 54788
rect 1995 54757 2007 54760
rect 1949 54751 2007 54757
rect 2406 54748 2412 54760
rect 2464 54748 2470 54800
rect 1674 54655 1732 54661
rect 1674 54652 1686 54655
rect 1596 54624 1686 54652
rect 1397 54615 1455 54621
rect 1674 54621 1686 54624
rect 1720 54621 1732 54655
rect 1674 54615 1732 54621
rect 1811 54655 1869 54661
rect 1811 54621 1823 54655
rect 1857 54652 1869 54655
rect 2314 54652 2320 54664
rect 1857 54624 2320 54652
rect 1857 54621 1869 54624
rect 1811 54615 1869 54621
rect 1412 54516 1440 54615
rect 2314 54612 2320 54624
rect 2372 54612 2378 54664
rect 2501 54655 2559 54661
rect 2501 54621 2513 54655
rect 2547 54652 2559 54655
rect 6270 54652 6276 54664
rect 2547 54624 6276 54652
rect 2547 54621 2559 54624
rect 2501 54615 2559 54621
rect 6270 54612 6276 54624
rect 6328 54612 6334 54664
rect 6822 54612 6828 54664
rect 6880 54652 6886 54664
rect 9493 54655 9551 54661
rect 9493 54652 9505 54655
rect 6880 54624 9505 54652
rect 6880 54612 6886 54624
rect 9493 54621 9505 54624
rect 9539 54621 9551 54655
rect 10134 54652 10140 54664
rect 10095 54624 10140 54652
rect 9493 54615 9551 54621
rect 10134 54612 10140 54624
rect 10192 54612 10198 54664
rect 1578 54584 1584 54596
rect 1539 54556 1584 54584
rect 1578 54544 1584 54556
rect 1636 54544 1642 54596
rect 6178 54584 6184 54596
rect 1688 54556 6184 54584
rect 1688 54516 1716 54556
rect 6178 54544 6184 54556
rect 6236 54544 6242 54596
rect 1412 54488 1716 54516
rect 2685 54519 2743 54525
rect 2685 54485 2697 54519
rect 2731 54516 2743 54519
rect 2774 54516 2780 54528
rect 2731 54488 2780 54516
rect 2731 54485 2743 54488
rect 2685 54479 2743 54485
rect 2774 54476 2780 54488
rect 2832 54476 2838 54528
rect 9309 54519 9367 54525
rect 9309 54485 9321 54519
rect 9355 54516 9367 54519
rect 9674 54516 9680 54528
rect 9355 54488 9680 54516
rect 9355 54485 9367 54488
rect 9309 54479 9367 54485
rect 9674 54476 9680 54488
rect 9732 54476 9738 54528
rect 9950 54516 9956 54528
rect 9911 54488 9956 54516
rect 9950 54476 9956 54488
rect 10008 54476 10014 54528
rect 1104 54426 10856 54448
rect 1104 54374 4214 54426
rect 4266 54374 4278 54426
rect 4330 54374 4342 54426
rect 4394 54374 4406 54426
rect 4458 54374 4470 54426
rect 4522 54374 7478 54426
rect 7530 54374 7542 54426
rect 7594 54374 7606 54426
rect 7658 54374 7670 54426
rect 7722 54374 7734 54426
rect 7786 54374 10856 54426
rect 1104 54352 10856 54374
rect 1394 54272 1400 54324
rect 1452 54312 1458 54324
rect 1670 54312 1676 54324
rect 1452 54284 1676 54312
rect 1452 54272 1458 54284
rect 1670 54272 1676 54284
rect 1728 54272 1734 54324
rect 8294 54244 8300 54256
rect 1412 54216 8300 54244
rect 1412 54185 1440 54216
rect 8294 54204 8300 54216
rect 8352 54204 8358 54256
rect 1397 54179 1455 54185
rect 1397 54145 1409 54179
rect 1443 54145 1455 54179
rect 1578 54176 1584 54188
rect 1539 54148 1584 54176
rect 1397 54139 1455 54145
rect 1578 54136 1584 54148
rect 1636 54136 1642 54188
rect 1673 54179 1731 54185
rect 1673 54145 1685 54179
rect 1719 54145 1731 54179
rect 1673 54139 1731 54145
rect 1770 54179 1828 54185
rect 1770 54145 1782 54179
rect 1816 54176 1828 54179
rect 2501 54179 2559 54185
rect 1816 54148 2176 54176
rect 1816 54145 1828 54148
rect 1770 54139 1828 54145
rect 566 54068 572 54120
rect 624 54108 630 54120
rect 1596 54108 1624 54136
rect 624 54080 1624 54108
rect 1688 54108 1716 54139
rect 2038 54108 2044 54120
rect 1688 54080 2044 54108
rect 624 54068 630 54080
rect 2038 54068 2044 54080
rect 2096 54068 2102 54120
rect 2148 54108 2176 54148
rect 2501 54145 2513 54179
rect 2547 54145 2559 54179
rect 9858 54176 9864 54188
rect 9819 54148 9864 54176
rect 2501 54139 2559 54145
rect 2314 54108 2320 54120
rect 2148 54080 2320 54108
rect 2314 54068 2320 54080
rect 2372 54068 2378 54120
rect 1302 54000 1308 54052
rect 1360 54040 1366 54052
rect 2516 54040 2544 54139
rect 9858 54136 9864 54148
rect 9916 54136 9922 54188
rect 10042 54040 10048 54052
rect 1360 54012 2544 54040
rect 10003 54012 10048 54040
rect 1360 54000 1366 54012
rect 10042 54000 10048 54012
rect 10100 54000 10106 54052
rect 1762 53932 1768 53984
rect 1820 53972 1826 53984
rect 1949 53975 2007 53981
rect 1949 53972 1961 53975
rect 1820 53944 1961 53972
rect 1820 53932 1826 53944
rect 1949 53941 1961 53944
rect 1995 53941 2007 53975
rect 1949 53935 2007 53941
rect 2038 53932 2044 53984
rect 2096 53972 2102 53984
rect 2685 53975 2743 53981
rect 2685 53972 2697 53975
rect 2096 53944 2697 53972
rect 2096 53932 2102 53944
rect 2685 53941 2697 53944
rect 2731 53941 2743 53975
rect 2685 53935 2743 53941
rect 1104 53882 10856 53904
rect 1104 53830 2582 53882
rect 2634 53830 2646 53882
rect 2698 53830 2710 53882
rect 2762 53830 2774 53882
rect 2826 53830 2838 53882
rect 2890 53830 5846 53882
rect 5898 53830 5910 53882
rect 5962 53830 5974 53882
rect 6026 53830 6038 53882
rect 6090 53830 6102 53882
rect 6154 53830 9110 53882
rect 9162 53830 9174 53882
rect 9226 53830 9238 53882
rect 9290 53830 9302 53882
rect 9354 53830 9366 53882
rect 9418 53830 10856 53882
rect 1104 53808 10856 53830
rect 2314 53592 2320 53644
rect 2372 53632 2378 53644
rect 2590 53632 2596 53644
rect 2372 53604 2596 53632
rect 2372 53592 2378 53604
rect 2590 53592 2596 53604
rect 2648 53592 2654 53644
rect 1397 53567 1455 53573
rect 1397 53533 1409 53567
rect 1443 53533 1455 53567
rect 1397 53527 1455 53533
rect 2133 53567 2191 53573
rect 2133 53533 2145 53567
rect 2179 53564 2191 53567
rect 4614 53564 4620 53576
rect 2179 53536 4620 53564
rect 2179 53533 2191 53536
rect 2133 53527 2191 53533
rect 1412 53496 1440 53527
rect 4614 53524 4620 53536
rect 4672 53524 4678 53576
rect 9674 53524 9680 53576
rect 9732 53564 9738 53576
rect 9861 53567 9919 53573
rect 9861 53564 9873 53567
rect 9732 53536 9873 53564
rect 9732 53524 9738 53536
rect 9861 53533 9873 53536
rect 9907 53533 9919 53567
rect 9861 53527 9919 53533
rect 5350 53496 5356 53508
rect 1412 53468 5356 53496
rect 5350 53456 5356 53468
rect 5408 53456 5414 53508
rect 1394 53388 1400 53440
rect 1452 53428 1458 53440
rect 1581 53431 1639 53437
rect 1581 53428 1593 53431
rect 1452 53400 1593 53428
rect 1452 53388 1458 53400
rect 1581 53397 1593 53400
rect 1627 53397 1639 53431
rect 2314 53428 2320 53440
rect 2275 53400 2320 53428
rect 1581 53391 1639 53397
rect 2314 53388 2320 53400
rect 2372 53388 2378 53440
rect 10042 53428 10048 53440
rect 10003 53400 10048 53428
rect 10042 53388 10048 53400
rect 10100 53388 10106 53440
rect 1104 53338 10856 53360
rect 1104 53286 4214 53338
rect 4266 53286 4278 53338
rect 4330 53286 4342 53338
rect 4394 53286 4406 53338
rect 4458 53286 4470 53338
rect 4522 53286 7478 53338
rect 7530 53286 7542 53338
rect 7594 53286 7606 53338
rect 7658 53286 7670 53338
rect 7722 53286 7734 53338
rect 7786 53286 10856 53338
rect 1104 53264 10856 53286
rect 2038 53184 2044 53236
rect 2096 53224 2102 53236
rect 2222 53224 2228 53236
rect 2096 53196 2228 53224
rect 2096 53184 2102 53196
rect 2222 53184 2228 53196
rect 2280 53184 2286 53236
rect 4706 53116 4712 53168
rect 4764 53156 4770 53168
rect 6822 53156 6828 53168
rect 4764 53128 6828 53156
rect 4764 53116 4770 53128
rect 6822 53116 6828 53128
rect 6880 53116 6886 53168
rect 658 53048 664 53100
rect 716 53088 722 53100
rect 1397 53091 1455 53097
rect 1397 53088 1409 53091
rect 716 53060 1409 53088
rect 716 53048 722 53060
rect 1397 53057 1409 53060
rect 1443 53057 1455 53091
rect 1397 53051 1455 53057
rect 2222 53048 2228 53100
rect 2280 53088 2286 53100
rect 2498 53088 2504 53100
rect 2280 53060 2504 53088
rect 2280 53048 2286 53060
rect 2498 53048 2504 53060
rect 2556 53048 2562 53100
rect 9861 53091 9919 53097
rect 9861 53057 9873 53091
rect 9907 53088 9919 53091
rect 9950 53088 9956 53100
rect 9907 53060 9956 53088
rect 9907 53057 9919 53060
rect 9861 53051 9919 53057
rect 9950 53048 9956 53060
rect 10008 53048 10014 53100
rect 1578 52884 1584 52896
rect 1539 52856 1584 52884
rect 1578 52844 1584 52856
rect 1636 52844 1642 52896
rect 2130 52844 2136 52896
rect 2188 52884 2194 52896
rect 2498 52884 2504 52896
rect 2188 52856 2504 52884
rect 2188 52844 2194 52856
rect 2498 52844 2504 52856
rect 2556 52844 2562 52896
rect 10042 52884 10048 52896
rect 10003 52856 10048 52884
rect 10042 52844 10048 52856
rect 10100 52844 10106 52896
rect 308 52788 428 52816
rect 1104 52794 10856 52816
rect 308 52476 336 52788
rect 1104 52742 2582 52794
rect 2634 52742 2646 52794
rect 2698 52742 2710 52794
rect 2762 52742 2774 52794
rect 2826 52742 2838 52794
rect 2890 52742 5846 52794
rect 5898 52742 5910 52794
rect 5962 52742 5974 52794
rect 6026 52742 6038 52794
rect 6090 52742 6102 52794
rect 6154 52742 9110 52794
rect 9162 52742 9174 52794
rect 9226 52742 9238 52794
rect 9290 52742 9302 52794
rect 9354 52742 9366 52794
rect 9418 52742 10856 52794
rect 1104 52720 10856 52742
rect 2133 52683 2191 52689
rect 2133 52649 2145 52683
rect 2179 52680 2191 52683
rect 4154 52680 4160 52692
rect 2179 52652 4160 52680
rect 2179 52649 2191 52652
rect 2133 52643 2191 52649
rect 4154 52640 4160 52652
rect 4212 52640 4218 52692
rect 5350 52544 5356 52556
rect 1412 52516 5356 52544
rect 474 52476 480 52488
rect 308 52448 480 52476
rect 474 52436 480 52448
rect 532 52436 538 52488
rect 1412 52485 1440 52516
rect 5350 52504 5356 52516
rect 5408 52504 5414 52556
rect 1397 52479 1455 52485
rect 1397 52445 1409 52479
rect 1443 52445 1455 52479
rect 2314 52476 2320 52488
rect 2275 52448 2320 52476
rect 1397 52439 1455 52445
rect 2314 52436 2320 52448
rect 2372 52436 2378 52488
rect 1486 52300 1492 52352
rect 1544 52340 1550 52352
rect 1581 52343 1639 52349
rect 1581 52340 1593 52343
rect 1544 52312 1593 52340
rect 1544 52300 1550 52312
rect 1581 52309 1593 52312
rect 1627 52309 1639 52343
rect 1581 52303 1639 52309
rect 1104 52250 10856 52272
rect 1104 52198 4214 52250
rect 4266 52198 4278 52250
rect 4330 52198 4342 52250
rect 4394 52198 4406 52250
rect 4458 52198 4470 52250
rect 4522 52198 7478 52250
rect 7530 52198 7542 52250
rect 7594 52198 7606 52250
rect 7658 52198 7670 52250
rect 7722 52198 7734 52250
rect 7786 52198 10856 52250
rect 1104 52176 10856 52198
rect 1578 52096 1584 52148
rect 1636 52136 1642 52148
rect 1636 52108 1716 52136
rect 1636 52096 1642 52108
rect 1394 52000 1400 52012
rect 1355 51972 1400 52000
rect 1394 51960 1400 51972
rect 1452 51960 1458 52012
rect 1688 52000 1716 52108
rect 2866 52096 2872 52148
rect 2924 52136 2930 52148
rect 3053 52139 3111 52145
rect 3053 52136 3065 52139
rect 2924 52108 3065 52136
rect 2924 52096 2930 52108
rect 3053 52105 3065 52108
rect 3099 52105 3111 52139
rect 3053 52099 3111 52105
rect 1596 51972 1716 52000
rect 2133 52003 2191 52009
rect 1596 51873 1624 51972
rect 2133 51969 2145 52003
rect 2179 52000 2191 52003
rect 2869 52003 2927 52009
rect 2179 51972 2774 52000
rect 2179 51969 2191 51972
rect 2133 51963 2191 51969
rect 2746 51932 2774 51972
rect 2869 51969 2881 52003
rect 2915 52000 2927 52003
rect 5350 52000 5356 52012
rect 2915 51972 5356 52000
rect 2915 51969 2927 51972
rect 2869 51963 2927 51969
rect 5350 51960 5356 51972
rect 5408 51960 5414 52012
rect 9858 52000 9864 52012
rect 9819 51972 9864 52000
rect 9858 51960 9864 51972
rect 9916 51960 9922 52012
rect 6914 51932 6920 51944
rect 2746 51904 6920 51932
rect 6914 51892 6920 51904
rect 6972 51892 6978 51944
rect 1581 51867 1639 51873
rect 1581 51833 1593 51867
rect 1627 51833 1639 51867
rect 1581 51827 1639 51833
rect 1670 51756 1676 51808
rect 1728 51796 1734 51808
rect 2317 51799 2375 51805
rect 2317 51796 2329 51799
rect 1728 51768 2329 51796
rect 1728 51756 1734 51768
rect 2317 51765 2329 51768
rect 2363 51765 2375 51799
rect 10042 51796 10048 51808
rect 10003 51768 10048 51796
rect 2317 51759 2375 51765
rect 10042 51756 10048 51768
rect 10100 51756 10106 51808
rect 1104 51706 10856 51728
rect 1104 51654 2582 51706
rect 2634 51654 2646 51706
rect 2698 51654 2710 51706
rect 2762 51654 2774 51706
rect 2826 51654 2838 51706
rect 2890 51654 5846 51706
rect 5898 51654 5910 51706
rect 5962 51654 5974 51706
rect 6026 51654 6038 51706
rect 6090 51654 6102 51706
rect 6154 51654 9110 51706
rect 9162 51654 9174 51706
rect 9226 51654 9238 51706
rect 9290 51654 9302 51706
rect 9354 51654 9366 51706
rect 9418 51654 10856 51706
rect 1104 51632 10856 51654
rect 2314 51552 2320 51604
rect 2372 51592 2378 51604
rect 2501 51595 2559 51601
rect 2501 51592 2513 51595
rect 2372 51564 2513 51592
rect 2372 51552 2378 51564
rect 2501 51561 2513 51564
rect 2547 51561 2559 51595
rect 2958 51592 2964 51604
rect 2919 51564 2964 51592
rect 2501 51555 2559 51561
rect 2958 51552 2964 51564
rect 3016 51552 3022 51604
rect 1302 51484 1308 51536
rect 1360 51524 1366 51536
rect 1670 51524 1676 51536
rect 1360 51496 1676 51524
rect 1360 51484 1366 51496
rect 1670 51484 1676 51496
rect 1728 51484 1734 51536
rect 3602 51456 3608 51468
rect 2976 51428 3608 51456
rect 1397 51391 1455 51397
rect 1397 51357 1409 51391
rect 1443 51388 1455 51391
rect 2225 51391 2283 51397
rect 1443 51360 2084 51388
rect 1443 51357 1455 51360
rect 1397 51351 1455 51357
rect 566 51212 572 51264
rect 624 51252 630 51264
rect 1578 51252 1584 51264
rect 624 51224 1072 51252
rect 1539 51224 1584 51252
rect 624 51212 630 51224
rect 106 51076 112 51128
rect 164 51116 170 51128
rect 566 51116 572 51128
rect 164 51088 572 51116
rect 164 51076 170 51088
rect 566 51076 572 51088
rect 624 51076 630 51128
rect 1044 50980 1072 51224
rect 1578 51212 1584 51224
rect 1636 51212 1642 51264
rect 2056 51252 2084 51360
rect 2225 51357 2237 51391
rect 2271 51357 2283 51391
rect 2225 51351 2283 51357
rect 2317 51391 2375 51397
rect 2317 51357 2329 51391
rect 2363 51388 2375 51391
rect 2590 51388 2596 51400
rect 2363 51360 2596 51388
rect 2363 51357 2375 51360
rect 2317 51351 2375 51357
rect 2240 51320 2268 51351
rect 2590 51348 2596 51360
rect 2648 51388 2654 51400
rect 2976 51388 3004 51428
rect 3602 51416 3608 51428
rect 3660 51416 3666 51468
rect 3142 51388 3148 51400
rect 2648 51360 3004 51388
rect 3103 51360 3148 51388
rect 2648 51348 2654 51360
rect 3142 51348 3148 51360
rect 3200 51348 3206 51400
rect 9674 51348 9680 51400
rect 9732 51388 9738 51400
rect 9861 51391 9919 51397
rect 9861 51388 9873 51391
rect 9732 51360 9873 51388
rect 9732 51348 9738 51360
rect 9861 51357 9873 51360
rect 9907 51357 9919 51391
rect 9861 51351 9919 51357
rect 2774 51320 2780 51332
rect 2240 51292 2780 51320
rect 2774 51280 2780 51292
rect 2832 51280 2838 51332
rect 6638 51252 6644 51264
rect 2056 51224 6644 51252
rect 6638 51212 6644 51224
rect 6696 51212 6702 51264
rect 10042 51252 10048 51264
rect 10003 51224 10048 51252
rect 10042 51212 10048 51224
rect 10100 51212 10106 51264
rect 1104 51162 10856 51184
rect 1104 51110 4214 51162
rect 4266 51110 4278 51162
rect 4330 51110 4342 51162
rect 4394 51110 4406 51162
rect 4458 51110 4470 51162
rect 4522 51110 7478 51162
rect 7530 51110 7542 51162
rect 7594 51110 7606 51162
rect 7658 51110 7670 51162
rect 7722 51110 7734 51162
rect 7786 51110 10856 51162
rect 1104 51088 10856 51110
rect 1118 51008 1124 51060
rect 1176 51048 1182 51060
rect 1176 51020 1717 51048
rect 1176 51008 1182 51020
rect 1689 50989 1717 51020
rect 2130 51008 2136 51060
rect 2188 51048 2194 51060
rect 2314 51048 2320 51060
rect 2188 51020 2320 51048
rect 2188 51008 2194 51020
rect 2314 51008 2320 51020
rect 2372 51008 2378 51060
rect 2869 51051 2927 51057
rect 2869 51017 2881 51051
rect 2915 51048 2927 51051
rect 3142 51048 3148 51060
rect 2915 51020 3148 51048
rect 2915 51017 2927 51020
rect 2869 51011 2927 51017
rect 3142 51008 3148 51020
rect 3200 51008 3206 51060
rect 5074 51048 5080 51060
rect 3252 51020 5080 51048
rect 1581 50983 1639 50989
rect 1581 50980 1593 50983
rect 1044 50952 1593 50980
rect 382 50464 388 50516
rect 440 50504 446 50516
rect 1044 50504 1072 50952
rect 1581 50949 1593 50952
rect 1627 50949 1639 50983
rect 1581 50943 1639 50949
rect 1669 50983 1727 50989
rect 1669 50949 1681 50983
rect 1715 50949 1727 50983
rect 3252 50980 3280 51020
rect 5074 51008 5080 51020
rect 5132 51008 5138 51060
rect 5166 51008 5172 51060
rect 5224 51008 5230 51060
rect 9858 51008 9864 51060
rect 9916 51048 9922 51060
rect 9953 51051 10011 51057
rect 9953 51048 9965 51051
rect 9916 51020 9965 51048
rect 9916 51008 9922 51020
rect 9953 51017 9965 51020
rect 9999 51017 10011 51051
rect 9953 51011 10011 51017
rect 5184 50980 5212 51008
rect 1669 50943 1727 50949
rect 2056 50952 3280 50980
rect 5000 50952 5212 50980
rect 9646 50952 10180 50980
rect 1397 50915 1455 50921
rect 1397 50881 1409 50915
rect 1443 50881 1455 50915
rect 1397 50875 1455 50881
rect 1412 50844 1440 50875
rect 1762 50872 1768 50924
rect 1820 50912 1826 50924
rect 1820 50884 1865 50912
rect 1820 50872 1826 50884
rect 2056 50844 2084 50952
rect 2130 50872 2136 50924
rect 2188 50872 2194 50924
rect 2685 50915 2743 50921
rect 2685 50912 2697 50915
rect 2608 50884 2697 50912
rect 1412 50816 2084 50844
rect 1118 50736 1124 50788
rect 1176 50776 1182 50788
rect 1486 50776 1492 50788
rect 1176 50748 1492 50776
rect 1176 50736 1182 50748
rect 1486 50736 1492 50748
rect 1544 50736 1550 50788
rect 2148 50776 2176 50872
rect 2608 50856 2636 50884
rect 2685 50881 2697 50884
rect 2731 50881 2743 50915
rect 2685 50875 2743 50881
rect 3513 50915 3571 50921
rect 3513 50881 3525 50915
rect 3559 50912 3571 50915
rect 4154 50912 4160 50924
rect 3559 50884 4160 50912
rect 3559 50881 3571 50884
rect 3513 50875 3571 50881
rect 4154 50872 4160 50884
rect 4212 50912 4218 50924
rect 4798 50912 4804 50924
rect 4212 50884 4804 50912
rect 4212 50872 4218 50884
rect 4798 50872 4804 50884
rect 4856 50872 4862 50924
rect 5000 50856 5028 50952
rect 5350 50872 5356 50924
rect 5408 50872 5414 50924
rect 2501 50847 2559 50853
rect 2501 50813 2513 50847
rect 2547 50813 2559 50847
rect 2501 50807 2559 50813
rect 1688 50748 2176 50776
rect 2516 50776 2544 50807
rect 2590 50804 2596 50856
rect 2648 50804 2654 50856
rect 2774 50804 2780 50856
rect 2832 50844 2838 50856
rect 3329 50847 3387 50853
rect 3329 50844 3341 50847
rect 2832 50816 3341 50844
rect 2832 50804 2838 50816
rect 3329 50813 3341 50816
rect 3375 50844 3387 50847
rect 4062 50844 4068 50856
rect 3375 50816 4068 50844
rect 3375 50813 3387 50816
rect 3329 50807 3387 50813
rect 4062 50804 4068 50816
rect 4120 50804 4126 50856
rect 4982 50804 4988 50856
rect 5040 50804 5046 50856
rect 5166 50804 5172 50856
rect 5224 50844 5230 50856
rect 5368 50844 5396 50872
rect 5224 50816 5396 50844
rect 5224 50804 5230 50816
rect 5442 50804 5448 50856
rect 5500 50844 5506 50856
rect 6638 50844 6644 50856
rect 5500 50816 6644 50844
rect 5500 50804 5506 50816
rect 6638 50804 6644 50816
rect 6696 50804 6702 50856
rect 6178 50776 6184 50788
rect 2516 50748 6184 50776
rect 1394 50668 1400 50720
rect 1452 50708 1458 50720
rect 1688 50708 1716 50748
rect 6178 50736 6184 50748
rect 6236 50736 6242 50788
rect 1452 50680 1716 50708
rect 1949 50711 2007 50717
rect 1452 50668 1458 50680
rect 1949 50677 1961 50711
rect 1995 50708 2007 50711
rect 2958 50708 2964 50720
rect 1995 50680 2964 50708
rect 1995 50677 2007 50680
rect 1949 50671 2007 50677
rect 2958 50668 2964 50680
rect 3016 50668 3022 50720
rect 3697 50711 3755 50717
rect 3697 50677 3709 50711
rect 3743 50708 3755 50711
rect 9646 50708 9674 50952
rect 10152 50921 10180 50952
rect 10137 50915 10195 50921
rect 10137 50881 10149 50915
rect 10183 50881 10195 50915
rect 10137 50875 10195 50881
rect 3743 50680 9674 50708
rect 3743 50677 3755 50680
rect 3697 50671 3755 50677
rect 1104 50618 10856 50640
rect 1104 50566 2582 50618
rect 2634 50566 2646 50618
rect 2698 50566 2710 50618
rect 2762 50566 2774 50618
rect 2826 50566 2838 50618
rect 2890 50566 5846 50618
rect 5898 50566 5910 50618
rect 5962 50566 5974 50618
rect 6026 50566 6038 50618
rect 6090 50566 6102 50618
rect 6154 50566 9110 50618
rect 9162 50566 9174 50618
rect 9226 50566 9238 50618
rect 9290 50566 9302 50618
rect 9354 50566 9366 50618
rect 9418 50566 10856 50618
rect 1104 50544 10856 50566
rect 1578 50504 1584 50516
rect 440 50476 980 50504
rect 1044 50476 1584 50504
rect 440 50464 446 50476
rect 952 50436 980 50476
rect 1578 50464 1584 50476
rect 1636 50464 1642 50516
rect 1026 50436 1032 50448
rect 952 50408 1032 50436
rect 1026 50396 1032 50408
rect 1084 50396 1090 50448
rect 2866 50396 2872 50448
rect 2924 50436 2930 50448
rect 4154 50436 4160 50448
rect 2924 50408 4160 50436
rect 2924 50396 2930 50408
rect 4154 50396 4160 50408
rect 4212 50396 4218 50448
rect 106 50328 112 50380
rect 164 50368 170 50380
rect 382 50368 388 50380
rect 164 50340 388 50368
rect 164 50328 170 50340
rect 382 50328 388 50340
rect 440 50328 446 50380
rect 8478 50368 8484 50380
rect 1412 50340 8484 50368
rect 1412 50309 1440 50340
rect 8478 50328 8484 50340
rect 8536 50328 8542 50380
rect 1397 50303 1455 50309
rect 1397 50269 1409 50303
rect 1443 50269 1455 50303
rect 1578 50300 1584 50312
rect 1539 50272 1584 50300
rect 1397 50263 1455 50269
rect 1578 50260 1584 50272
rect 1636 50260 1642 50312
rect 1762 50300 1768 50312
rect 1723 50272 1768 50300
rect 1762 50260 1768 50272
rect 1820 50260 1826 50312
rect 2409 50303 2467 50309
rect 2409 50269 2421 50303
rect 2455 50300 2467 50303
rect 7098 50300 7104 50312
rect 2455 50272 7104 50300
rect 2455 50269 2467 50272
rect 2409 50263 2467 50269
rect 7098 50260 7104 50272
rect 7156 50260 7162 50312
rect 9858 50300 9864 50312
rect 9819 50272 9864 50300
rect 9858 50260 9864 50272
rect 9916 50260 9922 50312
rect 934 50192 940 50244
rect 992 50232 998 50244
rect 1673 50235 1731 50241
rect 1673 50232 1685 50235
rect 992 50204 1685 50232
rect 992 50192 998 50204
rect 1673 50201 1685 50204
rect 1719 50201 1731 50235
rect 1673 50195 1731 50201
rect 1486 50124 1492 50176
rect 1544 50164 1550 50176
rect 1949 50167 2007 50173
rect 1949 50164 1961 50167
rect 1544 50136 1961 50164
rect 1544 50124 1550 50136
rect 1949 50133 1961 50136
rect 1995 50133 2007 50167
rect 1949 50127 2007 50133
rect 2593 50167 2651 50173
rect 2593 50133 2605 50167
rect 2639 50164 2651 50167
rect 2774 50164 2780 50176
rect 2639 50136 2780 50164
rect 2639 50133 2651 50136
rect 2593 50127 2651 50133
rect 2774 50124 2780 50136
rect 2832 50124 2838 50176
rect 10042 50164 10048 50176
rect 10003 50136 10048 50164
rect 10042 50124 10048 50136
rect 10100 50124 10106 50176
rect 1104 50074 10856 50096
rect 1104 50022 4214 50074
rect 4266 50022 4278 50074
rect 4330 50022 4342 50074
rect 4394 50022 4406 50074
rect 4458 50022 4470 50074
rect 4522 50022 7478 50074
rect 7530 50022 7542 50074
rect 7594 50022 7606 50074
rect 7658 50022 7670 50074
rect 7722 50022 7734 50074
rect 7786 50022 10856 50074
rect 1104 50000 10856 50022
rect 9582 49920 9588 49972
rect 9640 49960 9646 49972
rect 10045 49963 10103 49969
rect 10045 49960 10057 49963
rect 9640 49932 10057 49960
rect 9640 49920 9646 49932
rect 10045 49929 10057 49932
rect 10091 49929 10103 49963
rect 10045 49923 10103 49929
rect 1670 49892 1676 49904
rect 1631 49864 1676 49892
rect 1670 49852 1676 49864
rect 1728 49852 1734 49904
rect 1118 49784 1124 49836
rect 1176 49824 1182 49836
rect 1397 49827 1455 49833
rect 1397 49824 1409 49827
rect 1176 49796 1409 49824
rect 1176 49784 1182 49796
rect 1397 49793 1409 49796
rect 1443 49793 1455 49827
rect 1578 49824 1584 49836
rect 1539 49796 1584 49824
rect 1397 49787 1455 49793
rect 1578 49784 1584 49796
rect 1636 49784 1642 49836
rect 1762 49824 1768 49836
rect 1723 49796 1768 49824
rect 1762 49784 1768 49796
rect 1820 49784 1826 49836
rect 2409 49827 2467 49833
rect 2409 49793 2421 49827
rect 2455 49824 2467 49827
rect 2498 49824 2504 49836
rect 2455 49796 2504 49824
rect 2455 49793 2467 49796
rect 2409 49787 2467 49793
rect 2498 49784 2504 49796
rect 2556 49784 2562 49836
rect 9861 49827 9919 49833
rect 9861 49793 9873 49827
rect 9907 49824 9919 49827
rect 9950 49824 9956 49836
rect 9907 49796 9956 49824
rect 9907 49793 9919 49796
rect 9861 49787 9919 49793
rect 9950 49784 9956 49796
rect 10008 49784 10014 49836
rect 2590 49756 2596 49768
rect 1872 49728 2596 49756
rect 1762 49648 1768 49700
rect 1820 49688 1826 49700
rect 1872 49688 1900 49728
rect 2590 49716 2596 49728
rect 2648 49716 2654 49768
rect 3786 49716 3792 49768
rect 3844 49756 3850 49768
rect 3970 49756 3976 49768
rect 3844 49728 3976 49756
rect 3844 49716 3850 49728
rect 3970 49716 3976 49728
rect 4028 49716 4034 49768
rect 1820 49660 1900 49688
rect 1949 49691 2007 49697
rect 1820 49648 1826 49660
rect 1949 49657 1961 49691
rect 1995 49657 2007 49691
rect 1949 49651 2007 49657
rect 1118 49580 1124 49632
rect 1176 49620 1182 49632
rect 1964 49620 1992 49651
rect 1176 49592 1992 49620
rect 1176 49580 1182 49592
rect 2498 49580 2504 49632
rect 2556 49620 2562 49632
rect 2593 49623 2651 49629
rect 2593 49620 2605 49623
rect 2556 49592 2605 49620
rect 2556 49580 2562 49592
rect 2593 49589 2605 49592
rect 2639 49589 2651 49623
rect 2593 49583 2651 49589
rect 3418 49580 3424 49632
rect 3476 49620 3482 49632
rect 3970 49620 3976 49632
rect 3476 49592 3976 49620
rect 3476 49580 3482 49592
rect 3970 49580 3976 49592
rect 4028 49580 4034 49632
rect 1104 49530 10856 49552
rect 1104 49478 2582 49530
rect 2634 49478 2646 49530
rect 2698 49478 2710 49530
rect 2762 49478 2774 49530
rect 2826 49478 2838 49530
rect 2890 49478 5846 49530
rect 5898 49478 5910 49530
rect 5962 49478 5974 49530
rect 6026 49478 6038 49530
rect 6090 49478 6102 49530
rect 6154 49478 9110 49530
rect 9162 49478 9174 49530
rect 9226 49478 9238 49530
rect 9290 49478 9302 49530
rect 9354 49478 9366 49530
rect 9418 49478 10856 49530
rect 1104 49456 10856 49478
rect 14 49376 20 49428
rect 72 49416 78 49428
rect 2406 49416 2412 49428
rect 72 49388 2412 49416
rect 72 49376 78 49388
rect 2406 49376 2412 49388
rect 2464 49376 2470 49428
rect 3510 49376 3516 49428
rect 3568 49416 3574 49428
rect 3878 49416 3884 49428
rect 3568 49388 3884 49416
rect 3568 49376 3574 49388
rect 3878 49376 3884 49388
rect 3936 49376 3942 49428
rect 9217 49419 9275 49425
rect 9217 49385 9229 49419
rect 9263 49416 9275 49419
rect 9674 49416 9680 49428
rect 9263 49388 9680 49416
rect 9263 49385 9275 49388
rect 9217 49379 9275 49385
rect 9674 49376 9680 49388
rect 9732 49376 9738 49428
rect 1394 49308 1400 49360
rect 1452 49348 1458 49360
rect 1670 49348 1676 49360
rect 1452 49320 1676 49348
rect 1452 49308 1458 49320
rect 1670 49308 1676 49320
rect 1728 49308 1734 49360
rect 2682 49308 2688 49360
rect 2740 49348 2746 49360
rect 4522 49348 4528 49360
rect 2740 49320 4528 49348
rect 2740 49308 2746 49320
rect 4522 49308 4528 49320
rect 4580 49308 4586 49360
rect 2866 49280 2872 49292
rect 1412 49252 2872 49280
rect 1412 49221 1440 49252
rect 2866 49240 2872 49252
rect 2924 49240 2930 49292
rect 1397 49215 1455 49221
rect 1397 49181 1409 49215
rect 1443 49181 1455 49215
rect 1397 49175 1455 49181
rect 2133 49215 2191 49221
rect 2133 49181 2145 49215
rect 2179 49212 2191 49215
rect 2179 49184 2774 49212
rect 2179 49181 2191 49184
rect 2133 49175 2191 49181
rect 2746 49144 2774 49184
rect 6546 49172 6552 49224
rect 6604 49212 6610 49224
rect 9401 49215 9459 49221
rect 9401 49212 9413 49215
rect 6604 49184 9413 49212
rect 6604 49172 6610 49184
rect 9401 49181 9413 49184
rect 9447 49181 9459 49215
rect 9401 49175 9459 49181
rect 9490 49172 9496 49224
rect 9548 49212 9554 49224
rect 9861 49215 9919 49221
rect 9861 49212 9873 49215
rect 9548 49184 9873 49212
rect 9548 49172 9554 49184
rect 9861 49181 9873 49184
rect 9907 49181 9919 49215
rect 9861 49175 9919 49181
rect 6730 49144 6736 49156
rect 2746 49116 6736 49144
rect 6730 49104 6736 49116
rect 6788 49104 6794 49156
rect 1394 49036 1400 49088
rect 1452 49076 1458 49088
rect 1581 49079 1639 49085
rect 1581 49076 1593 49079
rect 1452 49048 1593 49076
rect 1452 49036 1458 49048
rect 1581 49045 1593 49048
rect 1627 49045 1639 49079
rect 2314 49076 2320 49088
rect 2275 49048 2320 49076
rect 1581 49039 1639 49045
rect 2314 49036 2320 49048
rect 2372 49036 2378 49088
rect 10042 49076 10048 49088
rect 10003 49048 10048 49076
rect 10042 49036 10048 49048
rect 10100 49036 10106 49088
rect 1104 48986 10856 49008
rect 1104 48934 4214 48986
rect 4266 48934 4278 48986
rect 4330 48934 4342 48986
rect 4394 48934 4406 48986
rect 4458 48934 4470 48986
rect 4522 48934 7478 48986
rect 7530 48934 7542 48986
rect 7594 48934 7606 48986
rect 7658 48934 7670 48986
rect 7722 48934 7734 48986
rect 7786 48934 10856 48986
rect 1104 48912 10856 48934
rect 9858 48832 9864 48884
rect 9916 48872 9922 48884
rect 9953 48875 10011 48881
rect 9953 48872 9965 48875
rect 9916 48844 9965 48872
rect 9916 48832 9922 48844
rect 9953 48841 9965 48844
rect 9999 48841 10011 48875
rect 9953 48835 10011 48841
rect 2682 48804 2688 48816
rect 1412 48776 2688 48804
rect 1412 48745 1440 48776
rect 2682 48764 2688 48776
rect 2740 48764 2746 48816
rect 2958 48764 2964 48816
rect 3016 48804 3022 48816
rect 3016 48776 3188 48804
rect 3016 48764 3022 48776
rect 3160 48748 3188 48776
rect 3344 48776 3832 48804
rect 1397 48739 1455 48745
rect 1397 48705 1409 48739
rect 1443 48705 1455 48739
rect 1397 48699 1455 48705
rect 2593 48739 2651 48745
rect 2593 48705 2605 48739
rect 2639 48736 2651 48739
rect 2774 48736 2780 48748
rect 2639 48708 2780 48736
rect 2639 48705 2651 48708
rect 2593 48699 2651 48705
rect 2774 48696 2780 48708
rect 2832 48696 2838 48748
rect 3142 48696 3148 48748
rect 3200 48736 3206 48748
rect 3344 48736 3372 48776
rect 3804 48745 3832 48776
rect 3605 48739 3663 48745
rect 3605 48736 3617 48739
rect 3200 48708 3372 48736
rect 3436 48708 3617 48736
rect 3200 48696 3206 48708
rect 2317 48671 2375 48677
rect 2317 48637 2329 48671
rect 2363 48668 2375 48671
rect 2958 48668 2964 48680
rect 2363 48640 2964 48668
rect 2363 48637 2375 48640
rect 2317 48631 2375 48637
rect 2958 48628 2964 48640
rect 3016 48628 3022 48680
rect 1118 48532 1124 48544
rect 1044 48504 1124 48532
rect 1044 48056 1072 48504
rect 1118 48492 1124 48504
rect 1176 48492 1182 48544
rect 1578 48532 1584 48544
rect 1539 48504 1584 48532
rect 1578 48492 1584 48504
rect 1636 48492 1642 48544
rect 3436 48532 3464 48708
rect 3605 48705 3617 48708
rect 3651 48705 3663 48739
rect 3605 48699 3663 48705
rect 3789 48739 3847 48745
rect 3789 48705 3801 48739
rect 3835 48705 3847 48739
rect 10134 48736 10140 48748
rect 10095 48708 10140 48736
rect 3789 48699 3847 48705
rect 10134 48696 10140 48708
rect 10192 48696 10198 48748
rect 3973 48603 4031 48609
rect 3973 48569 3985 48603
rect 4019 48569 4031 48603
rect 3973 48563 4031 48569
rect 3510 48532 3516 48544
rect 3436 48504 3516 48532
rect 3510 48492 3516 48504
rect 3568 48492 3574 48544
rect 3988 48532 4016 48563
rect 6546 48532 6552 48544
rect 3988 48504 6552 48532
rect 6546 48492 6552 48504
rect 6604 48492 6610 48544
rect 1104 48442 10856 48464
rect 1104 48390 2582 48442
rect 2634 48390 2646 48442
rect 2698 48390 2710 48442
rect 2762 48390 2774 48442
rect 2826 48390 2838 48442
rect 2890 48390 5846 48442
rect 5898 48390 5910 48442
rect 5962 48390 5974 48442
rect 6026 48390 6038 48442
rect 6090 48390 6102 48442
rect 6154 48390 9110 48442
rect 9162 48390 9174 48442
rect 9226 48390 9238 48442
rect 9290 48390 9302 48442
rect 9354 48390 9366 48442
rect 9418 48390 10856 48442
rect 1104 48368 10856 48390
rect 1762 48288 1768 48340
rect 1820 48288 1826 48340
rect 4522 48328 4528 48340
rect 2700 48326 4528 48328
rect 1780 48260 1808 48288
rect 2682 48274 2688 48326
rect 2740 48300 4528 48326
rect 2740 48274 2746 48300
rect 4522 48288 4528 48300
rect 4580 48288 4586 48340
rect 1780 48232 2636 48260
rect 2608 48136 2636 48232
rect 2774 48220 2780 48272
rect 2832 48260 2838 48272
rect 6178 48260 6184 48272
rect 2832 48232 2877 48260
rect 4540 48232 6184 48260
rect 2832 48220 2838 48232
rect 4540 48192 4568 48232
rect 6178 48220 6184 48232
rect 6236 48260 6242 48272
rect 7190 48260 7196 48272
rect 6236 48232 7196 48260
rect 6236 48220 6242 48232
rect 7190 48220 7196 48232
rect 7248 48220 7254 48272
rect 9217 48263 9275 48269
rect 9217 48229 9229 48263
rect 9263 48260 9275 48263
rect 9490 48260 9496 48272
rect 9263 48232 9496 48260
rect 9263 48229 9275 48232
rect 9217 48223 9275 48229
rect 9490 48220 9496 48232
rect 9548 48220 9554 48272
rect 4356 48164 4568 48192
rect 4617 48195 4675 48201
rect 1394 48124 1400 48136
rect 1355 48096 1400 48124
rect 1394 48084 1400 48096
rect 1452 48084 1458 48136
rect 2406 48124 2412 48136
rect 2367 48096 2412 48124
rect 2406 48084 2412 48096
rect 2464 48084 2470 48136
rect 2590 48124 2596 48136
rect 2551 48096 2596 48124
rect 2590 48084 2596 48096
rect 2648 48084 2654 48136
rect 4356 48133 4384 48164
rect 4617 48161 4629 48195
rect 4663 48192 4675 48195
rect 4663 48164 9444 48192
rect 4663 48161 4675 48164
rect 4617 48155 4675 48161
rect 9416 48133 9444 48164
rect 4341 48127 4399 48133
rect 4341 48093 4353 48127
rect 4387 48093 4399 48127
rect 4341 48087 4399 48093
rect 4433 48127 4491 48133
rect 4433 48093 4445 48127
rect 4479 48093 4491 48127
rect 4433 48087 4491 48093
rect 5077 48127 5135 48133
rect 5077 48093 5089 48127
rect 5123 48093 5135 48127
rect 5077 48087 5135 48093
rect 5261 48127 5319 48133
rect 5261 48093 5273 48127
rect 5307 48093 5319 48127
rect 5261 48087 5319 48093
rect 5445 48127 5503 48133
rect 5445 48093 5457 48127
rect 5491 48124 5503 48127
rect 7009 48127 7067 48133
rect 7009 48124 7021 48127
rect 5491 48096 7021 48124
rect 5491 48093 5503 48096
rect 5445 48087 5503 48093
rect 7009 48093 7021 48096
rect 7055 48093 7067 48127
rect 7009 48087 7067 48093
rect 9401 48127 9459 48133
rect 9401 48093 9413 48127
rect 9447 48093 9459 48127
rect 9401 48087 9459 48093
rect 9861 48127 9919 48133
rect 9861 48093 9873 48127
rect 9907 48093 9919 48127
rect 9861 48087 9919 48093
rect 2958 48056 2964 48068
rect 1044 48028 2964 48056
rect 2958 48016 2964 48028
rect 3016 48016 3022 48068
rect 1578 47988 1584 48000
rect 1539 47960 1584 47988
rect 1578 47948 1584 47960
rect 1636 47948 1642 48000
rect 4448 47988 4476 48087
rect 4522 48016 4528 48068
rect 4580 48056 4586 48068
rect 5092 48056 5120 48087
rect 4580 48028 5120 48056
rect 5276 48056 5304 48087
rect 6178 48056 6184 48068
rect 5276 48028 6184 48056
rect 4580 48016 4586 48028
rect 5276 47988 5304 48028
rect 6178 48016 6184 48028
rect 6236 48016 6242 48068
rect 9876 48056 9904 48087
rect 6840 48028 9904 48056
rect 6840 47997 6868 48028
rect 4448 47960 5304 47988
rect 6825 47991 6883 47997
rect 6825 47957 6837 47991
rect 6871 47957 6883 47991
rect 10042 47988 10048 48000
rect 10003 47960 10048 47988
rect 6825 47951 6883 47957
rect 10042 47948 10048 47960
rect 10100 47948 10106 48000
rect 1104 47898 10856 47920
rect 1104 47846 4214 47898
rect 4266 47846 4278 47898
rect 4330 47846 4342 47898
rect 4394 47846 4406 47898
rect 4458 47846 4470 47898
rect 4522 47846 7478 47898
rect 7530 47846 7542 47898
rect 7594 47846 7606 47898
rect 7658 47846 7670 47898
rect 7722 47846 7734 47898
rect 7786 47846 10856 47898
rect 1104 47824 10856 47846
rect 3510 47784 3516 47796
rect 1504 47756 3516 47784
rect 1504 47657 1532 47756
rect 3510 47744 3516 47756
rect 3568 47744 3574 47796
rect 2590 47716 2596 47728
rect 1596 47688 2596 47716
rect 1596 47657 1624 47688
rect 2590 47676 2596 47688
rect 2648 47676 2654 47728
rect 3878 47716 3884 47728
rect 3436 47688 3884 47716
rect 1489 47651 1547 47657
rect 1489 47617 1501 47651
rect 1535 47617 1547 47651
rect 1489 47611 1547 47617
rect 1581 47651 1639 47657
rect 1581 47617 1593 47651
rect 1627 47617 1639 47651
rect 1581 47611 1639 47617
rect 2501 47651 2559 47657
rect 2501 47617 2513 47651
rect 2547 47648 2559 47651
rect 3436 47648 3464 47688
rect 3878 47676 3884 47688
rect 3936 47676 3942 47728
rect 2547 47620 3464 47648
rect 3513 47651 3571 47657
rect 2547 47617 2559 47620
rect 2501 47611 2559 47617
rect 3513 47617 3525 47651
rect 3559 47617 3571 47651
rect 3513 47611 3571 47617
rect 1596 47580 1624 47611
rect 1044 47552 1624 47580
rect 2225 47583 2283 47589
rect 1044 47172 1072 47552
rect 2225 47549 2237 47583
rect 2271 47580 2283 47583
rect 2406 47580 2412 47592
rect 2271 47552 2412 47580
rect 2271 47549 2283 47552
rect 2225 47543 2283 47549
rect 2406 47540 2412 47552
rect 2464 47540 2470 47592
rect 3142 47540 3148 47592
rect 3200 47580 3206 47592
rect 3418 47580 3424 47592
rect 3200 47552 3424 47580
rect 3200 47540 3206 47552
rect 3418 47540 3424 47552
rect 3476 47540 3482 47592
rect 3528 47580 3556 47611
rect 7466 47608 7472 47660
rect 7524 47648 7530 47660
rect 9861 47651 9919 47657
rect 9861 47648 9873 47651
rect 7524 47620 9873 47648
rect 7524 47608 7530 47620
rect 9861 47617 9873 47620
rect 9907 47617 9919 47651
rect 9861 47611 9919 47617
rect 3878 47580 3884 47592
rect 3528 47552 3884 47580
rect 3878 47540 3884 47552
rect 3936 47540 3942 47592
rect 1486 47404 1492 47456
rect 1544 47444 1550 47456
rect 1765 47447 1823 47453
rect 1765 47444 1777 47447
rect 1544 47416 1777 47444
rect 1544 47404 1550 47416
rect 1765 47413 1777 47416
rect 1811 47413 1823 47447
rect 3694 47444 3700 47456
rect 3655 47416 3700 47444
rect 1765 47407 1823 47413
rect 3694 47404 3700 47416
rect 3752 47404 3758 47456
rect 10042 47444 10048 47456
rect 10003 47416 10048 47444
rect 10042 47404 10048 47416
rect 10100 47404 10106 47456
rect 1104 47354 10856 47376
rect 1104 47302 2582 47354
rect 2634 47302 2646 47354
rect 2698 47302 2710 47354
rect 2762 47302 2774 47354
rect 2826 47302 2838 47354
rect 2890 47302 5846 47354
rect 5898 47302 5910 47354
rect 5962 47302 5974 47354
rect 6026 47302 6038 47354
rect 6090 47302 6102 47354
rect 6154 47302 9110 47354
rect 9162 47302 9174 47354
rect 9226 47302 9238 47354
rect 9290 47302 9302 47354
rect 9354 47302 9366 47354
rect 9418 47302 10856 47354
rect 1104 47280 10856 47302
rect 2406 47200 2412 47252
rect 2464 47240 2470 47252
rect 3145 47243 3203 47249
rect 3145 47240 3157 47243
rect 2464 47212 3157 47240
rect 2464 47200 2470 47212
rect 3145 47209 3157 47212
rect 3191 47209 3203 47243
rect 7282 47240 7288 47252
rect 3145 47203 3203 47209
rect 3804 47212 7288 47240
rect 1044 47144 2452 47172
rect 2424 47116 2452 47144
rect 1486 47104 1492 47116
rect 1447 47076 1492 47104
rect 1486 47064 1492 47076
rect 1544 47064 1550 47116
rect 1762 47104 1768 47116
rect 1723 47076 1768 47104
rect 1762 47064 1768 47076
rect 1820 47064 1826 47116
rect 2406 47064 2412 47116
rect 2464 47104 2470 47116
rect 2464 47076 3004 47104
rect 2464 47064 2470 47076
rect 2976 47045 3004 47076
rect 3804 47045 3832 47212
rect 7282 47200 7288 47212
rect 7340 47200 7346 47252
rect 7466 47240 7472 47252
rect 7427 47212 7472 47240
rect 7466 47200 7472 47212
rect 7524 47200 7530 47252
rect 9950 47240 9956 47252
rect 9911 47212 9956 47240
rect 9950 47200 9956 47212
rect 10008 47200 10014 47252
rect 4614 47132 4620 47184
rect 4672 47172 4678 47184
rect 5166 47172 5172 47184
rect 4672 47144 5172 47172
rect 4672 47132 4678 47144
rect 5166 47132 5172 47144
rect 5224 47132 5230 47184
rect 5810 47104 5816 47116
rect 5184 47076 5816 47104
rect 2869 47039 2927 47045
rect 2869 47005 2881 47039
rect 2915 47005 2927 47039
rect 2869 46999 2927 47005
rect 2961 47039 3019 47045
rect 2961 47005 2973 47039
rect 3007 47005 3019 47039
rect 2961 46999 3019 47005
rect 3789 47039 3847 47045
rect 3789 47005 3801 47039
rect 3835 47005 3847 47039
rect 3789 46999 3847 47005
rect 1486 46928 1492 46980
rect 1544 46968 1550 46980
rect 1670 46968 1676 46980
rect 1544 46940 1676 46968
rect 1544 46928 1550 46940
rect 1670 46928 1676 46940
rect 1728 46928 1734 46980
rect 2884 46968 2912 46999
rect 4522 46996 4528 47048
rect 4580 47036 4586 47048
rect 5184 47045 5212 47076
rect 5810 47064 5816 47076
rect 5868 47104 5874 47116
rect 6178 47104 6184 47116
rect 5868 47076 6184 47104
rect 5868 47064 5874 47076
rect 6178 47064 6184 47076
rect 6236 47064 6242 47116
rect 4985 47039 5043 47045
rect 4985 47036 4997 47039
rect 4580 47008 4997 47036
rect 4580 46996 4586 47008
rect 4985 47005 4997 47008
rect 5031 47005 5043 47039
rect 4985 46999 5043 47005
rect 5169 47039 5227 47045
rect 5169 47005 5181 47039
rect 5215 47005 5227 47039
rect 5169 46999 5227 47005
rect 5353 47039 5411 47045
rect 5353 47005 5365 47039
rect 5399 47036 5411 47039
rect 7653 47039 7711 47045
rect 7653 47036 7665 47039
rect 5399 47008 7665 47036
rect 5399 47005 5411 47008
rect 5353 46999 5411 47005
rect 7653 47005 7665 47008
rect 7699 47005 7711 47039
rect 7653 46999 7711 47005
rect 10137 47039 10195 47045
rect 10137 47005 10149 47039
rect 10183 47005 10195 47039
rect 10137 46999 10195 47005
rect 4540 46968 4568 46996
rect 10152 46968 10180 46999
rect 2884 46940 4568 46968
rect 5184 46940 10180 46968
rect 5184 46912 5212 46940
rect 3970 46900 3976 46912
rect 3931 46872 3976 46900
rect 3970 46860 3976 46872
rect 4028 46860 4034 46912
rect 5166 46860 5172 46912
rect 5224 46860 5230 46912
rect 1104 46810 10856 46832
rect 1104 46758 4214 46810
rect 4266 46758 4278 46810
rect 4330 46758 4342 46810
rect 4394 46758 4406 46810
rect 4458 46758 4470 46810
rect 4522 46758 7478 46810
rect 7530 46758 7542 46810
rect 7594 46758 7606 46810
rect 7658 46758 7670 46810
rect 7722 46758 7734 46810
rect 7786 46758 10856 46810
rect 1104 46736 10856 46758
rect 106 46656 112 46708
rect 164 46696 170 46708
rect 1394 46696 1400 46708
rect 164 46668 1400 46696
rect 164 46656 170 46668
rect 1394 46656 1400 46668
rect 1452 46656 1458 46708
rect 1762 46656 1768 46708
rect 1820 46696 1826 46708
rect 1946 46696 1952 46708
rect 1820 46668 1952 46696
rect 1820 46656 1826 46668
rect 1946 46656 1952 46668
rect 2004 46656 2010 46708
rect 3237 46699 3295 46705
rect 3237 46665 3249 46699
rect 3283 46696 3295 46699
rect 10134 46696 10140 46708
rect 3283 46668 10140 46696
rect 3283 46665 3295 46668
rect 3237 46659 3295 46665
rect 10134 46656 10140 46668
rect 10192 46656 10198 46708
rect 106 46520 112 46572
rect 164 46560 170 46572
rect 1581 46563 1639 46569
rect 1581 46560 1593 46563
rect 164 46532 1593 46560
rect 164 46520 170 46532
rect 1581 46529 1593 46532
rect 1627 46529 1639 46563
rect 1581 46523 1639 46529
rect 1765 46563 1823 46569
rect 1765 46529 1777 46563
rect 1811 46560 1823 46563
rect 2406 46560 2412 46572
rect 1811 46532 2412 46560
rect 1811 46529 1823 46532
rect 1765 46523 1823 46529
rect 1596 46492 1624 46523
rect 2406 46520 2412 46532
rect 2464 46520 2470 46572
rect 3053 46563 3111 46569
rect 3053 46529 3065 46563
rect 3099 46529 3111 46563
rect 3694 46560 3700 46572
rect 3655 46532 3700 46560
rect 3053 46523 3111 46529
rect 2869 46495 2927 46501
rect 2869 46492 2881 46495
rect 1596 46464 2881 46492
rect 2869 46461 2881 46464
rect 2915 46461 2927 46495
rect 3068 46492 3096 46523
rect 3694 46520 3700 46532
rect 3752 46520 3758 46572
rect 5718 46520 5724 46572
rect 5776 46560 5782 46572
rect 6546 46560 6552 46572
rect 5776 46532 6552 46560
rect 5776 46520 5782 46532
rect 6546 46520 6552 46532
rect 6604 46520 6610 46572
rect 7006 46520 7012 46572
rect 7064 46560 7070 46572
rect 9861 46563 9919 46569
rect 9861 46560 9873 46563
rect 7064 46532 9873 46560
rect 7064 46520 7070 46532
rect 9861 46529 9873 46532
rect 9907 46529 9919 46563
rect 9861 46523 9919 46529
rect 3326 46492 3332 46504
rect 3068 46464 3332 46492
rect 2869 46455 2927 46461
rect 3326 46452 3332 46464
rect 3384 46492 3390 46504
rect 4154 46492 4160 46504
rect 3384 46464 4160 46492
rect 3384 46452 3390 46464
rect 4154 46452 4160 46464
rect 4212 46452 4218 46504
rect 5626 46452 5632 46504
rect 5684 46492 5690 46504
rect 6178 46492 6184 46504
rect 5684 46464 6184 46492
rect 5684 46452 5690 46464
rect 6178 46452 6184 46464
rect 6236 46452 6242 46504
rect 3878 46424 3884 46436
rect 3839 46396 3884 46424
rect 3878 46384 3884 46396
rect 3936 46384 3942 46436
rect 10042 46424 10048 46436
rect 10003 46396 10048 46424
rect 10042 46384 10048 46396
rect 10100 46384 10106 46436
rect 1394 46316 1400 46368
rect 1452 46356 1458 46368
rect 1949 46359 2007 46365
rect 1949 46356 1961 46359
rect 1452 46328 1961 46356
rect 1452 46316 1458 46328
rect 1949 46325 1961 46328
rect 1995 46325 2007 46359
rect 1949 46319 2007 46325
rect 4982 46316 4988 46368
rect 5040 46356 5046 46368
rect 6638 46356 6644 46368
rect 5040 46328 6644 46356
rect 5040 46316 5046 46328
rect 6638 46316 6644 46328
rect 6696 46316 6702 46368
rect 1104 46266 10856 46288
rect 1104 46214 2582 46266
rect 2634 46214 2646 46266
rect 2698 46214 2710 46266
rect 2762 46214 2774 46266
rect 2826 46214 2838 46266
rect 2890 46214 5846 46266
rect 5898 46214 5910 46266
rect 5962 46214 5974 46266
rect 6026 46214 6038 46266
rect 6090 46214 6102 46266
rect 6154 46214 9110 46266
rect 9162 46214 9174 46266
rect 9226 46214 9238 46266
rect 9290 46214 9302 46266
rect 9354 46214 9366 46266
rect 9418 46214 10856 46266
rect 1104 46192 10856 46214
rect 3050 46044 3056 46096
rect 3108 46084 3114 46096
rect 3234 46084 3240 46096
rect 3108 46056 3240 46084
rect 3108 46044 3114 46056
rect 3234 46044 3240 46056
rect 3292 46044 3298 46096
rect 4522 46044 4528 46096
rect 4580 46084 4586 46096
rect 4706 46084 4712 46096
rect 4580 46056 4712 46084
rect 4580 46044 4586 46056
rect 4706 46044 4712 46056
rect 4764 46044 4770 46096
rect 1394 46016 1400 46028
rect 1355 45988 1400 46016
rect 1394 45976 1400 45988
rect 1452 45976 1458 46028
rect 1670 46016 1676 46028
rect 1631 45988 1676 46016
rect 1670 45976 1676 45988
rect 1728 45976 1734 46028
rect 2682 45948 2688 45960
rect 2643 45920 2688 45948
rect 2682 45908 2688 45920
rect 2740 45908 2746 45960
rect 3786 45948 3792 45960
rect 3747 45920 3792 45948
rect 3786 45908 3792 45920
rect 3844 45908 3850 45960
rect 9858 45948 9864 45960
rect 9819 45920 9864 45948
rect 9858 45908 9864 45920
rect 9916 45908 9922 45960
rect 3050 45840 3056 45892
rect 3108 45880 3114 45892
rect 4154 45880 4160 45892
rect 3108 45852 4160 45880
rect 3108 45840 3114 45852
rect 4154 45840 4160 45852
rect 4212 45840 4218 45892
rect 2866 45812 2872 45824
rect 2827 45784 2872 45812
rect 2866 45772 2872 45784
rect 2924 45772 2930 45824
rect 3970 45812 3976 45824
rect 3931 45784 3976 45812
rect 3970 45772 3976 45784
rect 4028 45772 4034 45824
rect 5534 45772 5540 45824
rect 5592 45812 5598 45824
rect 5718 45812 5724 45824
rect 5592 45784 5724 45812
rect 5592 45772 5598 45784
rect 5718 45772 5724 45784
rect 5776 45772 5782 45824
rect 10042 45812 10048 45824
rect 10003 45784 10048 45812
rect 10042 45772 10048 45784
rect 10100 45772 10106 45824
rect 1104 45722 10856 45744
rect 1104 45670 4214 45722
rect 4266 45670 4278 45722
rect 4330 45670 4342 45722
rect 4394 45670 4406 45722
rect 4458 45670 4470 45722
rect 4522 45670 7478 45722
rect 7530 45670 7542 45722
rect 7594 45670 7606 45722
rect 7658 45670 7670 45722
rect 7722 45670 7734 45722
rect 7786 45670 10856 45722
rect 1104 45648 10856 45670
rect 566 45608 572 45620
rect 32 45580 572 45608
rect 32 45280 60 45580
rect 566 45568 572 45580
rect 624 45568 630 45620
rect 1026 45568 1032 45620
rect 1084 45568 1090 45620
rect 1044 45540 1072 45568
rect 1044 45512 2176 45540
rect 290 45432 296 45484
rect 348 45432 354 45484
rect 1026 45432 1032 45484
rect 1084 45472 1090 45484
rect 1486 45472 1492 45484
rect 1084 45444 1492 45472
rect 1084 45432 1090 45444
rect 1486 45432 1492 45444
rect 1544 45432 1550 45484
rect 2148 45481 2176 45512
rect 2866 45500 2872 45552
rect 2924 45540 2930 45552
rect 3786 45540 3792 45552
rect 2924 45512 3792 45540
rect 2924 45500 2930 45512
rect 3786 45500 3792 45512
rect 3844 45500 3850 45552
rect 2133 45475 2191 45481
rect 2133 45441 2145 45475
rect 2179 45441 2191 45475
rect 2133 45435 2191 45441
rect 308 45404 336 45432
rect 566 45404 572 45416
rect 308 45376 572 45404
rect 566 45364 572 45376
rect 624 45364 630 45416
rect 1854 45404 1860 45416
rect 1815 45376 1860 45404
rect 1854 45364 1860 45376
rect 1912 45364 1918 45416
rect 14 45228 20 45280
rect 72 45228 78 45280
rect 106 45228 112 45280
rect 164 45268 170 45280
rect 290 45268 296 45280
rect 164 45240 296 45268
rect 164 45228 170 45240
rect 290 45228 296 45240
rect 348 45228 354 45280
rect 1104 45178 10856 45200
rect 1104 45126 2582 45178
rect 2634 45126 2646 45178
rect 2698 45126 2710 45178
rect 2762 45126 2774 45178
rect 2826 45126 2838 45178
rect 2890 45126 5846 45178
rect 5898 45126 5910 45178
rect 5962 45126 5974 45178
rect 6026 45126 6038 45178
rect 6090 45126 6102 45178
rect 6154 45126 9110 45178
rect 9162 45126 9174 45178
rect 9226 45126 9238 45178
rect 9290 45126 9302 45178
rect 9354 45126 9366 45178
rect 9418 45126 10856 45178
rect 1104 45104 10856 45126
rect 106 45024 112 45076
rect 164 45064 170 45076
rect 1302 45064 1308 45076
rect 164 45036 1308 45064
rect 164 45024 170 45036
rect 1302 45024 1308 45036
rect 1360 45024 1366 45076
rect 1578 45064 1584 45076
rect 1539 45036 1584 45064
rect 1578 45024 1584 45036
rect 1636 45024 1642 45076
rect 1854 45024 1860 45076
rect 1912 45064 1918 45076
rect 2501 45067 2559 45073
rect 2501 45064 2513 45067
rect 1912 45036 2513 45064
rect 1912 45024 1918 45036
rect 2501 45033 2513 45036
rect 2547 45033 2559 45067
rect 2501 45027 2559 45033
rect 5629 45067 5687 45073
rect 5629 45033 5641 45067
rect 5675 45064 5687 45067
rect 7006 45064 7012 45076
rect 5675 45036 7012 45064
rect 5675 45033 5687 45036
rect 5629 45027 5687 45033
rect 7006 45024 7012 45036
rect 7064 45024 7070 45076
rect 1394 44860 1400 44872
rect 1355 44832 1400 44860
rect 1394 44820 1400 44832
rect 1452 44820 1458 44872
rect 2225 44863 2283 44869
rect 2225 44829 2237 44863
rect 2271 44829 2283 44863
rect 2225 44823 2283 44829
rect 2317 44863 2375 44869
rect 2317 44829 2329 44863
rect 2363 44860 2375 44863
rect 2406 44860 2412 44872
rect 2363 44832 2412 44860
rect 2363 44829 2375 44832
rect 2317 44823 2375 44829
rect 2240 44792 2268 44823
rect 2406 44820 2412 44832
rect 2464 44860 2470 44872
rect 2590 44860 2596 44872
rect 2464 44832 2596 44860
rect 2464 44820 2470 44832
rect 2590 44820 2596 44832
rect 2648 44820 2654 44872
rect 4890 44820 4896 44872
rect 4948 44860 4954 44872
rect 5813 44863 5871 44869
rect 5813 44860 5825 44863
rect 4948 44832 5825 44860
rect 4948 44820 4954 44832
rect 5813 44829 5825 44832
rect 5859 44829 5871 44863
rect 5813 44823 5871 44829
rect 8294 44820 8300 44872
rect 8352 44860 8358 44872
rect 9861 44863 9919 44869
rect 9861 44860 9873 44863
rect 8352 44832 9873 44860
rect 8352 44820 8358 44832
rect 9861 44829 9873 44832
rect 9907 44829 9919 44863
rect 9861 44823 9919 44829
rect 3970 44792 3976 44804
rect 2240 44764 3976 44792
rect 3970 44752 3976 44764
rect 4028 44752 4034 44804
rect 1854 44684 1860 44736
rect 1912 44724 1918 44736
rect 3878 44724 3884 44736
rect 1912 44696 3884 44724
rect 1912 44684 1918 44696
rect 3878 44684 3884 44696
rect 3936 44684 3942 44736
rect 10042 44724 10048 44736
rect 10003 44696 10048 44724
rect 10042 44684 10048 44696
rect 10100 44684 10106 44736
rect 1104 44634 10856 44656
rect 1104 44582 4214 44634
rect 4266 44582 4278 44634
rect 4330 44582 4342 44634
rect 4394 44582 4406 44634
rect 4458 44582 4470 44634
rect 4522 44582 7478 44634
rect 7530 44582 7542 44634
rect 7594 44582 7606 44634
rect 7658 44582 7670 44634
rect 7722 44582 7734 44634
rect 7786 44582 10856 44634
rect 1104 44560 10856 44582
rect 1578 44520 1584 44532
rect 1539 44492 1584 44520
rect 1578 44480 1584 44492
rect 1636 44480 1642 44532
rect 3050 44520 3056 44532
rect 2976 44492 3056 44520
rect 2976 44393 3004 44492
rect 3050 44480 3056 44492
rect 3108 44480 3114 44532
rect 4890 44520 4896 44532
rect 4851 44492 4896 44520
rect 4890 44480 4896 44492
rect 4948 44480 4954 44532
rect 1397 44387 1455 44393
rect 1397 44353 1409 44387
rect 1443 44353 1455 44387
rect 1397 44347 1455 44353
rect 2961 44387 3019 44393
rect 2961 44353 2973 44387
rect 3007 44353 3019 44387
rect 2961 44347 3019 44353
rect 3605 44387 3663 44393
rect 3605 44353 3617 44387
rect 3651 44384 3663 44387
rect 3786 44384 3792 44396
rect 3651 44356 3792 44384
rect 3651 44353 3663 44356
rect 3605 44347 3663 44353
rect 290 44276 296 44328
rect 348 44316 354 44328
rect 1412 44316 1440 44347
rect 348 44288 1440 44316
rect 2777 44319 2835 44325
rect 348 44276 354 44288
rect 2777 44285 2789 44319
rect 2823 44285 2835 44319
rect 2976 44316 3004 44347
rect 3786 44344 3792 44356
rect 3844 44344 3850 44396
rect 4246 44344 4252 44396
rect 4304 44384 4310 44396
rect 4709 44387 4767 44393
rect 4709 44384 4721 44387
rect 4304 44356 4721 44384
rect 4304 44344 4310 44356
rect 4709 44353 4721 44356
rect 4755 44384 4767 44387
rect 4890 44384 4896 44396
rect 4755 44356 4896 44384
rect 4755 44353 4767 44356
rect 4709 44347 4767 44353
rect 4890 44344 4896 44356
rect 4948 44384 4954 44396
rect 5626 44384 5632 44396
rect 4948 44356 5632 44384
rect 4948 44344 4954 44356
rect 5626 44344 5632 44356
rect 5684 44344 5690 44396
rect 9490 44344 9496 44396
rect 9548 44384 9554 44396
rect 9861 44387 9919 44393
rect 9861 44384 9873 44387
rect 9548 44356 9873 44384
rect 9548 44344 9554 44356
rect 9861 44353 9873 44356
rect 9907 44353 9919 44387
rect 9861 44347 9919 44353
rect 3878 44316 3884 44328
rect 2976 44288 3884 44316
rect 2777 44279 2835 44285
rect 2792 44248 2820 44279
rect 3878 44276 3884 44288
rect 3936 44276 3942 44328
rect 3970 44276 3976 44328
rect 4028 44316 4034 44328
rect 4525 44319 4583 44325
rect 4525 44316 4537 44319
rect 4028 44288 4537 44316
rect 4028 44276 4034 44288
rect 4525 44285 4537 44288
rect 4571 44285 4583 44319
rect 4525 44279 4583 44285
rect 2958 44248 2964 44260
rect 2792 44220 2964 44248
rect 2958 44208 2964 44220
rect 3016 44208 3022 44260
rect 3145 44251 3203 44257
rect 3145 44217 3157 44251
rect 3191 44248 3203 44251
rect 5166 44248 5172 44260
rect 3191 44220 5172 44248
rect 3191 44217 3203 44220
rect 3145 44211 3203 44217
rect 5166 44208 5172 44220
rect 5224 44208 5230 44260
rect 3786 44180 3792 44192
rect 3747 44152 3792 44180
rect 3786 44140 3792 44152
rect 3844 44140 3850 44192
rect 10042 44180 10048 44192
rect 10003 44152 10048 44180
rect 10042 44140 10048 44152
rect 10100 44140 10106 44192
rect 1104 44090 10856 44112
rect 1104 44038 2582 44090
rect 2634 44038 2646 44090
rect 2698 44038 2710 44090
rect 2762 44038 2774 44090
rect 2826 44038 2838 44090
rect 2890 44038 5846 44090
rect 5898 44038 5910 44090
rect 5962 44038 5974 44090
rect 6026 44038 6038 44090
rect 6090 44038 6102 44090
rect 6154 44038 9110 44090
rect 9162 44038 9174 44090
rect 9226 44038 9238 44090
rect 9290 44038 9302 44090
rect 9354 44038 9366 44090
rect 9418 44038 10856 44090
rect 1104 44016 10856 44038
rect 9217 43979 9275 43985
rect 1872 43948 5212 43976
rect 1872 43772 1900 43948
rect 2222 43868 2228 43920
rect 2280 43868 2286 43920
rect 2501 43911 2559 43917
rect 2501 43877 2513 43911
rect 2547 43908 2559 43911
rect 5184 43908 5212 43948
rect 9217 43945 9229 43979
rect 9263 43976 9275 43979
rect 9490 43976 9496 43988
rect 9263 43948 9496 43976
rect 9263 43945 9275 43948
rect 9217 43939 9275 43945
rect 9490 43936 9496 43948
rect 9548 43936 9554 43988
rect 9766 43908 9772 43920
rect 2547 43880 4660 43908
rect 5184 43880 9772 43908
rect 2547 43877 2559 43880
rect 2501 43871 2559 43877
rect 2130 43840 2136 43852
rect 2056 43812 2136 43840
rect 1949 43775 2007 43781
rect 1949 43772 1961 43775
rect 1872 43744 1961 43772
rect 1949 43741 1961 43744
rect 1995 43741 2007 43775
rect 1949 43735 2007 43741
rect 1486 43664 1492 43716
rect 1544 43704 1550 43716
rect 2056 43704 2084 43812
rect 2130 43800 2136 43812
rect 2188 43800 2194 43852
rect 2240 43781 2268 43868
rect 2866 43800 2872 43852
rect 2924 43840 2930 43852
rect 3142 43840 3148 43852
rect 2924 43812 3148 43840
rect 2924 43800 2930 43812
rect 3142 43800 3148 43812
rect 3200 43800 3206 43852
rect 2225 43775 2283 43781
rect 2225 43741 2237 43775
rect 2271 43741 2283 43775
rect 2225 43735 2283 43741
rect 2317 43775 2375 43781
rect 2317 43741 2329 43775
rect 2363 43772 2375 43775
rect 2498 43772 2504 43784
rect 2363 43744 2504 43772
rect 2363 43741 2375 43744
rect 2317 43735 2375 43741
rect 2498 43732 2504 43744
rect 2556 43732 2562 43784
rect 2961 43775 3019 43781
rect 2961 43741 2973 43775
rect 3007 43772 3019 43775
rect 3418 43772 3424 43784
rect 3007 43744 3424 43772
rect 3007 43741 3019 43744
rect 2961 43735 3019 43741
rect 3418 43732 3424 43744
rect 3476 43732 3482 43784
rect 3878 43772 3884 43784
rect 3839 43744 3884 43772
rect 3878 43732 3884 43744
rect 3936 43732 3942 43784
rect 3973 43775 4031 43781
rect 3973 43741 3985 43775
rect 4019 43772 4031 43775
rect 4246 43772 4252 43784
rect 4019 43744 4252 43772
rect 4019 43741 4031 43744
rect 3973 43735 4031 43741
rect 4246 43732 4252 43744
rect 4304 43732 4310 43784
rect 4632 43781 4660 43880
rect 9766 43868 9772 43880
rect 9824 43868 9830 43920
rect 4617 43775 4675 43781
rect 4617 43741 4629 43775
rect 4663 43741 4675 43775
rect 4617 43735 4675 43741
rect 9401 43775 9459 43781
rect 9401 43741 9413 43775
rect 9447 43741 9459 43775
rect 9401 43735 9459 43741
rect 9861 43775 9919 43781
rect 9861 43741 9873 43775
rect 9907 43772 9919 43775
rect 9950 43772 9956 43784
rect 9907 43744 9956 43772
rect 9907 43741 9919 43744
rect 9861 43735 9919 43741
rect 1544 43676 2084 43704
rect 2133 43707 2191 43713
rect 1544 43664 1550 43676
rect 2133 43673 2145 43707
rect 2179 43704 2191 43707
rect 2774 43704 2780 43716
rect 2179 43676 2780 43704
rect 2179 43673 2191 43676
rect 2133 43667 2191 43673
rect 2774 43664 2780 43676
rect 2832 43664 2838 43716
rect 4157 43707 4215 43713
rect 4157 43673 4169 43707
rect 4203 43704 4215 43707
rect 9416 43704 9444 43735
rect 9950 43732 9956 43744
rect 10008 43732 10014 43784
rect 4203 43676 9444 43704
rect 4203 43673 4215 43676
rect 4157 43667 4215 43673
rect 2222 43596 2228 43648
rect 2280 43636 2286 43648
rect 2958 43636 2964 43648
rect 2280 43608 2964 43636
rect 2280 43596 2286 43608
rect 2958 43596 2964 43608
rect 3016 43596 3022 43648
rect 3142 43636 3148 43648
rect 3103 43608 3148 43636
rect 3142 43596 3148 43608
rect 3200 43596 3206 43648
rect 3418 43596 3424 43648
rect 3476 43636 3482 43648
rect 4801 43639 4859 43645
rect 4801 43636 4813 43639
rect 3476 43608 4813 43636
rect 3476 43596 3482 43608
rect 4801 43605 4813 43608
rect 4847 43605 4859 43639
rect 10042 43636 10048 43648
rect 10003 43608 10048 43636
rect 4801 43599 4859 43605
rect 10042 43596 10048 43608
rect 10100 43596 10106 43648
rect 1104 43546 10856 43568
rect 1104 43494 4214 43546
rect 4266 43494 4278 43546
rect 4330 43494 4342 43546
rect 4394 43494 4406 43546
rect 4458 43494 4470 43546
rect 4522 43494 7478 43546
rect 7530 43494 7542 43546
rect 7594 43494 7606 43546
rect 7658 43494 7670 43546
rect 7722 43494 7734 43546
rect 7786 43494 10856 43546
rect 1104 43472 10856 43494
rect 1578 43432 1584 43444
rect 1539 43404 1584 43432
rect 1578 43392 1584 43404
rect 1636 43392 1642 43444
rect 9950 43432 9956 43444
rect 9911 43404 9956 43432
rect 9950 43392 9956 43404
rect 10008 43392 10014 43444
rect 2746 43336 3832 43364
rect 2746 43308 2774 43336
rect 1397 43299 1455 43305
rect 1397 43296 1409 43299
rect 1228 43268 1409 43296
rect 1228 43160 1256 43268
rect 1397 43265 1409 43268
rect 1443 43265 1455 43299
rect 1397 43259 1455 43265
rect 1486 43256 1492 43308
rect 1544 43296 1550 43308
rect 2133 43299 2191 43305
rect 2133 43296 2145 43299
rect 1544 43268 2145 43296
rect 1544 43256 1550 43268
rect 2133 43265 2145 43268
rect 2179 43265 2191 43299
rect 2498 43296 2504 43308
rect 2133 43259 2191 43265
rect 2424 43268 2504 43296
rect 2424 43240 2452 43268
rect 2498 43256 2504 43268
rect 2556 43256 2562 43308
rect 2682 43256 2688 43308
rect 2740 43268 2774 43308
rect 3804 43305 3832 43336
rect 2869 43299 2927 43305
rect 2740 43256 2746 43268
rect 2869 43265 2881 43299
rect 2915 43296 2927 43299
rect 3789 43299 3847 43305
rect 2915 43268 3556 43296
rect 2915 43265 2927 43268
rect 2869 43259 2927 43265
rect 1302 43188 1308 43240
rect 1360 43228 1366 43240
rect 1670 43228 1676 43240
rect 1360 43200 1676 43228
rect 1360 43188 1366 43200
rect 1670 43188 1676 43200
rect 1728 43188 1734 43240
rect 2406 43188 2412 43240
rect 2464 43188 2470 43240
rect 2774 43188 2780 43240
rect 2832 43228 2838 43240
rect 3145 43231 3203 43237
rect 3145 43228 3157 43231
rect 2832 43200 3157 43228
rect 2832 43188 2838 43200
rect 3145 43197 3157 43200
rect 3191 43228 3203 43231
rect 3418 43228 3424 43240
rect 3191 43200 3424 43228
rect 3191 43197 3203 43200
rect 3145 43191 3203 43197
rect 3418 43188 3424 43200
rect 3476 43188 3482 43240
rect 3528 43228 3556 43268
rect 3789 43265 3801 43299
rect 3835 43265 3847 43299
rect 10134 43296 10140 43308
rect 10095 43268 10140 43296
rect 3789 43259 3847 43265
rect 10134 43256 10140 43268
rect 10192 43256 10198 43308
rect 4154 43228 4160 43240
rect 3528 43200 4160 43228
rect 3804 43172 3832 43200
rect 4154 43188 4160 43200
rect 4212 43188 4218 43240
rect 1486 43160 1492 43172
rect 1228 43132 1492 43160
rect 1486 43120 1492 43132
rect 1544 43120 1550 43172
rect 3786 43120 3792 43172
rect 3844 43120 3850 43172
rect 2317 43095 2375 43101
rect 2317 43061 2329 43095
rect 2363 43092 2375 43095
rect 3050 43092 3056 43104
rect 2363 43064 3056 43092
rect 2363 43061 2375 43064
rect 2317 43055 2375 43061
rect 3050 43052 3056 43064
rect 3108 43052 3114 43104
rect 3970 43092 3976 43104
rect 3931 43064 3976 43092
rect 3970 43052 3976 43064
rect 4028 43052 4034 43104
rect 1104 43002 10856 43024
rect 1104 42950 2582 43002
rect 2634 42950 2646 43002
rect 2698 42950 2710 43002
rect 2762 42950 2774 43002
rect 2826 42950 2838 43002
rect 2890 42950 5846 43002
rect 5898 42950 5910 43002
rect 5962 42950 5974 43002
rect 6026 42950 6038 43002
rect 6090 42950 6102 43002
rect 6154 42950 9110 43002
rect 9162 42950 9174 43002
rect 9226 42950 9238 43002
rect 9290 42950 9302 43002
rect 9354 42950 9366 43002
rect 9418 42950 10856 43002
rect 1104 42928 10856 42950
rect 566 42780 572 42832
rect 624 42820 630 42832
rect 624 42792 1808 42820
rect 624 42780 630 42792
rect 1780 42761 1808 42792
rect 1765 42755 1823 42761
rect 1765 42721 1777 42755
rect 1811 42721 1823 42755
rect 1765 42715 1823 42721
rect 3142 42712 3148 42764
rect 3200 42752 3206 42764
rect 3510 42752 3516 42764
rect 3200 42724 3516 42752
rect 3200 42712 3206 42724
rect 3510 42712 3516 42724
rect 3568 42712 3574 42764
rect 1486 42684 1492 42696
rect 1447 42656 1492 42684
rect 1486 42644 1492 42656
rect 1544 42644 1550 42696
rect 2777 42687 2835 42693
rect 2777 42653 2789 42687
rect 2823 42684 2835 42687
rect 2958 42684 2964 42696
rect 2823 42656 2964 42684
rect 2823 42653 2835 42656
rect 2777 42647 2835 42653
rect 2958 42644 2964 42656
rect 3016 42644 3022 42696
rect 3786 42684 3792 42696
rect 3747 42656 3792 42684
rect 3786 42644 3792 42656
rect 3844 42644 3850 42696
rect 9766 42644 9772 42696
rect 9824 42684 9830 42696
rect 9861 42687 9919 42693
rect 9861 42684 9873 42687
rect 9824 42656 9873 42684
rect 9824 42644 9830 42656
rect 9861 42653 9873 42656
rect 9907 42653 9919 42687
rect 9861 42647 9919 42653
rect 2958 42548 2964 42560
rect 2919 42520 2964 42548
rect 2958 42508 2964 42520
rect 3016 42508 3022 42560
rect 3418 42508 3424 42560
rect 3476 42548 3482 42560
rect 3973 42551 4031 42557
rect 3973 42548 3985 42551
rect 3476 42520 3985 42548
rect 3476 42508 3482 42520
rect 3973 42517 3985 42520
rect 4019 42517 4031 42551
rect 10042 42548 10048 42560
rect 10003 42520 10048 42548
rect 3973 42511 4031 42517
rect 10042 42508 10048 42520
rect 10100 42508 10106 42560
rect 1104 42458 10856 42480
rect 1104 42406 4214 42458
rect 4266 42406 4278 42458
rect 4330 42406 4342 42458
rect 4394 42406 4406 42458
rect 4458 42406 4470 42458
rect 4522 42406 7478 42458
rect 7530 42406 7542 42458
rect 7594 42406 7606 42458
rect 7658 42406 7670 42458
rect 7722 42406 7734 42458
rect 7786 42406 10856 42458
rect 1104 42384 10856 42406
rect 1486 42304 1492 42356
rect 1544 42344 1550 42356
rect 3053 42347 3111 42353
rect 3053 42344 3065 42347
rect 1544 42316 3065 42344
rect 1544 42304 1550 42316
rect 3053 42313 3065 42316
rect 3099 42313 3111 42347
rect 3053 42307 3111 42313
rect 4249 42347 4307 42353
rect 4249 42313 4261 42347
rect 4295 42344 4307 42347
rect 10134 42344 10140 42356
rect 4295 42316 10140 42344
rect 4295 42313 4307 42316
rect 4249 42307 4307 42313
rect 10134 42304 10140 42316
rect 10192 42304 10198 42356
rect 1302 42236 1308 42288
rect 1360 42276 1366 42288
rect 1762 42276 1768 42288
rect 1360 42248 1768 42276
rect 1360 42236 1366 42248
rect 1762 42236 1768 42248
rect 1820 42236 1826 42288
rect 2682 42236 2688 42288
rect 2740 42276 2746 42288
rect 4430 42276 4436 42288
rect 2740 42248 2912 42276
rect 2740 42236 2746 42248
rect 1673 42211 1731 42217
rect 1673 42177 1685 42211
rect 1719 42208 1731 42211
rect 2774 42208 2780 42220
rect 1719 42180 2780 42208
rect 1719 42177 1731 42180
rect 1673 42171 1731 42177
rect 2774 42168 2780 42180
rect 2832 42168 2838 42220
rect 2884 42217 2912 42248
rect 4080 42248 4436 42276
rect 2869 42211 2927 42217
rect 2869 42177 2881 42211
rect 2915 42177 2927 42211
rect 3970 42208 3976 42220
rect 3931 42180 3976 42208
rect 2869 42171 2927 42177
rect 1394 42140 1400 42152
rect 1355 42112 1400 42140
rect 1394 42100 1400 42112
rect 1452 42100 1458 42152
rect 2222 42100 2228 42152
rect 2280 42100 2286 42152
rect 2685 42143 2743 42149
rect 2685 42109 2697 42143
rect 2731 42109 2743 42143
rect 2685 42103 2743 42109
rect 566 42032 572 42084
rect 624 42072 630 42084
rect 2240 42072 2268 42100
rect 2700 42072 2728 42103
rect 624 42044 2728 42072
rect 624 42032 630 42044
rect 2222 41964 2228 42016
rect 2280 42004 2286 42016
rect 2884 42004 2912 42171
rect 3970 42168 3976 42180
rect 4028 42168 4034 42220
rect 4080 42217 4108 42248
rect 4430 42236 4436 42248
rect 4488 42276 4494 42288
rect 4890 42276 4896 42288
rect 4488 42248 4896 42276
rect 4488 42236 4494 42248
rect 4890 42236 4896 42248
rect 4948 42236 4954 42288
rect 4065 42211 4123 42217
rect 4065 42177 4077 42211
rect 4111 42177 4123 42211
rect 4065 42171 4123 42177
rect 4709 42211 4767 42217
rect 4709 42177 4721 42211
rect 4755 42208 4767 42211
rect 5258 42208 5264 42220
rect 4755 42180 5264 42208
rect 4755 42177 4767 42180
rect 4709 42171 4767 42177
rect 5258 42168 5264 42180
rect 5316 42168 5322 42220
rect 5626 42208 5632 42220
rect 5587 42180 5632 42208
rect 5626 42168 5632 42180
rect 5684 42168 5690 42220
rect 9490 42168 9496 42220
rect 9548 42208 9554 42220
rect 9861 42211 9919 42217
rect 9861 42208 9873 42211
rect 9548 42180 9873 42208
rect 9548 42168 9554 42180
rect 9861 42177 9873 42180
rect 9907 42177 9919 42211
rect 9861 42171 9919 42177
rect 3786 42032 3792 42084
rect 3844 42072 3850 42084
rect 4893 42075 4951 42081
rect 4893 42072 4905 42075
rect 3844 42044 4905 42072
rect 3844 42032 3850 42044
rect 4893 42041 4905 42044
rect 4939 42041 4951 42075
rect 4893 42035 4951 42041
rect 5445 42075 5503 42081
rect 5445 42041 5457 42075
rect 5491 42072 5503 42075
rect 8294 42072 8300 42084
rect 5491 42044 8300 42072
rect 5491 42041 5503 42044
rect 5445 42035 5503 42041
rect 8294 42032 8300 42044
rect 8352 42032 8358 42084
rect 10042 42004 10048 42016
rect 2280 41976 2912 42004
rect 10003 41976 10048 42004
rect 2280 41964 2286 41976
rect 10042 41964 10048 41976
rect 10100 41964 10106 42016
rect 1104 41914 10856 41936
rect 1104 41862 2582 41914
rect 2634 41862 2646 41914
rect 2698 41862 2710 41914
rect 2762 41862 2774 41914
rect 2826 41862 2838 41914
rect 2890 41862 5846 41914
rect 5898 41862 5910 41914
rect 5962 41862 5974 41914
rect 6026 41862 6038 41914
rect 6090 41862 6102 41914
rect 6154 41862 9110 41914
rect 9162 41862 9174 41914
rect 9226 41862 9238 41914
rect 9290 41862 9302 41914
rect 9354 41862 9366 41914
rect 9418 41862 10856 41914
rect 1104 41840 10856 41862
rect 4617 41803 4675 41809
rect 4617 41769 4629 41803
rect 4663 41800 4675 41803
rect 5626 41800 5632 41812
rect 4663 41772 5632 41800
rect 4663 41769 4675 41772
rect 4617 41763 4675 41769
rect 5626 41760 5632 41772
rect 5684 41760 5690 41812
rect 2774 41732 2780 41744
rect 1780 41704 2780 41732
rect 1780 41673 1808 41704
rect 2774 41692 2780 41704
rect 2832 41692 2838 41744
rect 1765 41667 1823 41673
rect 1765 41633 1777 41667
rect 1811 41633 1823 41667
rect 1765 41627 1823 41633
rect 4154 41624 4160 41676
rect 4212 41664 4218 41676
rect 4249 41667 4307 41673
rect 4249 41664 4261 41667
rect 4212 41636 4261 41664
rect 4212 41624 4218 41636
rect 4249 41633 4261 41636
rect 4295 41664 4307 41667
rect 5258 41664 5264 41676
rect 4295 41636 5264 41664
rect 4295 41633 4307 41636
rect 4249 41627 4307 41633
rect 5258 41624 5264 41636
rect 5316 41624 5322 41676
rect 1302 41556 1308 41608
rect 1360 41596 1366 41608
rect 2041 41599 2099 41605
rect 2041 41596 2053 41599
rect 1360 41568 2053 41596
rect 1360 41556 1366 41568
rect 2041 41565 2053 41568
rect 2087 41565 2099 41599
rect 2041 41559 2099 41565
rect 3418 41556 3424 41608
rect 3476 41596 3482 41608
rect 4062 41596 4068 41608
rect 3476 41568 4068 41596
rect 3476 41556 3482 41568
rect 4062 41556 4068 41568
rect 4120 41556 4126 41608
rect 4430 41596 4436 41608
rect 4391 41568 4436 41596
rect 4430 41556 4436 41568
rect 4488 41596 4494 41608
rect 5074 41596 5080 41608
rect 4488 41568 5080 41596
rect 4488 41556 4494 41568
rect 5074 41556 5080 41568
rect 5132 41556 5138 41608
rect 1026 41488 1032 41540
rect 1084 41528 1090 41540
rect 1084 41500 1440 41528
rect 1084 41488 1090 41500
rect 1412 41460 1440 41500
rect 1946 41488 1952 41540
rect 2004 41528 2010 41540
rect 2682 41528 2688 41540
rect 2004 41500 2688 41528
rect 2004 41488 2010 41500
rect 2682 41488 2688 41500
rect 2740 41488 2746 41540
rect 3786 41528 3792 41540
rect 3528 41500 3792 41528
rect 3528 41472 3556 41500
rect 3786 41488 3792 41500
rect 3844 41488 3850 41540
rect 1762 41460 1768 41472
rect 1412 41432 1768 41460
rect 1762 41420 1768 41432
rect 1820 41420 1826 41472
rect 3510 41420 3516 41472
rect 3568 41420 3574 41472
rect 1104 41370 10856 41392
rect 1104 41318 4214 41370
rect 4266 41318 4278 41370
rect 4330 41318 4342 41370
rect 4394 41318 4406 41370
rect 4458 41318 4470 41370
rect 4522 41318 7478 41370
rect 7530 41318 7542 41370
rect 7594 41318 7606 41370
rect 7658 41318 7670 41370
rect 7722 41318 7734 41370
rect 7786 41318 10856 41370
rect 1104 41296 10856 41318
rect 1394 41216 1400 41268
rect 1452 41256 1458 41268
rect 1949 41259 2007 41265
rect 1949 41256 1961 41259
rect 1452 41228 1961 41256
rect 1452 41216 1458 41228
rect 1949 41225 1961 41228
rect 1995 41225 2007 41259
rect 1949 41219 2007 41225
rect 2406 41216 2412 41268
rect 2464 41256 2470 41268
rect 2590 41256 2596 41268
rect 2464 41228 2596 41256
rect 2464 41216 2470 41228
rect 2590 41216 2596 41228
rect 2648 41216 2654 41268
rect 2774 41256 2780 41268
rect 2735 41228 2780 41256
rect 2774 41216 2780 41228
rect 2832 41216 2838 41268
rect 3510 41216 3516 41268
rect 3568 41256 3574 41268
rect 3568 41228 3924 41256
rect 3568 41216 3574 41228
rect 3896 41200 3924 41228
rect 6178 41216 6184 41268
rect 6236 41216 6242 41268
rect 1118 41148 1124 41200
rect 1176 41188 1182 41200
rect 1670 41188 1676 41200
rect 1176 41160 1676 41188
rect 1176 41148 1182 41160
rect 1670 41148 1676 41160
rect 1728 41148 1734 41200
rect 3878 41148 3884 41200
rect 3936 41148 3942 41200
rect 4338 41148 4344 41200
rect 4396 41188 4402 41200
rect 6196 41188 6224 41216
rect 4396 41160 6224 41188
rect 4396 41148 4402 41160
rect 1394 41080 1400 41132
rect 1452 41120 1458 41132
rect 1765 41123 1823 41129
rect 1452 41092 1716 41120
rect 1452 41080 1458 41092
rect 1581 41055 1639 41061
rect 1581 41021 1593 41055
rect 1627 41021 1639 41055
rect 1688 41052 1716 41092
rect 1765 41089 1777 41123
rect 1811 41120 1823 41123
rect 1946 41120 1952 41132
rect 1811 41092 1952 41120
rect 1811 41089 1823 41092
rect 1765 41083 1823 41089
rect 1946 41080 1952 41092
rect 2004 41120 2010 41132
rect 2222 41120 2228 41132
rect 2004 41092 2228 41120
rect 2004 41080 2010 41092
rect 2222 41080 2228 41092
rect 2280 41120 2286 41132
rect 2593 41123 2651 41129
rect 2593 41120 2605 41123
rect 2280 41092 2605 41120
rect 2280 41080 2286 41092
rect 2593 41089 2605 41092
rect 2639 41089 2651 41123
rect 2593 41083 2651 41089
rect 2682 41080 2688 41132
rect 2740 41120 2746 41132
rect 3237 41123 3295 41129
rect 3237 41120 3249 41123
rect 2740 41092 3249 41120
rect 2740 41080 2746 41092
rect 3237 41089 3249 41092
rect 3283 41089 3295 41123
rect 4522 41120 4528 41132
rect 4435 41092 4528 41120
rect 3237 41083 3295 41089
rect 4522 41080 4528 41092
rect 4580 41120 4586 41132
rect 4709 41123 4767 41129
rect 4580 41092 4660 41120
rect 4580 41080 4586 41092
rect 2409 41055 2467 41061
rect 2409 41052 2421 41055
rect 1688 41024 2421 41052
rect 1581 41015 1639 41021
rect 2409 41021 2421 41024
rect 2455 41052 2467 41055
rect 4341 41055 4399 41061
rect 4341 41052 4353 41055
rect 2455 41024 4353 41052
rect 2455 41021 2467 41024
rect 2409 41015 2467 41021
rect 4341 41021 4353 41024
rect 4387 41021 4399 41055
rect 4632 41052 4660 41092
rect 4709 41089 4721 41123
rect 4755 41120 4767 41123
rect 5721 41123 5779 41129
rect 5721 41120 5733 41123
rect 4755 41092 5733 41120
rect 4755 41089 4767 41092
rect 4709 41083 4767 41089
rect 5721 41089 5733 41092
rect 5767 41089 5779 41123
rect 5721 41083 5779 41089
rect 6178 41080 6184 41132
rect 6236 41120 6242 41132
rect 9861 41123 9919 41129
rect 9861 41120 9873 41123
rect 6236 41092 9873 41120
rect 6236 41080 6242 41092
rect 9861 41089 9873 41092
rect 9907 41089 9919 41123
rect 9861 41083 9919 41089
rect 5074 41052 5080 41064
rect 4632 41024 5080 41052
rect 4341 41015 4399 41021
rect 1596 40984 1624 41015
rect 5074 41012 5080 41024
rect 5132 41012 5138 41064
rect 5350 41012 5356 41064
rect 5408 41052 5414 41064
rect 5626 41052 5632 41064
rect 5408 41024 5632 41052
rect 5408 41012 5414 41024
rect 5626 41012 5632 41024
rect 5684 41012 5690 41064
rect 4062 40984 4068 40996
rect 1596 40956 4068 40984
rect 4062 40944 4068 40956
rect 4120 40944 4126 40996
rect 5537 40987 5595 40993
rect 5537 40953 5549 40987
rect 5583 40984 5595 40987
rect 9858 40984 9864 40996
rect 5583 40956 9864 40984
rect 5583 40953 5595 40956
rect 5537 40947 5595 40953
rect 9858 40944 9864 40956
rect 9916 40944 9922 40996
rect 10042 40984 10048 40996
rect 10003 40956 10048 40984
rect 10042 40944 10048 40956
rect 10100 40944 10106 40996
rect 3418 40916 3424 40928
rect 3379 40888 3424 40916
rect 3418 40876 3424 40888
rect 3476 40876 3482 40928
rect 5074 40876 5080 40928
rect 5132 40916 5138 40928
rect 7282 40916 7288 40928
rect 5132 40888 7288 40916
rect 5132 40876 5138 40888
rect 7282 40876 7288 40888
rect 7340 40876 7346 40928
rect 1104 40826 10856 40848
rect 1104 40774 2582 40826
rect 2634 40774 2646 40826
rect 2698 40774 2710 40826
rect 2762 40774 2774 40826
rect 2826 40774 2838 40826
rect 2890 40774 5846 40826
rect 5898 40774 5910 40826
rect 5962 40774 5974 40826
rect 6026 40774 6038 40826
rect 6090 40774 6102 40826
rect 6154 40774 9110 40826
rect 9162 40774 9174 40826
rect 9226 40774 9238 40826
rect 9290 40774 9302 40826
rect 9354 40774 9366 40826
rect 9418 40774 10856 40826
rect 1104 40752 10856 40774
rect 3786 40672 3792 40724
rect 3844 40712 3850 40724
rect 4062 40712 4068 40724
rect 3844 40684 4068 40712
rect 3844 40672 3850 40684
rect 4062 40672 4068 40684
rect 4120 40672 4126 40724
rect 9217 40715 9275 40721
rect 9217 40681 9229 40715
rect 9263 40712 9275 40715
rect 9490 40712 9496 40724
rect 9263 40684 9496 40712
rect 9263 40681 9275 40684
rect 9217 40675 9275 40681
rect 9490 40672 9496 40684
rect 9548 40672 9554 40724
rect 2222 40604 2228 40656
rect 2280 40644 2286 40656
rect 3970 40644 3976 40656
rect 2280 40616 3976 40644
rect 2280 40604 2286 40616
rect 3970 40604 3976 40616
rect 4028 40604 4034 40656
rect 4706 40604 4712 40656
rect 4764 40644 4770 40656
rect 5626 40644 5632 40656
rect 4764 40616 5632 40644
rect 4764 40604 4770 40616
rect 5626 40604 5632 40616
rect 5684 40604 5690 40656
rect 14 40536 20 40588
rect 72 40576 78 40588
rect 2317 40579 2375 40585
rect 2317 40576 2329 40579
rect 72 40548 2329 40576
rect 72 40536 78 40548
rect 2317 40545 2329 40548
rect 2363 40545 2375 40579
rect 2317 40539 2375 40545
rect 2041 40511 2099 40517
rect 2041 40477 2053 40511
rect 2087 40477 2099 40511
rect 2041 40471 2099 40477
rect 3789 40511 3847 40517
rect 3789 40477 3801 40511
rect 3835 40508 3847 40511
rect 4338 40508 4344 40520
rect 3835 40480 4344 40508
rect 3835 40477 3847 40480
rect 3789 40471 3847 40477
rect 14 40400 20 40452
rect 72 40440 78 40452
rect 566 40440 572 40452
rect 72 40412 572 40440
rect 72 40400 78 40412
rect 566 40400 572 40412
rect 624 40400 630 40452
rect 2056 40372 2084 40471
rect 4338 40468 4344 40480
rect 4396 40468 4402 40520
rect 4982 40468 4988 40520
rect 5040 40508 5046 40520
rect 9401 40511 9459 40517
rect 9401 40508 9413 40511
rect 5040 40480 9413 40508
rect 5040 40468 5046 40480
rect 9401 40477 9413 40480
rect 9447 40477 9459 40511
rect 9858 40508 9864 40520
rect 9819 40480 9864 40508
rect 9401 40471 9459 40477
rect 9858 40468 9864 40480
rect 9916 40468 9922 40520
rect 4522 40400 4528 40452
rect 4580 40440 4586 40452
rect 4706 40440 4712 40452
rect 4580 40412 4712 40440
rect 4580 40400 4586 40412
rect 4706 40400 4712 40412
rect 4764 40400 4770 40452
rect 3142 40372 3148 40384
rect 2056 40344 3148 40372
rect 3142 40332 3148 40344
rect 3200 40332 3206 40384
rect 3234 40332 3240 40384
rect 3292 40372 3298 40384
rect 3418 40372 3424 40384
rect 3292 40344 3424 40372
rect 3292 40332 3298 40344
rect 3418 40332 3424 40344
rect 3476 40332 3482 40384
rect 3970 40372 3976 40384
rect 3931 40344 3976 40372
rect 3970 40332 3976 40344
rect 4028 40332 4034 40384
rect 10042 40372 10048 40384
rect 10003 40344 10048 40372
rect 10042 40332 10048 40344
rect 10100 40332 10106 40384
rect 1104 40282 10856 40304
rect 1104 40230 4214 40282
rect 4266 40230 4278 40282
rect 4330 40230 4342 40282
rect 4394 40230 4406 40282
rect 4458 40230 4470 40282
rect 4522 40230 7478 40282
rect 7530 40230 7542 40282
rect 7594 40230 7606 40282
rect 7658 40230 7670 40282
rect 7722 40230 7734 40282
rect 7786 40230 10856 40282
rect 1104 40208 10856 40230
rect 2222 40168 2228 40180
rect 1688 40140 2228 40168
rect 1688 40041 1716 40140
rect 2222 40128 2228 40140
rect 2280 40128 2286 40180
rect 6365 40171 6423 40177
rect 3712 40140 6316 40168
rect 1946 40100 1952 40112
rect 1780 40072 1952 40100
rect 1780 40041 1808 40072
rect 1946 40060 1952 40072
rect 2004 40100 2010 40112
rect 2958 40100 2964 40112
rect 2004 40072 2964 40100
rect 2004 40060 2010 40072
rect 2958 40060 2964 40072
rect 3016 40060 3022 40112
rect 3712 40041 3740 40140
rect 4338 40060 4344 40112
rect 4396 40100 4402 40112
rect 4706 40100 4712 40112
rect 4396 40072 4712 40100
rect 4396 40060 4402 40072
rect 4706 40060 4712 40072
rect 4764 40060 4770 40112
rect 6288 40100 6316 40140
rect 6365 40137 6377 40171
rect 6411 40168 6423 40171
rect 9858 40168 9864 40180
rect 6411 40140 9864 40168
rect 6411 40137 6423 40140
rect 6365 40131 6423 40137
rect 9858 40128 9864 40140
rect 9916 40128 9922 40180
rect 6638 40100 6644 40112
rect 6288 40072 6644 40100
rect 6638 40060 6644 40072
rect 6696 40060 6702 40112
rect 1673 40035 1731 40041
rect 1673 40001 1685 40035
rect 1719 40001 1731 40035
rect 1673 39995 1731 40001
rect 1765 40035 1823 40041
rect 1765 40001 1777 40035
rect 1811 40001 1823 40035
rect 1765 39995 1823 40001
rect 3697 40035 3755 40041
rect 3697 40001 3709 40035
rect 3743 40001 3755 40035
rect 3697 39995 3755 40001
rect 4433 40035 4491 40041
rect 4433 40001 4445 40035
rect 4479 40032 4491 40035
rect 5718 40032 5724 40044
rect 4479 40004 5724 40032
rect 4479 40001 4491 40004
rect 4433 39995 4491 40001
rect 5718 39992 5724 40004
rect 5776 39992 5782 40044
rect 6546 40032 6552 40044
rect 6507 40004 6552 40032
rect 6546 39992 6552 40004
rect 6604 39992 6610 40044
rect 9858 40032 9864 40044
rect 9819 40004 9864 40032
rect 9858 39992 9864 40004
rect 9916 39992 9922 40044
rect 1949 39967 2007 39973
rect 1949 39933 1961 39967
rect 1995 39964 2007 39967
rect 2409 39967 2467 39973
rect 2409 39964 2421 39967
rect 1995 39936 2421 39964
rect 1995 39933 2007 39936
rect 1949 39927 2007 39933
rect 2409 39933 2421 39936
rect 2455 39933 2467 39967
rect 2409 39927 2467 39933
rect 2590 39924 2596 39976
rect 2648 39964 2654 39976
rect 2685 39967 2743 39973
rect 2685 39964 2697 39967
rect 2648 39936 2697 39964
rect 2648 39924 2654 39936
rect 2685 39933 2697 39936
rect 2731 39933 2743 39967
rect 2685 39927 2743 39933
rect 3326 39856 3332 39908
rect 3384 39896 3390 39908
rect 4617 39899 4675 39905
rect 4617 39896 4629 39899
rect 3384 39868 4629 39896
rect 3384 39856 3390 39868
rect 4617 39865 4629 39868
rect 4663 39865 4675 39899
rect 4617 39859 4675 39865
rect 3881 39831 3939 39837
rect 3881 39797 3893 39831
rect 3927 39828 3939 39831
rect 4246 39828 4252 39840
rect 3927 39800 4252 39828
rect 3927 39797 3939 39800
rect 3881 39791 3939 39797
rect 4246 39788 4252 39800
rect 4304 39788 4310 39840
rect 10042 39828 10048 39840
rect 10003 39800 10048 39828
rect 10042 39788 10048 39800
rect 10100 39788 10106 39840
rect 1104 39738 10856 39760
rect 1104 39686 2582 39738
rect 2634 39686 2646 39738
rect 2698 39686 2710 39738
rect 2762 39686 2774 39738
rect 2826 39686 2838 39738
rect 2890 39686 5846 39738
rect 5898 39686 5910 39738
rect 5962 39686 5974 39738
rect 6026 39686 6038 39738
rect 6090 39686 6102 39738
rect 6154 39686 9110 39738
rect 9162 39686 9174 39738
rect 9226 39686 9238 39738
rect 9290 39686 9302 39738
rect 9354 39686 9366 39738
rect 9418 39686 10856 39738
rect 1104 39664 10856 39686
rect 3142 39624 3148 39636
rect 3103 39596 3148 39624
rect 3142 39584 3148 39596
rect 3200 39584 3206 39636
rect 5353 39627 5411 39633
rect 5353 39593 5365 39627
rect 5399 39624 5411 39627
rect 6178 39624 6184 39636
rect 5399 39596 6184 39624
rect 5399 39593 5411 39596
rect 5353 39587 5411 39593
rect 6178 39584 6184 39596
rect 6236 39584 6242 39636
rect 9766 39584 9772 39636
rect 9824 39624 9830 39636
rect 9953 39627 10011 39633
rect 9953 39624 9965 39627
rect 9824 39596 9965 39624
rect 9824 39584 9830 39596
rect 9953 39593 9965 39596
rect 9999 39593 10011 39627
rect 9953 39587 10011 39593
rect 2222 39516 2228 39568
rect 2280 39556 2286 39568
rect 3326 39556 3332 39568
rect 2280 39528 3332 39556
rect 2280 39516 2286 39528
rect 3326 39516 3332 39528
rect 3384 39516 3390 39568
rect 3786 39516 3792 39568
rect 3844 39556 3850 39568
rect 4801 39559 4859 39565
rect 4801 39556 4813 39559
rect 3844 39528 4813 39556
rect 3844 39516 3850 39528
rect 4801 39525 4813 39528
rect 4847 39525 4859 39559
rect 4801 39519 4859 39525
rect 1489 39491 1547 39497
rect 1489 39488 1501 39491
rect 1044 39460 1501 39488
rect 1044 39080 1072 39460
rect 1489 39457 1501 39460
rect 1535 39457 1547 39491
rect 5718 39488 5724 39500
rect 1489 39451 1547 39457
rect 4356 39460 5724 39488
rect 4356 39432 4384 39460
rect 5718 39448 5724 39460
rect 5776 39448 5782 39500
rect 1118 39380 1124 39432
rect 1176 39420 1182 39432
rect 1765 39423 1823 39429
rect 1765 39420 1777 39423
rect 1176 39392 1777 39420
rect 1176 39380 1182 39392
rect 1765 39389 1777 39392
rect 1811 39389 1823 39423
rect 1765 39383 1823 39389
rect 2774 39380 2780 39432
rect 2832 39420 2838 39432
rect 2832 39392 2877 39420
rect 2832 39380 2838 39392
rect 2958 39380 2964 39432
rect 3016 39420 3022 39432
rect 3789 39423 3847 39429
rect 3016 39392 3061 39420
rect 3016 39380 3022 39392
rect 3789 39389 3801 39423
rect 3835 39389 3847 39423
rect 3789 39383 3847 39389
rect 3973 39423 4031 39429
rect 3973 39389 3985 39423
rect 4019 39420 4031 39423
rect 4338 39420 4344 39432
rect 4019 39392 4344 39420
rect 4019 39389 4031 39392
rect 3973 39383 4031 39389
rect 2498 39312 2504 39364
rect 2556 39352 2562 39364
rect 3804 39352 3832 39383
rect 4338 39380 4344 39392
rect 4396 39380 4402 39432
rect 4614 39420 4620 39432
rect 4575 39392 4620 39420
rect 4614 39380 4620 39392
rect 4672 39380 4678 39432
rect 5534 39420 5540 39432
rect 5495 39392 5540 39420
rect 5534 39380 5540 39392
rect 5592 39380 5598 39432
rect 10137 39423 10195 39429
rect 10137 39389 10149 39423
rect 10183 39389 10195 39423
rect 10137 39383 10195 39389
rect 2556 39324 3832 39352
rect 4157 39355 4215 39361
rect 2556 39312 2562 39324
rect 4157 39321 4169 39355
rect 4203 39352 4215 39355
rect 10152 39352 10180 39383
rect 4203 39324 10180 39352
rect 4203 39321 4215 39324
rect 4157 39315 4215 39321
rect 1104 39194 10856 39216
rect 1104 39142 4214 39194
rect 4266 39142 4278 39194
rect 4330 39142 4342 39194
rect 4394 39142 4406 39194
rect 4458 39142 4470 39194
rect 4522 39142 7478 39194
rect 7530 39142 7542 39194
rect 7594 39142 7606 39194
rect 7658 39142 7670 39194
rect 7722 39142 7734 39194
rect 7786 39142 10856 39194
rect 1104 39120 10856 39142
rect 1118 39080 1124 39092
rect 1044 39052 1124 39080
rect 1118 39040 1124 39052
rect 1176 39040 1182 39092
rect 1762 39040 1768 39092
rect 1820 39080 1826 39092
rect 1946 39080 1952 39092
rect 1820 39052 1952 39080
rect 1820 39040 1826 39052
rect 1946 39040 1952 39052
rect 2004 39040 2010 39092
rect 5077 39083 5135 39089
rect 5077 39049 5089 39083
rect 5123 39080 5135 39083
rect 6546 39080 6552 39092
rect 5123 39052 6552 39080
rect 5123 39049 5135 39052
rect 5077 39043 5135 39049
rect 6546 39040 6552 39052
rect 6604 39040 6610 39092
rect 3234 38972 3240 39024
rect 3292 38972 3298 39024
rect 3786 38972 3792 39024
rect 3844 39012 3850 39024
rect 5626 39012 5632 39024
rect 3844 38984 5632 39012
rect 3844 38972 3850 38984
rect 5626 38972 5632 38984
rect 5684 38972 5690 39024
rect 934 38904 940 38956
rect 992 38944 998 38956
rect 1765 38947 1823 38953
rect 1765 38944 1777 38947
rect 992 38916 1777 38944
rect 992 38904 998 38916
rect 1765 38913 1777 38916
rect 1811 38913 1823 38947
rect 1765 38907 1823 38913
rect 3053 38947 3111 38953
rect 3053 38913 3065 38947
rect 3099 38944 3111 38947
rect 3252 38944 3280 38972
rect 3099 38916 3280 38944
rect 3099 38913 3111 38916
rect 3053 38907 3111 38913
rect 4430 38904 4436 38956
rect 4488 38944 4494 38956
rect 4893 38947 4951 38953
rect 4893 38944 4905 38947
rect 4488 38916 4905 38944
rect 4488 38904 4494 38916
rect 4893 38913 4905 38916
rect 4939 38944 4951 38947
rect 5718 38944 5724 38956
rect 4939 38916 5724 38944
rect 4939 38913 4951 38916
rect 4893 38907 4951 38913
rect 5718 38904 5724 38916
rect 5776 38904 5782 38956
rect 9674 38904 9680 38956
rect 9732 38944 9738 38956
rect 9861 38947 9919 38953
rect 9861 38944 9873 38947
rect 9732 38916 9873 38944
rect 9732 38904 9738 38916
rect 9861 38913 9873 38916
rect 9907 38913 9919 38947
rect 9861 38907 9919 38913
rect 1489 38879 1547 38885
rect 1489 38845 1501 38879
rect 1535 38876 1547 38879
rect 1670 38876 1676 38888
rect 1535 38848 1676 38876
rect 1535 38845 1547 38848
rect 1489 38839 1547 38845
rect 1670 38836 1676 38848
rect 1728 38836 1734 38888
rect 2777 38879 2835 38885
rect 2777 38845 2789 38879
rect 2823 38845 2835 38879
rect 2777 38839 2835 38845
rect 2792 38808 2820 38839
rect 2958 38836 2964 38888
rect 3016 38876 3022 38888
rect 3016 38848 4108 38876
rect 3016 38836 3022 38848
rect 3050 38808 3056 38820
rect 2792 38780 3056 38808
rect 3050 38768 3056 38780
rect 3108 38768 3114 38820
rect 4080 38808 4108 38848
rect 4154 38836 4160 38888
rect 4212 38876 4218 38888
rect 4709 38879 4767 38885
rect 4709 38876 4721 38879
rect 4212 38848 4721 38876
rect 4212 38836 4218 38848
rect 4709 38845 4721 38848
rect 4755 38845 4767 38879
rect 4709 38839 4767 38845
rect 4246 38808 4252 38820
rect 4080 38780 4252 38808
rect 4246 38768 4252 38780
rect 4304 38768 4310 38820
rect 10042 38740 10048 38752
rect 10003 38712 10048 38740
rect 10042 38700 10048 38712
rect 10100 38700 10106 38752
rect 1104 38650 10856 38672
rect 1104 38598 2582 38650
rect 2634 38598 2646 38650
rect 2698 38598 2710 38650
rect 2762 38598 2774 38650
rect 2826 38598 2838 38650
rect 2890 38598 5846 38650
rect 5898 38598 5910 38650
rect 5962 38598 5974 38650
rect 6026 38598 6038 38650
rect 6090 38598 6102 38650
rect 6154 38598 9110 38650
rect 9162 38598 9174 38650
rect 9226 38598 9238 38650
rect 9290 38598 9302 38650
rect 9354 38598 9366 38650
rect 9418 38598 10856 38650
rect 1104 38576 10856 38598
rect 566 38496 572 38548
rect 624 38536 630 38548
rect 1394 38536 1400 38548
rect 624 38508 1400 38536
rect 624 38496 630 38508
rect 1394 38496 1400 38508
rect 1452 38496 1458 38548
rect 1486 38496 1492 38548
rect 1544 38496 1550 38548
rect 1670 38496 1676 38548
rect 1728 38496 1734 38548
rect 1762 38496 1768 38548
rect 1820 38536 1826 38548
rect 1820 38508 1900 38536
rect 1820 38496 1826 38508
rect 934 38360 940 38412
rect 992 38400 998 38412
rect 1302 38400 1308 38412
rect 992 38372 1308 38400
rect 992 38360 998 38372
rect 1302 38360 1308 38372
rect 1360 38360 1366 38412
rect 1118 38332 1124 38344
rect 768 38304 1124 38332
rect 768 37924 796 38304
rect 1118 38292 1124 38304
rect 1176 38292 1182 38344
rect 1397 38335 1455 38341
rect 1397 38301 1409 38335
rect 1443 38332 1455 38335
rect 1504 38332 1532 38496
rect 1688 38412 1716 38496
rect 1670 38360 1676 38412
rect 1728 38360 1734 38412
rect 1872 38400 1900 38508
rect 1946 38496 1952 38548
rect 2004 38496 2010 38548
rect 2038 38496 2044 38548
rect 2096 38496 2102 38548
rect 2130 38496 2136 38548
rect 2188 38496 2194 38548
rect 2222 38496 2228 38548
rect 2280 38496 2286 38548
rect 2869 38539 2927 38545
rect 2869 38505 2881 38539
rect 2915 38536 2927 38539
rect 2958 38536 2964 38548
rect 2915 38508 2964 38536
rect 2915 38505 2927 38508
rect 2869 38499 2927 38505
rect 2958 38496 2964 38508
rect 3016 38496 3022 38548
rect 3142 38536 3148 38548
rect 3068 38508 3148 38536
rect 1964 38412 1992 38496
rect 1780 38372 1900 38400
rect 1780 38344 1808 38372
rect 1946 38360 1952 38412
rect 2004 38360 2010 38412
rect 1443 38304 1532 38332
rect 1443 38301 1455 38304
rect 1397 38295 1455 38301
rect 1762 38292 1768 38344
rect 1820 38292 1826 38344
rect 1854 38264 1860 38276
rect 860 38236 1860 38264
rect 860 38128 888 38236
rect 1854 38224 1860 38236
rect 1912 38224 1918 38276
rect 2056 38208 2084 38496
rect 2148 38276 2176 38496
rect 2130 38224 2136 38276
rect 2188 38224 2194 38276
rect 2240 38208 2268 38496
rect 3068 38480 3096 38508
rect 3142 38496 3148 38508
rect 3200 38496 3206 38548
rect 4617 38539 4675 38545
rect 4617 38505 4629 38539
rect 4663 38536 4675 38539
rect 5534 38536 5540 38548
rect 4663 38508 5540 38536
rect 4663 38505 4675 38508
rect 4617 38499 4675 38505
rect 5534 38496 5540 38508
rect 5592 38496 5598 38548
rect 3050 38428 3056 38480
rect 3108 38428 3114 38480
rect 4246 38428 4252 38480
rect 4304 38428 4310 38480
rect 4264 38400 4292 38428
rect 2516 38372 4292 38400
rect 2516 38344 2544 38372
rect 2498 38292 2504 38344
rect 2556 38292 2562 38344
rect 2700 38341 2728 38372
rect 2593 38335 2651 38341
rect 2593 38301 2605 38335
rect 2639 38301 2651 38335
rect 2593 38295 2651 38301
rect 2685 38335 2743 38341
rect 2685 38301 2697 38335
rect 2731 38301 2743 38335
rect 2685 38295 2743 38301
rect 4249 38335 4307 38341
rect 4249 38301 4261 38335
rect 4295 38301 4307 38335
rect 4430 38332 4436 38344
rect 4391 38304 4436 38332
rect 4249 38295 4307 38301
rect 2314 38224 2320 38276
rect 2372 38264 2378 38276
rect 2608 38264 2636 38295
rect 2372 38236 2636 38264
rect 2372 38224 2378 38236
rect 2958 38224 2964 38276
rect 3016 38264 3022 38276
rect 4154 38264 4160 38276
rect 3016 38236 4160 38264
rect 3016 38224 3022 38236
rect 4154 38224 4160 38236
rect 4212 38224 4218 38276
rect 934 38156 940 38208
rect 992 38196 998 38208
rect 1581 38199 1639 38205
rect 1581 38196 1593 38199
rect 992 38168 1593 38196
rect 992 38156 998 38168
rect 1581 38165 1593 38168
rect 1627 38165 1639 38199
rect 1581 38159 1639 38165
rect 2038 38156 2044 38208
rect 2096 38156 2102 38208
rect 2222 38156 2228 38208
rect 2280 38156 2286 38208
rect 2682 38156 2688 38208
rect 2740 38196 2746 38208
rect 4264 38196 4292 38295
rect 4430 38292 4436 38304
rect 4488 38332 4494 38344
rect 5534 38332 5540 38344
rect 4488 38304 5540 38332
rect 4488 38292 4494 38304
rect 5534 38292 5540 38304
rect 5592 38292 5598 38344
rect 9861 38335 9919 38341
rect 9861 38301 9873 38335
rect 9907 38332 9919 38335
rect 9950 38332 9956 38344
rect 9907 38304 9956 38332
rect 9907 38301 9919 38304
rect 9861 38295 9919 38301
rect 9950 38292 9956 38304
rect 10008 38292 10014 38344
rect 10042 38196 10048 38208
rect 2740 38168 4292 38196
rect 10003 38168 10048 38196
rect 2740 38156 2746 38168
rect 10042 38156 10048 38168
rect 10100 38156 10106 38208
rect 860 38100 980 38128
rect 952 37992 980 38100
rect 1104 38106 10856 38128
rect 1104 38054 4214 38106
rect 4266 38054 4278 38106
rect 4330 38054 4342 38106
rect 4394 38054 4406 38106
rect 4458 38054 4470 38106
rect 4522 38054 7478 38106
rect 7530 38054 7542 38106
rect 7594 38054 7606 38106
rect 7658 38054 7670 38106
rect 7722 38054 7734 38106
rect 7786 38054 10856 38106
rect 1104 38032 10856 38054
rect 1118 37992 1124 38004
rect 952 37964 1124 37992
rect 1118 37952 1124 37964
rect 1176 37952 1182 38004
rect 1670 37952 1676 38004
rect 1728 37992 1734 38004
rect 1949 37995 2007 38001
rect 1949 37992 1961 37995
rect 1728 37964 1961 37992
rect 1728 37952 1734 37964
rect 1949 37961 1961 37964
rect 1995 37961 2007 37995
rect 2774 37992 2780 38004
rect 2735 37964 2780 37992
rect 1949 37955 2007 37961
rect 2774 37952 2780 37964
rect 2832 37952 2838 38004
rect 9858 37952 9864 38004
rect 9916 37992 9922 38004
rect 9953 37995 10011 38001
rect 9953 37992 9965 37995
rect 9916 37964 9965 37992
rect 9916 37952 9922 37964
rect 9953 37961 9965 37964
rect 9999 37961 10011 37995
rect 9953 37955 10011 37961
rect 1210 37924 1216 37936
rect 768 37896 1216 37924
rect 1210 37884 1216 37896
rect 1268 37884 1274 37936
rect 2958 37924 2964 37936
rect 1688 37896 2964 37924
rect 1688 37865 1716 37896
rect 2958 37884 2964 37896
rect 3016 37884 3022 37936
rect 1673 37859 1731 37865
rect 1673 37825 1685 37859
rect 1719 37825 1731 37859
rect 1673 37819 1731 37825
rect 1765 37859 1823 37865
rect 1765 37825 1777 37859
rect 1811 37856 1823 37859
rect 2590 37856 2596 37868
rect 1811 37828 2596 37856
rect 1811 37825 1823 37828
rect 1765 37819 1823 37825
rect 1394 37748 1400 37800
rect 1452 37788 1458 37800
rect 1780 37788 1808 37819
rect 2590 37816 2596 37828
rect 2648 37816 2654 37868
rect 3237 37859 3295 37865
rect 3237 37825 3249 37859
rect 3283 37856 3295 37859
rect 3786 37856 3792 37868
rect 3283 37828 3792 37856
rect 3283 37825 3295 37828
rect 3237 37819 3295 37825
rect 3786 37816 3792 37828
rect 3844 37816 3850 37868
rect 3973 37859 4031 37865
rect 3973 37825 3985 37859
rect 4019 37856 4031 37859
rect 6730 37856 6736 37868
rect 4019 37828 6736 37856
rect 4019 37825 4031 37828
rect 3973 37819 4031 37825
rect 6730 37816 6736 37828
rect 6788 37816 6794 37868
rect 10137 37859 10195 37865
rect 10137 37825 10149 37859
rect 10183 37856 10195 37859
rect 10226 37856 10232 37868
rect 10183 37828 10232 37856
rect 10183 37825 10195 37828
rect 10137 37819 10195 37825
rect 10226 37816 10232 37828
rect 10284 37816 10290 37868
rect 1452 37760 1808 37788
rect 1452 37748 1458 37760
rect 1946 37748 1952 37800
rect 2004 37788 2010 37800
rect 2314 37788 2320 37800
rect 2004 37760 2320 37788
rect 2004 37748 2010 37760
rect 2314 37748 2320 37760
rect 2372 37748 2378 37800
rect 2409 37791 2467 37797
rect 2409 37757 2421 37791
rect 2455 37788 2467 37791
rect 2682 37788 2688 37800
rect 2455 37760 2688 37788
rect 2455 37757 2467 37760
rect 2409 37751 2467 37757
rect 1670 37680 1676 37732
rect 1728 37720 1734 37732
rect 2424 37720 2452 37751
rect 2682 37748 2688 37760
rect 2740 37748 2746 37800
rect 1728 37692 2452 37720
rect 1728 37680 1734 37692
rect 3510 37680 3516 37732
rect 3568 37720 3574 37732
rect 4157 37723 4215 37729
rect 4157 37720 4169 37723
rect 3568 37692 4169 37720
rect 3568 37680 3574 37692
rect 4157 37689 4169 37692
rect 4203 37689 4215 37723
rect 4157 37683 4215 37689
rect 14 37612 20 37664
rect 72 37652 78 37664
rect 1946 37652 1952 37664
rect 72 37624 1952 37652
rect 72 37612 78 37624
rect 1946 37612 1952 37624
rect 2004 37612 2010 37664
rect 3418 37652 3424 37664
rect 3379 37624 3424 37652
rect 3418 37612 3424 37624
rect 3476 37612 3482 37664
rect 1104 37562 10856 37584
rect 1104 37510 2582 37562
rect 2634 37510 2646 37562
rect 2698 37510 2710 37562
rect 2762 37510 2774 37562
rect 2826 37510 2838 37562
rect 2890 37510 5846 37562
rect 5898 37510 5910 37562
rect 5962 37510 5974 37562
rect 6026 37510 6038 37562
rect 6090 37510 6102 37562
rect 6154 37510 9110 37562
rect 9162 37510 9174 37562
rect 9226 37510 9238 37562
rect 9290 37510 9302 37562
rect 9354 37510 9366 37562
rect 9418 37510 10856 37562
rect 1104 37488 10856 37510
rect 1486 37408 1492 37460
rect 1544 37448 1550 37460
rect 2222 37448 2228 37460
rect 1544 37420 2228 37448
rect 1544 37408 1550 37420
rect 2222 37408 2228 37420
rect 2280 37408 2286 37460
rect 2498 37408 2504 37460
rect 2556 37448 2562 37460
rect 2777 37451 2835 37457
rect 2777 37448 2789 37451
rect 2556 37420 2789 37448
rect 2556 37408 2562 37420
rect 2777 37417 2789 37420
rect 2823 37417 2835 37451
rect 2777 37411 2835 37417
rect 566 37340 572 37392
rect 624 37380 630 37392
rect 624 37352 1808 37380
rect 624 37340 630 37352
rect 1670 37312 1676 37324
rect 1044 37284 1676 37312
rect 1044 36700 1072 37284
rect 1670 37272 1676 37284
rect 1728 37272 1734 37324
rect 1780 37312 1808 37352
rect 1854 37340 1860 37392
rect 1912 37380 1918 37392
rect 3973 37383 4031 37389
rect 3973 37380 3985 37383
rect 1912 37352 3985 37380
rect 1912 37340 1918 37352
rect 3973 37349 3985 37352
rect 4019 37349 4031 37383
rect 3973 37343 4031 37349
rect 1780 37284 2728 37312
rect 1397 37247 1455 37253
rect 1397 37213 1409 37247
rect 1443 37244 1455 37247
rect 1486 37244 1492 37256
rect 1443 37216 1492 37244
rect 1443 37213 1455 37216
rect 1397 37207 1455 37213
rect 1486 37204 1492 37216
rect 1544 37204 1550 37256
rect 2700 37188 2728 37284
rect 5626 37272 5632 37324
rect 5684 37312 5690 37324
rect 7098 37312 7104 37324
rect 5684 37284 7104 37312
rect 5684 37272 5690 37284
rect 7098 37272 7104 37284
rect 7156 37272 7162 37324
rect 3694 37204 3700 37256
rect 3752 37244 3758 37256
rect 3789 37247 3847 37253
rect 3789 37244 3801 37247
rect 3752 37216 3801 37244
rect 3752 37204 3758 37216
rect 3789 37213 3801 37216
rect 3835 37213 3847 37247
rect 9858 37244 9864 37256
rect 9819 37216 9864 37244
rect 3789 37207 3847 37213
rect 9858 37204 9864 37216
rect 9916 37204 9922 37256
rect 2222 37136 2228 37188
rect 2280 37176 2286 37188
rect 2314 37176 2320 37188
rect 2280 37148 2320 37176
rect 2280 37136 2286 37148
rect 2314 37136 2320 37148
rect 2372 37136 2378 37188
rect 2682 37176 2688 37188
rect 2643 37148 2688 37176
rect 2682 37136 2688 37148
rect 2740 37136 2746 37188
rect 1578 37108 1584 37120
rect 1539 37080 1584 37108
rect 1578 37068 1584 37080
rect 1636 37068 1642 37120
rect 2958 37068 2964 37120
rect 3016 37108 3022 37120
rect 3694 37108 3700 37120
rect 3016 37080 3700 37108
rect 3016 37068 3022 37080
rect 3694 37068 3700 37080
rect 3752 37068 3758 37120
rect 10042 37108 10048 37120
rect 10003 37080 10048 37108
rect 10042 37068 10048 37080
rect 10100 37068 10106 37120
rect 1104 37018 10856 37040
rect 1104 36966 4214 37018
rect 4266 36966 4278 37018
rect 4330 36966 4342 37018
rect 4394 36966 4406 37018
rect 4458 36966 4470 37018
rect 4522 36966 7478 37018
rect 7530 36966 7542 37018
rect 7594 36966 7606 37018
rect 7658 36966 7670 37018
rect 7722 36966 7734 37018
rect 7786 36966 10856 37018
rect 1104 36944 10856 36966
rect 1118 36864 1124 36916
rect 1176 36904 1182 36916
rect 1857 36907 1915 36913
rect 1857 36904 1869 36907
rect 1176 36876 1869 36904
rect 1176 36864 1182 36876
rect 1857 36873 1869 36876
rect 1903 36873 1915 36907
rect 1857 36867 1915 36873
rect 2314 36864 2320 36916
rect 2372 36904 2378 36916
rect 2682 36904 2688 36916
rect 2372 36876 2688 36904
rect 2372 36864 2378 36876
rect 2682 36864 2688 36876
rect 2740 36864 2746 36916
rect 2961 36907 3019 36913
rect 2961 36873 2973 36907
rect 3007 36873 3019 36907
rect 2961 36867 3019 36873
rect 4617 36907 4675 36913
rect 4617 36873 4629 36907
rect 4663 36904 4675 36907
rect 4982 36904 4988 36916
rect 4663 36876 4988 36904
rect 4663 36873 4675 36876
rect 4617 36867 4675 36873
rect 1765 36839 1823 36845
rect 1765 36805 1777 36839
rect 1811 36836 1823 36839
rect 2866 36836 2872 36848
rect 1811 36808 2872 36836
rect 1811 36805 1823 36808
rect 1765 36799 1823 36805
rect 2866 36796 2872 36808
rect 2924 36796 2930 36848
rect 2976 36836 3004 36867
rect 4982 36864 4988 36876
rect 5040 36864 5046 36916
rect 4522 36836 4528 36848
rect 2976 36808 4528 36836
rect 2409 36771 2467 36777
rect 2409 36737 2421 36771
rect 2455 36768 2467 36771
rect 2498 36768 2504 36780
rect 2455 36740 2504 36768
rect 2455 36737 2467 36740
rect 2409 36731 2467 36737
rect 2498 36728 2504 36740
rect 2556 36728 2562 36780
rect 3252 36777 3280 36808
rect 4522 36796 4528 36808
rect 4580 36796 4586 36848
rect 3237 36771 3295 36777
rect 3237 36737 3249 36771
rect 3283 36737 3295 36771
rect 3237 36731 3295 36737
rect 4433 36771 4491 36777
rect 4433 36737 4445 36771
rect 4479 36768 4491 36771
rect 5534 36768 5540 36780
rect 4479 36740 5540 36768
rect 4479 36737 4491 36740
rect 4433 36731 4491 36737
rect 5534 36728 5540 36740
rect 5592 36768 5598 36780
rect 5718 36768 5724 36780
rect 5592 36740 5724 36768
rect 5592 36728 5598 36740
rect 5718 36728 5724 36740
rect 5776 36728 5782 36780
rect 9861 36771 9919 36777
rect 9861 36737 9873 36771
rect 9907 36768 9919 36771
rect 10134 36768 10140 36780
rect 9907 36740 10140 36768
rect 9907 36737 9919 36740
rect 9861 36731 9919 36737
rect 10134 36728 10140 36740
rect 10192 36728 10198 36780
rect 1118 36700 1124 36712
rect 1044 36672 1124 36700
rect 1118 36660 1124 36672
rect 1176 36660 1182 36712
rect 1854 36660 1860 36712
rect 1912 36700 1918 36712
rect 2225 36703 2283 36709
rect 2225 36700 2237 36703
rect 1912 36672 2237 36700
rect 1912 36660 1918 36672
rect 2225 36669 2237 36672
rect 2271 36700 2283 36703
rect 4249 36703 4307 36709
rect 4249 36700 4261 36703
rect 2271 36672 4261 36700
rect 2271 36669 2283 36672
rect 2225 36663 2283 36669
rect 4249 36669 4261 36672
rect 4295 36669 4307 36703
rect 4249 36663 4307 36669
rect 3418 36632 3424 36644
rect 3379 36604 3424 36632
rect 3418 36592 3424 36604
rect 3476 36592 3482 36644
rect 2498 36524 2504 36576
rect 2556 36564 2562 36576
rect 2593 36567 2651 36573
rect 2593 36564 2605 36567
rect 2556 36536 2605 36564
rect 2556 36524 2562 36536
rect 2593 36533 2605 36536
rect 2639 36533 2651 36567
rect 2593 36527 2651 36533
rect 3050 36524 3056 36576
rect 3108 36564 3114 36576
rect 3326 36564 3332 36576
rect 3108 36536 3332 36564
rect 3108 36524 3114 36536
rect 3326 36524 3332 36536
rect 3384 36524 3390 36576
rect 10042 36564 10048 36576
rect 10003 36536 10048 36564
rect 10042 36524 10048 36536
rect 10100 36524 10106 36576
rect 1104 36474 10856 36496
rect 1104 36422 2582 36474
rect 2634 36422 2646 36474
rect 2698 36422 2710 36474
rect 2762 36422 2774 36474
rect 2826 36422 2838 36474
rect 2890 36422 5846 36474
rect 5898 36422 5910 36474
rect 5962 36422 5974 36474
rect 6026 36422 6038 36474
rect 6090 36422 6102 36474
rect 6154 36422 9110 36474
rect 9162 36422 9174 36474
rect 9226 36422 9238 36474
rect 9290 36422 9302 36474
rect 9354 36422 9366 36474
rect 9418 36422 10856 36474
rect 1104 36400 10856 36422
rect 2961 36363 3019 36369
rect 2961 36329 2973 36363
rect 3007 36360 3019 36363
rect 6822 36360 6828 36372
rect 3007 36332 6828 36360
rect 3007 36329 3019 36332
rect 2961 36323 3019 36329
rect 6822 36320 6828 36332
rect 6880 36320 6886 36372
rect 9217 36363 9275 36369
rect 9217 36329 9229 36363
rect 9263 36360 9275 36363
rect 9674 36360 9680 36372
rect 9263 36332 9680 36360
rect 9263 36329 9275 36332
rect 9217 36323 9275 36329
rect 9674 36320 9680 36332
rect 9732 36320 9738 36372
rect 750 36184 756 36236
rect 808 36224 814 36236
rect 1765 36227 1823 36233
rect 1765 36224 1777 36227
rect 808 36196 1777 36224
rect 808 36184 814 36196
rect 1765 36193 1777 36196
rect 1811 36193 1823 36227
rect 1765 36187 1823 36193
rect 1486 36156 1492 36168
rect 1447 36128 1492 36156
rect 1486 36116 1492 36128
rect 1544 36116 1550 36168
rect 2498 36116 2504 36168
rect 2556 36156 2562 36168
rect 2869 36159 2927 36165
rect 2869 36156 2881 36159
rect 2556 36128 2881 36156
rect 2556 36116 2562 36128
rect 2869 36125 2881 36128
rect 2915 36125 2927 36159
rect 2869 36119 2927 36125
rect 5534 36116 5540 36168
rect 5592 36156 5598 36168
rect 9401 36159 9459 36165
rect 9401 36156 9413 36159
rect 5592 36128 9413 36156
rect 5592 36116 5598 36128
rect 9401 36125 9413 36128
rect 9447 36125 9459 36159
rect 9401 36119 9459 36125
rect 9766 36116 9772 36168
rect 9824 36156 9830 36168
rect 9861 36159 9919 36165
rect 9861 36156 9873 36159
rect 9824 36128 9873 36156
rect 9824 36116 9830 36128
rect 9861 36125 9873 36128
rect 9907 36125 9919 36159
rect 9861 36119 9919 36125
rect 10042 36020 10048 36032
rect 10003 35992 10048 36020
rect 10042 35980 10048 35992
rect 10100 35980 10106 36032
rect 1104 35930 10856 35952
rect 1104 35878 4214 35930
rect 4266 35878 4278 35930
rect 4330 35878 4342 35930
rect 4394 35878 4406 35930
rect 4458 35878 4470 35930
rect 4522 35878 7478 35930
rect 7530 35878 7542 35930
rect 7594 35878 7606 35930
rect 7658 35878 7670 35930
rect 7722 35878 7734 35930
rect 7786 35878 10856 35930
rect 1104 35856 10856 35878
rect 4985 35819 5043 35825
rect 4985 35785 4997 35819
rect 5031 35816 5043 35819
rect 5534 35816 5540 35828
rect 5031 35788 5540 35816
rect 5031 35785 5043 35788
rect 4985 35779 5043 35785
rect 5534 35776 5540 35788
rect 5592 35776 5598 35828
rect 9950 35816 9956 35828
rect 9911 35788 9956 35816
rect 9950 35776 9956 35788
rect 10008 35776 10014 35828
rect 3510 35708 3516 35760
rect 3568 35748 3574 35760
rect 3697 35751 3755 35757
rect 3697 35748 3709 35751
rect 3568 35720 3709 35748
rect 3568 35708 3574 35720
rect 3697 35717 3709 35720
rect 3743 35717 3755 35751
rect 3697 35711 3755 35717
rect 4065 35751 4123 35757
rect 4065 35717 4077 35751
rect 4111 35748 4123 35751
rect 4430 35748 4436 35760
rect 4111 35720 4436 35748
rect 4111 35717 4123 35720
rect 4065 35711 4123 35717
rect 4430 35708 4436 35720
rect 4488 35748 4494 35760
rect 5718 35748 5724 35760
rect 4488 35720 5724 35748
rect 4488 35708 4494 35720
rect 474 35640 480 35692
rect 532 35680 538 35692
rect 1397 35683 1455 35689
rect 1397 35680 1409 35683
rect 532 35652 1409 35680
rect 532 35640 538 35652
rect 1397 35649 1409 35652
rect 1443 35649 1455 35683
rect 1397 35643 1455 35649
rect 2133 35683 2191 35689
rect 2133 35649 2145 35683
rect 2179 35680 2191 35683
rect 3786 35680 3792 35692
rect 2179 35652 3792 35680
rect 2179 35649 2191 35652
rect 2133 35643 2191 35649
rect 3786 35640 3792 35652
rect 3844 35640 3850 35692
rect 4816 35689 4844 35720
rect 5718 35708 5724 35720
rect 5776 35708 5782 35760
rect 4801 35683 4859 35689
rect 4801 35649 4813 35683
rect 4847 35649 4859 35683
rect 4801 35643 4859 35649
rect 4890 35640 4896 35692
rect 4948 35680 4954 35692
rect 10137 35683 10195 35689
rect 10137 35680 10149 35683
rect 4948 35652 10149 35680
rect 4948 35640 4954 35652
rect 10137 35649 10149 35652
rect 10183 35649 10195 35683
rect 10137 35643 10195 35649
rect 4614 35612 4620 35624
rect 4575 35584 4620 35612
rect 4614 35572 4620 35584
rect 4672 35572 4678 35624
rect 2314 35544 2320 35556
rect 2275 35516 2320 35544
rect 2314 35504 2320 35516
rect 2372 35504 2378 35556
rect 1578 35476 1584 35488
rect 1539 35448 1584 35476
rect 1578 35436 1584 35448
rect 1636 35436 1642 35488
rect 1104 35386 10856 35408
rect 1104 35334 2582 35386
rect 2634 35334 2646 35386
rect 2698 35334 2710 35386
rect 2762 35334 2774 35386
rect 2826 35334 2838 35386
rect 2890 35334 5846 35386
rect 5898 35334 5910 35386
rect 5962 35334 5974 35386
rect 6026 35334 6038 35386
rect 6090 35334 6102 35386
rect 6154 35334 9110 35386
rect 9162 35334 9174 35386
rect 9226 35334 9238 35386
rect 9290 35334 9302 35386
rect 9354 35334 9366 35386
rect 9418 35334 10856 35386
rect 1104 35312 10856 35334
rect 1486 35232 1492 35284
rect 1544 35272 1550 35284
rect 1949 35275 2007 35281
rect 1949 35272 1961 35275
rect 1544 35244 1961 35272
rect 1544 35232 1550 35244
rect 1949 35241 1961 35244
rect 1995 35241 2007 35275
rect 4890 35272 4896 35284
rect 4851 35244 4896 35272
rect 1949 35235 2007 35241
rect 4890 35232 4896 35244
rect 4948 35232 4954 35284
rect 4614 35204 4620 35216
rect 1596 35176 4620 35204
rect 1486 35028 1492 35080
rect 1544 35068 1550 35080
rect 1596 35077 1624 35176
rect 4614 35164 4620 35176
rect 4672 35164 4678 35216
rect 5166 35204 5172 35216
rect 5000 35176 5172 35204
rect 3970 35096 3976 35148
rect 4028 35136 4034 35148
rect 4430 35136 4436 35148
rect 4028 35108 4436 35136
rect 4028 35096 4034 35108
rect 4430 35096 4436 35108
rect 4488 35136 4494 35148
rect 4488 35108 4752 35136
rect 4488 35096 4494 35108
rect 1581 35071 1639 35077
rect 1581 35068 1593 35071
rect 1544 35040 1593 35068
rect 1544 35028 1550 35040
rect 1581 35037 1593 35040
rect 1627 35037 1639 35071
rect 1581 35031 1639 35037
rect 1765 35071 1823 35077
rect 1765 35037 1777 35071
rect 1811 35037 1823 35071
rect 2406 35068 2412 35080
rect 2367 35040 2412 35068
rect 1765 35031 1823 35037
rect 1394 34960 1400 35012
rect 1452 35000 1458 35012
rect 1780 35000 1808 35031
rect 2406 35028 2412 35040
rect 2464 35028 2470 35080
rect 3694 35028 3700 35080
rect 3752 35068 3758 35080
rect 4724 35077 4752 35108
rect 5000 35080 5028 35176
rect 5166 35164 5172 35176
rect 5224 35164 5230 35216
rect 4525 35071 4583 35077
rect 4525 35068 4537 35071
rect 3752 35040 4537 35068
rect 3752 35028 3758 35040
rect 4525 35037 4537 35040
rect 4571 35037 4583 35071
rect 4525 35031 4583 35037
rect 4709 35071 4767 35077
rect 4709 35037 4721 35071
rect 4755 35037 4767 35071
rect 4709 35031 4767 35037
rect 4982 35028 4988 35080
rect 5040 35028 5046 35080
rect 5166 35028 5172 35080
rect 5224 35068 5230 35080
rect 9861 35071 9919 35077
rect 9861 35068 9873 35071
rect 5224 35040 9873 35068
rect 5224 35028 5230 35040
rect 9861 35037 9873 35040
rect 9907 35037 9919 35071
rect 9861 35031 9919 35037
rect 2498 35000 2504 35012
rect 1452 34972 2504 35000
rect 1452 34960 1458 34972
rect 2498 34960 2504 34972
rect 2556 34960 2562 35012
rect 2593 34935 2651 34941
rect 2593 34901 2605 34935
rect 2639 34932 2651 34935
rect 2774 34932 2780 34944
rect 2639 34904 2780 34932
rect 2639 34901 2651 34904
rect 2593 34895 2651 34901
rect 2774 34892 2780 34904
rect 2832 34892 2838 34944
rect 10042 34932 10048 34944
rect 10003 34904 10048 34932
rect 10042 34892 10048 34904
rect 10100 34892 10106 34944
rect 1104 34842 10856 34864
rect 1104 34790 4214 34842
rect 4266 34790 4278 34842
rect 4330 34790 4342 34842
rect 4394 34790 4406 34842
rect 4458 34790 4470 34842
rect 4522 34790 7478 34842
rect 7530 34790 7542 34842
rect 7594 34790 7606 34842
rect 7658 34790 7670 34842
rect 7722 34790 7734 34842
rect 7786 34790 10856 34842
rect 1104 34768 10856 34790
rect 1578 34728 1584 34740
rect 1539 34700 1584 34728
rect 1578 34688 1584 34700
rect 1636 34688 1642 34740
rect 9582 34688 9588 34740
rect 9640 34728 9646 34740
rect 10045 34731 10103 34737
rect 10045 34728 10057 34731
rect 9640 34700 10057 34728
rect 9640 34688 9646 34700
rect 10045 34697 10057 34700
rect 10091 34697 10103 34731
rect 10045 34691 10103 34697
rect 3970 34620 3976 34672
rect 4028 34620 4034 34672
rect 4341 34663 4399 34669
rect 4341 34629 4353 34663
rect 4387 34660 4399 34663
rect 10226 34660 10232 34672
rect 4387 34632 10232 34660
rect 4387 34629 4399 34632
rect 4341 34623 4399 34629
rect 10226 34620 10232 34632
rect 10284 34620 10290 34672
rect 382 34552 388 34604
rect 440 34592 446 34604
rect 1397 34595 1455 34601
rect 1397 34592 1409 34595
rect 440 34564 1409 34592
rect 440 34552 446 34564
rect 1397 34561 1409 34564
rect 1443 34561 1455 34595
rect 1397 34555 1455 34561
rect 2038 34552 2044 34604
rect 2096 34592 2102 34604
rect 2133 34595 2191 34601
rect 2133 34592 2145 34595
rect 2096 34564 2145 34592
rect 2096 34552 2102 34564
rect 2133 34561 2145 34564
rect 2179 34561 2191 34595
rect 2133 34555 2191 34561
rect 2869 34595 2927 34601
rect 2869 34561 2881 34595
rect 2915 34592 2927 34595
rect 2958 34592 2964 34604
rect 2915 34564 2964 34592
rect 2915 34561 2927 34564
rect 2869 34555 2927 34561
rect 2958 34552 2964 34564
rect 3016 34552 3022 34604
rect 3988 34592 4016 34620
rect 4154 34592 4160 34604
rect 3988 34564 4160 34592
rect 4154 34552 4160 34564
rect 4212 34552 4218 34604
rect 9674 34552 9680 34604
rect 9732 34592 9738 34604
rect 9861 34595 9919 34601
rect 9861 34592 9873 34595
rect 9732 34564 9873 34592
rect 9732 34552 9738 34564
rect 9861 34561 9873 34564
rect 9907 34561 9919 34595
rect 9861 34555 9919 34561
rect 3970 34524 3976 34536
rect 3931 34496 3976 34524
rect 3970 34484 3976 34496
rect 4028 34484 4034 34536
rect 2038 34416 2044 34468
rect 2096 34456 2102 34468
rect 2222 34456 2228 34468
rect 2096 34428 2228 34456
rect 2096 34416 2102 34428
rect 2222 34416 2228 34428
rect 2280 34416 2286 34468
rect 1394 34348 1400 34400
rect 1452 34388 1458 34400
rect 2317 34391 2375 34397
rect 2317 34388 2329 34391
rect 1452 34360 2329 34388
rect 1452 34348 1458 34360
rect 2317 34357 2329 34360
rect 2363 34357 2375 34391
rect 3050 34388 3056 34400
rect 3011 34360 3056 34388
rect 2317 34351 2375 34357
rect 3050 34348 3056 34360
rect 3108 34348 3114 34400
rect 1104 34298 10856 34320
rect 1104 34246 2582 34298
rect 2634 34246 2646 34298
rect 2698 34246 2710 34298
rect 2762 34246 2774 34298
rect 2826 34246 2838 34298
rect 2890 34246 5846 34298
rect 5898 34246 5910 34298
rect 5962 34246 5974 34298
rect 6026 34246 6038 34298
rect 6090 34246 6102 34298
rect 6154 34246 9110 34298
rect 9162 34246 9174 34298
rect 9226 34246 9238 34298
rect 9290 34246 9302 34298
rect 9354 34246 9366 34298
rect 9418 34246 10856 34298
rect 1104 34224 10856 34246
rect 9858 34144 9864 34196
rect 9916 34184 9922 34196
rect 9953 34187 10011 34193
rect 9953 34184 9965 34187
rect 9916 34156 9965 34184
rect 9916 34144 9922 34156
rect 9953 34153 9965 34156
rect 9999 34153 10011 34187
rect 9953 34147 10011 34153
rect 198 34076 204 34128
rect 256 34116 262 34128
rect 2041 34119 2099 34125
rect 2041 34116 2053 34119
rect 256 34088 2053 34116
rect 256 34076 262 34088
rect 2041 34085 2053 34088
rect 2087 34085 2099 34119
rect 2041 34079 2099 34085
rect 3789 34119 3847 34125
rect 3789 34085 3801 34119
rect 3835 34116 3847 34119
rect 10134 34116 10140 34128
rect 3835 34088 10140 34116
rect 3835 34085 3847 34088
rect 3789 34079 3847 34085
rect 10134 34076 10140 34088
rect 10192 34076 10198 34128
rect 2406 33940 2412 33992
rect 2464 33980 2470 33992
rect 2685 33983 2743 33989
rect 2685 33980 2697 33983
rect 2464 33952 2697 33980
rect 2464 33940 2470 33952
rect 2685 33949 2697 33952
rect 2731 33949 2743 33983
rect 2685 33943 2743 33949
rect 2866 33940 2872 33992
rect 2924 33991 2930 33992
rect 2924 33985 2947 33991
rect 2935 33982 2947 33985
rect 3053 33983 3111 33989
rect 2935 33954 3015 33982
rect 2935 33951 2947 33954
rect 2924 33945 2947 33951
rect 2924 33940 2930 33945
rect 1857 33915 1915 33921
rect 1857 33881 1869 33915
rect 1903 33912 1915 33915
rect 2222 33912 2228 33924
rect 1903 33884 2228 33912
rect 1903 33881 1915 33884
rect 1857 33875 1915 33881
rect 2222 33872 2228 33884
rect 2280 33872 2286 33924
rect 2314 33872 2320 33924
rect 2372 33912 2378 33924
rect 2976 33912 3004 33954
rect 3053 33949 3065 33983
rect 3099 33980 3111 33983
rect 3973 33983 4031 33989
rect 3973 33980 3985 33983
rect 3099 33952 3985 33980
rect 3099 33949 3111 33952
rect 3053 33943 3111 33949
rect 3973 33949 3985 33952
rect 4019 33949 4031 33983
rect 10134 33980 10140 33992
rect 10095 33952 10140 33980
rect 3973 33943 4031 33949
rect 10134 33940 10140 33952
rect 10192 33940 10198 33992
rect 3786 33912 3792 33924
rect 2372 33884 2774 33912
rect 2976 33884 3792 33912
rect 2372 33872 2378 33884
rect 2746 33844 2774 33884
rect 3786 33872 3792 33884
rect 3844 33872 3850 33924
rect 3970 33844 3976 33856
rect 2746 33816 3976 33844
rect 3970 33804 3976 33816
rect 4028 33804 4034 33856
rect 1104 33754 10856 33776
rect 1104 33702 4214 33754
rect 4266 33702 4278 33754
rect 4330 33702 4342 33754
rect 4394 33702 4406 33754
rect 4458 33702 4470 33754
rect 4522 33702 7478 33754
rect 7530 33702 7542 33754
rect 7594 33702 7606 33754
rect 7658 33702 7670 33754
rect 7722 33702 7734 33754
rect 7786 33702 10856 33754
rect 1104 33680 10856 33702
rect 2222 33640 2228 33652
rect 2183 33612 2228 33640
rect 2222 33600 2228 33612
rect 2280 33600 2286 33652
rect 2869 33643 2927 33649
rect 2869 33609 2881 33643
rect 2915 33640 2927 33643
rect 3234 33640 3240 33652
rect 2915 33612 3240 33640
rect 2915 33609 2927 33612
rect 2869 33603 2927 33609
rect 3234 33600 3240 33612
rect 3292 33600 3298 33652
rect 4525 33643 4583 33649
rect 4525 33609 4537 33643
rect 4571 33640 4583 33643
rect 10134 33640 10140 33652
rect 4571 33612 10140 33640
rect 4571 33609 4583 33612
rect 4525 33603 4583 33609
rect 10134 33600 10140 33612
rect 10192 33600 10198 33652
rect 2314 33572 2320 33584
rect 1964 33544 2320 33572
rect 1964 33513 1992 33544
rect 2314 33532 2320 33544
rect 2372 33532 2378 33584
rect 2498 33532 2504 33584
rect 2556 33532 2562 33584
rect 1949 33507 2007 33513
rect 1949 33473 1961 33507
rect 1995 33473 2007 33507
rect 1949 33467 2007 33473
rect 2041 33507 2099 33513
rect 2041 33473 2053 33507
rect 2087 33504 2099 33507
rect 2222 33504 2228 33516
rect 2087 33476 2228 33504
rect 2087 33473 2099 33476
rect 2041 33467 2099 33473
rect 2222 33464 2228 33476
rect 2280 33504 2286 33516
rect 2516 33504 2544 33532
rect 2280 33476 2544 33504
rect 2777 33507 2835 33513
rect 2280 33464 2286 33476
rect 2777 33473 2789 33507
rect 2823 33504 2835 33507
rect 2958 33504 2964 33516
rect 2823 33476 2964 33504
rect 2823 33473 2835 33476
rect 2777 33467 2835 33473
rect 2958 33464 2964 33476
rect 3016 33464 3022 33516
rect 3050 33464 3056 33516
rect 3108 33504 3114 33516
rect 3234 33504 3240 33516
rect 3108 33476 3240 33504
rect 3108 33464 3114 33476
rect 3234 33464 3240 33476
rect 3292 33464 3298 33516
rect 3786 33464 3792 33516
rect 3844 33504 3850 33516
rect 4341 33507 4399 33513
rect 4341 33504 4353 33507
rect 3844 33476 4353 33504
rect 3844 33464 3850 33476
rect 4341 33473 4353 33476
rect 4387 33473 4399 33507
rect 4341 33467 4399 33473
rect 5534 33464 5540 33516
rect 5592 33504 5598 33516
rect 9861 33507 9919 33513
rect 9861 33504 9873 33507
rect 5592 33476 9873 33504
rect 5592 33464 5598 33476
rect 9861 33473 9873 33476
rect 9907 33473 9919 33507
rect 9861 33467 9919 33473
rect 2498 33396 2504 33448
rect 2556 33436 2562 33448
rect 4157 33439 4215 33445
rect 4157 33436 4169 33439
rect 2556 33408 4169 33436
rect 2556 33396 2562 33408
rect 4157 33405 4169 33408
rect 4203 33405 4215 33439
rect 4157 33399 4215 33405
rect 2866 33328 2872 33380
rect 2924 33368 2930 33380
rect 3050 33368 3056 33380
rect 2924 33340 3056 33368
rect 2924 33328 2930 33340
rect 3050 33328 3056 33340
rect 3108 33328 3114 33380
rect 10042 33368 10048 33380
rect 10003 33340 10048 33368
rect 10042 33328 10048 33340
rect 10100 33328 10106 33380
rect 1104 33210 10856 33232
rect 1104 33158 2582 33210
rect 2634 33158 2646 33210
rect 2698 33158 2710 33210
rect 2762 33158 2774 33210
rect 2826 33158 2838 33210
rect 2890 33158 5846 33210
rect 5898 33158 5910 33210
rect 5962 33158 5974 33210
rect 6026 33158 6038 33210
rect 6090 33158 6102 33210
rect 6154 33158 9110 33210
rect 9162 33158 9174 33210
rect 9226 33158 9238 33210
rect 9290 33158 9302 33210
rect 9354 33158 9366 33210
rect 9418 33158 10856 33210
rect 1104 33136 10856 33158
rect 3789 33099 3847 33105
rect 3789 33065 3801 33099
rect 3835 33096 3847 33099
rect 9674 33096 9680 33108
rect 3835 33068 9680 33096
rect 3835 33065 3847 33068
rect 3789 33059 3847 33065
rect 9674 33056 9680 33068
rect 9732 33056 9738 33108
rect 1486 32920 1492 32972
rect 1544 32960 1550 32972
rect 1544 32932 2268 32960
rect 1544 32920 1550 32932
rect 1397 32895 1455 32901
rect 1397 32861 1409 32895
rect 1443 32892 1455 32895
rect 1670 32892 1676 32904
rect 1443 32864 1676 32892
rect 1443 32861 1455 32864
rect 1397 32855 1455 32861
rect 1670 32852 1676 32864
rect 1728 32852 1734 32904
rect 2130 32892 2136 32904
rect 2091 32864 2136 32892
rect 2130 32852 2136 32864
rect 2188 32852 2194 32904
rect 2240 32892 2268 32932
rect 2869 32895 2927 32901
rect 2869 32892 2881 32895
rect 2240 32864 2881 32892
rect 2869 32861 2881 32864
rect 2915 32861 2927 32895
rect 2869 32855 2927 32861
rect 3786 32852 3792 32904
rect 3844 32892 3850 32904
rect 3973 32895 4031 32901
rect 3973 32892 3985 32895
rect 3844 32864 3985 32892
rect 3844 32852 3850 32864
rect 3973 32861 3985 32864
rect 4019 32861 4031 32895
rect 9858 32892 9864 32904
rect 9819 32864 9864 32892
rect 3973 32855 4031 32861
rect 9858 32852 9864 32864
rect 9916 32852 9922 32904
rect 1581 32759 1639 32765
rect 1581 32756 1593 32759
rect 1044 32728 1593 32756
rect 1044 32552 1072 32728
rect 1581 32725 1593 32728
rect 1627 32725 1639 32759
rect 2314 32756 2320 32768
rect 2275 32728 2320 32756
rect 1581 32719 1639 32725
rect 2314 32716 2320 32728
rect 2372 32716 2378 32768
rect 2774 32716 2780 32768
rect 2832 32756 2838 32768
rect 3053 32759 3111 32765
rect 3053 32756 3065 32759
rect 2832 32728 3065 32756
rect 2832 32716 2838 32728
rect 3053 32725 3065 32728
rect 3099 32725 3111 32759
rect 3053 32719 3111 32725
rect 4982 32716 4988 32768
rect 5040 32756 5046 32768
rect 5718 32756 5724 32768
rect 5040 32728 5724 32756
rect 5040 32716 5046 32728
rect 5718 32716 5724 32728
rect 5776 32716 5782 32768
rect 10042 32756 10048 32768
rect 10003 32728 10048 32756
rect 10042 32716 10048 32728
rect 10100 32716 10106 32768
rect 1104 32666 10856 32688
rect 1104 32614 4214 32666
rect 4266 32614 4278 32666
rect 4330 32614 4342 32666
rect 4394 32614 4406 32666
rect 4458 32614 4470 32666
rect 4522 32614 7478 32666
rect 7530 32614 7542 32666
rect 7594 32614 7606 32666
rect 7658 32614 7670 32666
rect 7722 32614 7734 32666
rect 7786 32614 10856 32666
rect 1104 32592 10856 32614
rect 1578 32552 1584 32564
rect 1044 32524 1584 32552
rect 1578 32512 1584 32524
rect 1636 32512 1642 32564
rect 2409 32555 2467 32561
rect 2409 32521 2421 32555
rect 2455 32552 2467 32555
rect 2958 32552 2964 32564
rect 2455 32524 2964 32552
rect 2455 32521 2467 32524
rect 2409 32515 2467 32521
rect 2958 32512 2964 32524
rect 3016 32512 3022 32564
rect 3605 32555 3663 32561
rect 3605 32521 3617 32555
rect 3651 32552 3663 32555
rect 9858 32552 9864 32564
rect 3651 32524 9864 32552
rect 3651 32521 3663 32524
rect 3605 32515 3663 32521
rect 9858 32512 9864 32524
rect 9916 32512 9922 32564
rect 3878 32484 3884 32496
rect 2884 32456 3884 32484
rect 2222 32416 2228 32428
rect 2183 32388 2228 32416
rect 2222 32376 2228 32388
rect 2280 32376 2286 32428
rect 2884 32425 2912 32456
rect 3878 32444 3884 32456
rect 3936 32444 3942 32496
rect 2869 32419 2927 32425
rect 2869 32385 2881 32419
rect 2915 32385 2927 32419
rect 2869 32379 2927 32385
rect 3789 32419 3847 32425
rect 3789 32385 3801 32419
rect 3835 32385 3847 32419
rect 3789 32379 3847 32385
rect 4433 32419 4491 32425
rect 4433 32385 4445 32419
rect 4479 32416 4491 32419
rect 4982 32416 4988 32428
rect 4479 32388 4988 32416
rect 4479 32385 4491 32388
rect 4433 32379 4491 32385
rect 934 32308 940 32360
rect 992 32348 998 32360
rect 2041 32351 2099 32357
rect 2041 32348 2053 32351
rect 992 32320 2053 32348
rect 992 32308 998 32320
rect 2041 32317 2053 32320
rect 2087 32348 2099 32351
rect 3694 32348 3700 32360
rect 2087 32320 3700 32348
rect 2087 32317 2099 32320
rect 2041 32311 2099 32317
rect 3694 32308 3700 32320
rect 3752 32308 3758 32360
rect 3050 32280 3056 32292
rect 3011 32252 3056 32280
rect 3050 32240 3056 32252
rect 3108 32240 3114 32292
rect 3418 32172 3424 32224
rect 3476 32212 3482 32224
rect 3694 32212 3700 32224
rect 3476 32184 3700 32212
rect 3476 32172 3482 32184
rect 3694 32172 3700 32184
rect 3752 32172 3758 32224
rect 3804 32212 3832 32379
rect 4982 32376 4988 32388
rect 5040 32376 5046 32428
rect 4249 32283 4307 32289
rect 4249 32249 4261 32283
rect 4295 32280 4307 32283
rect 5166 32280 5172 32292
rect 4295 32252 5172 32280
rect 4295 32249 4307 32252
rect 4249 32243 4307 32249
rect 5166 32240 5172 32252
rect 5224 32240 5230 32292
rect 4706 32212 4712 32224
rect 3804 32184 4712 32212
rect 4706 32172 4712 32184
rect 4764 32172 4770 32224
rect 1104 32122 10856 32144
rect 1104 32070 2582 32122
rect 2634 32070 2646 32122
rect 2698 32070 2710 32122
rect 2762 32070 2774 32122
rect 2826 32070 2838 32122
rect 2890 32070 5846 32122
rect 5898 32070 5910 32122
rect 5962 32070 5974 32122
rect 6026 32070 6038 32122
rect 6090 32070 6102 32122
rect 6154 32070 9110 32122
rect 9162 32070 9174 32122
rect 9226 32070 9238 32122
rect 9290 32070 9302 32122
rect 9354 32070 9366 32122
rect 9418 32070 10856 32122
rect 1104 32048 10856 32070
rect 842 31968 848 32020
rect 900 32008 906 32020
rect 1949 32011 2007 32017
rect 1949 32008 1961 32011
rect 900 31980 1961 32008
rect 900 31968 906 31980
rect 1949 31977 1961 31980
rect 1995 31977 2007 32011
rect 1949 31971 2007 31977
rect 2498 31968 2504 32020
rect 2556 32008 2562 32020
rect 4246 32008 4252 32020
rect 2556 31980 2636 32008
rect 2556 31968 2562 31980
rect 2608 31952 2636 31980
rect 2792 31980 4252 32008
rect 1854 31900 1860 31952
rect 1912 31940 1918 31952
rect 1912 31912 2544 31940
rect 1912 31900 1918 31912
rect 2516 31884 2544 31912
rect 2590 31900 2596 31952
rect 2648 31900 2654 31952
rect 2792 31949 2820 31980
rect 4246 31968 4252 31980
rect 4304 31968 4310 32020
rect 4525 32011 4583 32017
rect 4525 31977 4537 32011
rect 4571 32008 4583 32011
rect 9766 32008 9772 32020
rect 4571 31980 9772 32008
rect 4571 31977 4583 31980
rect 4525 31971 4583 31977
rect 9766 31968 9772 31980
rect 9824 31968 9830 32020
rect 2777 31943 2835 31949
rect 2777 31909 2789 31943
rect 2823 31909 2835 31943
rect 3970 31940 3976 31952
rect 3931 31912 3976 31940
rect 2777 31903 2835 31909
rect 3970 31900 3976 31912
rect 4028 31900 4034 31952
rect 10042 31940 10048 31952
rect 10003 31912 10048 31940
rect 10042 31900 10048 31912
rect 10100 31900 10106 31952
rect 658 31832 664 31884
rect 716 31872 722 31884
rect 716 31844 2176 31872
rect 716 31832 722 31844
rect 2148 31816 2176 31844
rect 2222 31832 2228 31884
rect 2280 31832 2286 31884
rect 2498 31832 2504 31884
rect 2556 31832 2562 31884
rect 4614 31832 4620 31884
rect 4672 31872 4678 31884
rect 4672 31844 4844 31872
rect 4672 31832 4678 31844
rect 1118 31764 1124 31816
rect 1176 31804 1182 31816
rect 1394 31804 1400 31816
rect 1176 31776 1400 31804
rect 1176 31764 1182 31776
rect 1394 31764 1400 31776
rect 1452 31764 1458 31816
rect 2130 31764 2136 31816
rect 2188 31764 2194 31816
rect 2240 31804 2268 31832
rect 3789 31807 3847 31813
rect 3789 31804 3801 31807
rect 2240 31776 3801 31804
rect 3789 31773 3801 31776
rect 3835 31773 3847 31807
rect 3789 31767 3847 31773
rect 4709 31807 4767 31813
rect 4709 31773 4721 31807
rect 4755 31773 4767 31807
rect 4816 31804 4844 31844
rect 5350 31832 5356 31884
rect 5408 31872 5414 31884
rect 5626 31872 5632 31884
rect 5408 31844 5632 31872
rect 5408 31832 5414 31844
rect 5626 31832 5632 31844
rect 5684 31832 5690 31884
rect 9861 31807 9919 31813
rect 9861 31804 9873 31807
rect 4816 31776 9873 31804
rect 4709 31767 4767 31773
rect 9861 31773 9873 31776
rect 9907 31773 9919 31807
rect 9861 31767 9919 31773
rect 1578 31696 1584 31748
rect 1636 31696 1642 31748
rect 1854 31736 1860 31748
rect 1815 31708 1860 31736
rect 1854 31696 1860 31708
rect 1912 31696 1918 31748
rect 2222 31696 2228 31748
rect 2280 31736 2286 31748
rect 2593 31739 2651 31745
rect 2593 31736 2605 31739
rect 2280 31708 2605 31736
rect 2280 31696 2286 31708
rect 2593 31705 2605 31708
rect 2639 31705 2651 31739
rect 2593 31699 2651 31705
rect 3050 31696 3056 31748
rect 3108 31736 3114 31748
rect 4724 31736 4752 31767
rect 3108 31708 4752 31736
rect 3108 31696 3114 31708
rect 1118 31628 1124 31680
rect 1176 31668 1182 31680
rect 1596 31668 1624 31696
rect 1176 31640 1624 31668
rect 1176 31628 1182 31640
rect 2314 31628 2320 31680
rect 2372 31668 2378 31680
rect 2682 31668 2688 31680
rect 2372 31640 2688 31668
rect 2372 31628 2378 31640
rect 2682 31628 2688 31640
rect 2740 31628 2746 31680
rect 1104 31578 10856 31600
rect 1104 31526 4214 31578
rect 4266 31526 4278 31578
rect 4330 31526 4342 31578
rect 4394 31526 4406 31578
rect 4458 31526 4470 31578
rect 4522 31526 7478 31578
rect 7530 31526 7542 31578
rect 7594 31526 7606 31578
rect 7658 31526 7670 31578
rect 7722 31526 7734 31578
rect 7786 31526 10856 31578
rect 1104 31504 10856 31526
rect 1854 31424 1860 31476
rect 1912 31464 1918 31476
rect 1949 31467 2007 31473
rect 1949 31464 1961 31467
rect 1912 31436 1961 31464
rect 1912 31424 1918 31436
rect 1949 31433 1961 31436
rect 1995 31433 2007 31467
rect 1949 31427 2007 31433
rect 2314 31424 2320 31476
rect 2372 31464 2378 31476
rect 2498 31464 2504 31476
rect 2372 31436 2504 31464
rect 2372 31424 2378 31436
rect 2498 31424 2504 31436
rect 2556 31424 2562 31476
rect 3050 31424 3056 31476
rect 3108 31464 3114 31476
rect 3881 31467 3939 31473
rect 3881 31464 3893 31467
rect 3108 31436 3893 31464
rect 3108 31424 3114 31436
rect 3881 31433 3893 31436
rect 3927 31433 3939 31467
rect 3881 31427 3939 31433
rect 2682 31356 2688 31408
rect 2740 31356 2746 31408
rect 658 31288 664 31340
rect 716 31328 722 31340
rect 1765 31331 1823 31337
rect 1765 31328 1777 31331
rect 716 31300 1777 31328
rect 716 31288 722 31300
rect 1765 31297 1777 31300
rect 1811 31328 1823 31331
rect 2700 31328 2728 31356
rect 1811 31300 2728 31328
rect 2869 31331 2927 31337
rect 1811 31297 1823 31300
rect 1765 31291 1823 31297
rect 2869 31297 2881 31331
rect 2915 31328 2927 31331
rect 2958 31328 2964 31340
rect 2915 31300 2964 31328
rect 2915 31297 2927 31300
rect 2869 31291 2927 31297
rect 2958 31288 2964 31300
rect 3016 31328 3022 31340
rect 3697 31331 3755 31337
rect 3697 31328 3709 31331
rect 3016 31300 3709 31328
rect 3016 31288 3022 31300
rect 3697 31297 3709 31300
rect 3743 31297 3755 31331
rect 3697 31291 3755 31297
rect 5350 31288 5356 31340
rect 5408 31328 5414 31340
rect 5626 31328 5632 31340
rect 5408 31300 5632 31328
rect 5408 31288 5414 31300
rect 5626 31288 5632 31300
rect 5684 31288 5690 31340
rect 9858 31328 9864 31340
rect 9819 31300 9864 31328
rect 9858 31288 9864 31300
rect 9916 31288 9922 31340
rect 842 31220 848 31272
rect 900 31260 906 31272
rect 1581 31263 1639 31269
rect 1581 31260 1593 31263
rect 900 31232 1593 31260
rect 900 31220 906 31232
rect 1581 31229 1593 31232
rect 1627 31260 1639 31263
rect 2685 31263 2743 31269
rect 2685 31260 2697 31263
rect 1627 31232 2697 31260
rect 1627 31229 1639 31232
rect 1581 31223 1639 31229
rect 2685 31229 2697 31232
rect 2731 31229 2743 31263
rect 2685 31223 2743 31229
rect 3513 31263 3571 31269
rect 3513 31229 3525 31263
rect 3559 31260 3571 31263
rect 3878 31260 3884 31272
rect 3559 31232 3884 31260
rect 3559 31229 3571 31232
rect 3513 31223 3571 31229
rect 3878 31220 3884 31232
rect 3936 31220 3942 31272
rect 2406 31152 2412 31204
rect 2464 31192 2470 31204
rect 2590 31192 2596 31204
rect 2464 31164 2596 31192
rect 2464 31152 2470 31164
rect 2590 31152 2596 31164
rect 2648 31152 2654 31204
rect 3053 31195 3111 31201
rect 3053 31161 3065 31195
rect 3099 31192 3111 31195
rect 4890 31192 4896 31204
rect 3099 31164 4896 31192
rect 3099 31161 3111 31164
rect 3053 31155 3111 31161
rect 4890 31152 4896 31164
rect 4948 31152 4954 31204
rect 10042 31124 10048 31136
rect 10003 31096 10048 31124
rect 10042 31084 10048 31096
rect 10100 31084 10106 31136
rect 1104 31034 10856 31056
rect 1104 30982 2582 31034
rect 2634 30982 2646 31034
rect 2698 30982 2710 31034
rect 2762 30982 2774 31034
rect 2826 30982 2838 31034
rect 2890 30982 5846 31034
rect 5898 30982 5910 31034
rect 5962 30982 5974 31034
rect 6026 30982 6038 31034
rect 6090 30982 6102 31034
rect 6154 30982 9110 31034
rect 9162 30982 9174 31034
rect 9226 30982 9238 31034
rect 9290 30982 9302 31034
rect 9354 30982 9366 31034
rect 9418 30982 10856 31034
rect 1104 30960 10856 30982
rect 1949 30923 2007 30929
rect 1949 30889 1961 30923
rect 1995 30920 2007 30923
rect 3326 30920 3332 30932
rect 1995 30892 3332 30920
rect 1995 30889 2007 30892
rect 1949 30883 2007 30889
rect 3326 30880 3332 30892
rect 3384 30880 3390 30932
rect 4706 30812 4712 30864
rect 4764 30852 4770 30864
rect 4890 30852 4896 30864
rect 4764 30824 4896 30852
rect 4764 30812 4770 30824
rect 4890 30812 4896 30824
rect 4948 30812 4954 30864
rect 1762 30676 1768 30728
rect 1820 30716 1826 30728
rect 2501 30719 2559 30725
rect 2501 30716 2513 30719
rect 1820 30688 2513 30716
rect 1820 30676 1826 30688
rect 2501 30685 2513 30688
rect 2547 30685 2559 30719
rect 2501 30679 2559 30685
rect 4522 30676 4528 30728
rect 4580 30716 4586 30728
rect 4706 30716 4712 30728
rect 4580 30688 4712 30716
rect 4580 30676 4586 30688
rect 4706 30676 4712 30688
rect 4764 30676 4770 30728
rect 8294 30676 8300 30728
rect 8352 30716 8358 30728
rect 9861 30719 9919 30725
rect 9861 30716 9873 30719
rect 8352 30688 9873 30716
rect 8352 30676 8358 30688
rect 9861 30685 9873 30688
rect 9907 30685 9919 30719
rect 9861 30679 9919 30685
rect 1854 30648 1860 30660
rect 1815 30620 1860 30648
rect 1854 30608 1860 30620
rect 1912 30608 1918 30660
rect 2685 30583 2743 30589
rect 2685 30549 2697 30583
rect 2731 30580 2743 30583
rect 2774 30580 2780 30592
rect 2731 30552 2780 30580
rect 2731 30549 2743 30552
rect 2685 30543 2743 30549
rect 2774 30540 2780 30552
rect 2832 30540 2838 30592
rect 10042 30580 10048 30592
rect 10003 30552 10048 30580
rect 10042 30540 10048 30552
rect 10100 30540 10106 30592
rect 1104 30490 10856 30512
rect 1104 30438 4214 30490
rect 4266 30438 4278 30490
rect 4330 30438 4342 30490
rect 4394 30438 4406 30490
rect 4458 30438 4470 30490
rect 4522 30438 7478 30490
rect 7530 30438 7542 30490
rect 7594 30438 7606 30490
rect 7658 30438 7670 30490
rect 7722 30438 7734 30490
rect 7786 30438 10856 30490
rect 1104 30416 10856 30438
rect 3786 30336 3792 30388
rect 3844 30336 3850 30388
rect 1118 30268 1124 30320
rect 1176 30308 1182 30320
rect 1857 30311 1915 30317
rect 1857 30308 1869 30311
rect 1176 30280 1869 30308
rect 1176 30268 1182 30280
rect 1857 30277 1869 30280
rect 1903 30277 1915 30311
rect 1857 30271 1915 30277
rect 2038 30268 2044 30320
rect 2096 30308 2102 30320
rect 2685 30311 2743 30317
rect 2096 30280 2636 30308
rect 2096 30268 2102 30280
rect 1670 30240 1676 30252
rect 1631 30212 1676 30240
rect 1670 30200 1676 30212
rect 1728 30200 1734 30252
rect 2501 30243 2559 30249
rect 2501 30209 2513 30243
rect 2547 30209 2559 30243
rect 2608 30240 2636 30280
rect 2685 30277 2697 30311
rect 2731 30308 2743 30311
rect 3804 30308 3832 30336
rect 2731 30280 3832 30308
rect 2731 30277 2743 30280
rect 2685 30271 2743 30277
rect 4522 30268 4528 30320
rect 4580 30308 4586 30320
rect 5718 30308 5724 30320
rect 4580 30280 5724 30308
rect 4580 30268 4586 30280
rect 5718 30268 5724 30280
rect 5776 30268 5782 30320
rect 3145 30243 3203 30249
rect 3145 30240 3157 30243
rect 2608 30212 3157 30240
rect 2501 30203 2559 30209
rect 3145 30209 3157 30212
rect 3191 30209 3203 30243
rect 3145 30203 3203 30209
rect 2314 30172 2320 30184
rect 2275 30144 2320 30172
rect 2314 30132 2320 30144
rect 2372 30132 2378 30184
rect 2516 30172 2544 30203
rect 3786 30200 3792 30252
rect 3844 30240 3850 30252
rect 4065 30243 4123 30249
rect 4065 30240 4077 30243
rect 3844 30212 4077 30240
rect 3844 30200 3850 30212
rect 4065 30209 4077 30212
rect 4111 30209 4123 30243
rect 4065 30203 4123 30209
rect 4709 30243 4767 30249
rect 4709 30209 4721 30243
rect 4755 30240 4767 30243
rect 5626 30240 5632 30252
rect 4755 30212 5632 30240
rect 4755 30209 4767 30212
rect 4709 30203 4767 30209
rect 5626 30200 5632 30212
rect 5684 30200 5690 30252
rect 2958 30172 2964 30184
rect 2516 30144 2964 30172
rect 2958 30132 2964 30144
rect 3016 30132 3022 30184
rect 3326 30104 3332 30116
rect 3287 30076 3332 30104
rect 3326 30064 3332 30076
rect 3384 30064 3390 30116
rect 4525 30107 4583 30113
rect 4525 30073 4537 30107
rect 4571 30104 4583 30107
rect 4614 30104 4620 30116
rect 4571 30076 4620 30104
rect 4571 30073 4583 30076
rect 4525 30067 4583 30073
rect 4614 30064 4620 30076
rect 4672 30064 4678 30116
rect 842 29996 848 30048
rect 900 30036 906 30048
rect 1854 30036 1860 30048
rect 900 30008 1860 30036
rect 900 29996 906 30008
rect 1854 29996 1860 30008
rect 1912 29996 1918 30048
rect 3881 30039 3939 30045
rect 3881 30005 3893 30039
rect 3927 30036 3939 30039
rect 9858 30036 9864 30048
rect 3927 30008 9864 30036
rect 3927 30005 3939 30008
rect 3881 29999 3939 30005
rect 9858 29996 9864 30008
rect 9916 29996 9922 30048
rect 1104 29946 10856 29968
rect 1104 29894 2582 29946
rect 2634 29894 2646 29946
rect 2698 29894 2710 29946
rect 2762 29894 2774 29946
rect 2826 29894 2838 29946
rect 2890 29894 5846 29946
rect 5898 29894 5910 29946
rect 5962 29894 5974 29946
rect 6026 29894 6038 29946
rect 6090 29894 6102 29946
rect 6154 29894 9110 29946
rect 9162 29894 9174 29946
rect 9226 29894 9238 29946
rect 9290 29894 9302 29946
rect 9354 29894 9366 29946
rect 9418 29894 10856 29946
rect 1104 29872 10856 29894
rect 750 29792 756 29844
rect 808 29832 814 29844
rect 2685 29835 2743 29841
rect 2685 29832 2697 29835
rect 808 29804 2697 29832
rect 808 29792 814 29804
rect 2685 29801 2697 29804
rect 2731 29801 2743 29835
rect 2685 29795 2743 29801
rect 7653 29835 7711 29841
rect 7653 29801 7665 29835
rect 7699 29832 7711 29835
rect 8294 29832 8300 29844
rect 7699 29804 8300 29832
rect 7699 29801 7711 29804
rect 7653 29795 7711 29801
rect 8294 29792 8300 29804
rect 8352 29792 8358 29844
rect 2041 29631 2099 29637
rect 2041 29597 2053 29631
rect 2087 29628 2099 29631
rect 6914 29628 6920 29640
rect 2087 29600 6920 29628
rect 2087 29597 2099 29600
rect 2041 29591 2099 29597
rect 6914 29588 6920 29600
rect 6972 29588 6978 29640
rect 7834 29628 7840 29640
rect 7795 29600 7840 29628
rect 7834 29588 7840 29600
rect 7892 29588 7898 29640
rect 10134 29628 10140 29640
rect 10095 29600 10140 29628
rect 10134 29588 10140 29600
rect 10192 29588 10198 29640
rect 1857 29563 1915 29569
rect 1857 29529 1869 29563
rect 1903 29529 1915 29563
rect 1857 29523 1915 29529
rect 2593 29563 2651 29569
rect 2593 29529 2605 29563
rect 2639 29560 2651 29563
rect 2774 29560 2780 29572
rect 2639 29532 2780 29560
rect 2639 29529 2651 29532
rect 2593 29523 2651 29529
rect 1872 29492 1900 29523
rect 2774 29520 2780 29532
rect 2832 29520 2838 29572
rect 3050 29492 3056 29504
rect 1872 29464 3056 29492
rect 3050 29452 3056 29464
rect 3108 29452 3114 29504
rect 1104 29402 10856 29424
rect 1104 29350 4214 29402
rect 4266 29350 4278 29402
rect 4330 29350 4342 29402
rect 4394 29350 4406 29402
rect 4458 29350 4470 29402
rect 4522 29350 7478 29402
rect 7530 29350 7542 29402
rect 7594 29350 7606 29402
rect 7658 29350 7670 29402
rect 7722 29350 7734 29402
rect 7786 29350 10856 29402
rect 1104 29328 10856 29350
rect 106 29248 112 29300
rect 164 29288 170 29300
rect 2133 29291 2191 29297
rect 2133 29288 2145 29291
rect 164 29260 2145 29288
rect 164 29248 170 29260
rect 2133 29257 2145 29260
rect 2179 29257 2191 29291
rect 2133 29251 2191 29257
rect 2869 29291 2927 29297
rect 2869 29257 2881 29291
rect 2915 29288 2927 29291
rect 3142 29288 3148 29300
rect 2915 29260 3148 29288
rect 2915 29257 2927 29260
rect 2869 29251 2927 29257
rect 3142 29248 3148 29260
rect 3200 29248 3206 29300
rect 2041 29223 2099 29229
rect 2041 29189 2053 29223
rect 2087 29220 2099 29223
rect 2087 29192 3188 29220
rect 2087 29189 2099 29192
rect 2041 29183 2099 29189
rect 3160 29164 3188 29192
rect 2777 29155 2835 29161
rect 2777 29121 2789 29155
rect 2823 29152 2835 29155
rect 2958 29152 2964 29164
rect 2823 29124 2964 29152
rect 2823 29121 2835 29124
rect 2777 29115 2835 29121
rect 2958 29112 2964 29124
rect 3016 29112 3022 29164
rect 3142 29112 3148 29164
rect 3200 29112 3206 29164
rect 10134 29016 10140 29028
rect 10095 28988 10140 29016
rect 10134 28976 10140 28988
rect 10192 28976 10198 29028
rect 1104 28858 10856 28880
rect 1104 28806 2582 28858
rect 2634 28806 2646 28858
rect 2698 28806 2710 28858
rect 2762 28806 2774 28858
rect 2826 28806 2838 28858
rect 2890 28806 5846 28858
rect 5898 28806 5910 28858
rect 5962 28806 5974 28858
rect 6026 28806 6038 28858
rect 6090 28806 6102 28858
rect 6154 28806 9110 28858
rect 9162 28806 9174 28858
rect 9226 28806 9238 28858
rect 9290 28806 9302 28858
rect 9354 28806 9366 28858
rect 9418 28806 10856 28858
rect 1104 28784 10856 28806
rect 1949 28747 2007 28753
rect 1949 28713 1961 28747
rect 1995 28744 2007 28747
rect 6454 28744 6460 28756
rect 1995 28716 6460 28744
rect 1995 28713 2007 28716
rect 1949 28707 2007 28713
rect 6454 28704 6460 28716
rect 6512 28704 6518 28756
rect 2866 28636 2872 28688
rect 2924 28676 2930 28688
rect 3050 28676 3056 28688
rect 2924 28648 3056 28676
rect 2924 28636 2930 28648
rect 3050 28636 3056 28648
rect 3108 28636 3114 28688
rect 4062 28676 4068 28688
rect 4023 28648 4068 28676
rect 4062 28636 4068 28648
rect 4120 28636 4126 28688
rect 2777 28611 2835 28617
rect 2777 28577 2789 28611
rect 2823 28608 2835 28611
rect 6362 28608 6368 28620
rect 2823 28580 6368 28608
rect 2823 28577 2835 28580
rect 2777 28571 2835 28577
rect 6362 28568 6368 28580
rect 6420 28568 6426 28620
rect 1857 28543 1915 28549
rect 1857 28509 1869 28543
rect 1903 28540 1915 28543
rect 3050 28540 3056 28552
rect 1903 28512 3056 28540
rect 1903 28509 1915 28512
rect 1857 28503 1915 28509
rect 3050 28500 3056 28512
rect 3108 28500 3114 28552
rect 2593 28475 2651 28481
rect 2593 28441 2605 28475
rect 2639 28472 2651 28475
rect 2639 28444 2774 28472
rect 2639 28441 2651 28444
rect 2593 28435 2651 28441
rect 2746 28404 2774 28444
rect 3326 28432 3332 28484
rect 3384 28472 3390 28484
rect 3881 28475 3939 28481
rect 3881 28472 3893 28475
rect 3384 28444 3893 28472
rect 3384 28432 3390 28444
rect 3881 28441 3893 28444
rect 3927 28441 3939 28475
rect 3881 28435 3939 28441
rect 2958 28404 2964 28416
rect 2746 28376 2964 28404
rect 2958 28364 2964 28376
rect 3016 28364 3022 28416
rect 1104 28314 10856 28336
rect 1104 28262 4214 28314
rect 4266 28262 4278 28314
rect 4330 28262 4342 28314
rect 4394 28262 4406 28314
rect 4458 28262 4470 28314
rect 4522 28262 7478 28314
rect 7530 28262 7542 28314
rect 7594 28262 7606 28314
rect 7658 28262 7670 28314
rect 7722 28262 7734 28314
rect 7786 28262 10856 28314
rect 1104 28240 10856 28262
rect 1394 28160 1400 28212
rect 1452 28200 1458 28212
rect 1670 28200 1676 28212
rect 1452 28172 1676 28200
rect 1452 28160 1458 28172
rect 1670 28160 1676 28172
rect 1728 28160 1734 28212
rect 3053 28203 3111 28209
rect 3053 28169 3065 28203
rect 3099 28200 3111 28203
rect 3142 28200 3148 28212
rect 3099 28172 3148 28200
rect 3099 28169 3111 28172
rect 3053 28163 3111 28169
rect 3142 28160 3148 28172
rect 3200 28160 3206 28212
rect 3326 28160 3332 28212
rect 3384 28200 3390 28212
rect 3602 28200 3608 28212
rect 3384 28172 3608 28200
rect 3384 28160 3390 28172
rect 3602 28160 3608 28172
rect 3660 28160 3666 28212
rect 4249 28203 4307 28209
rect 4249 28169 4261 28203
rect 4295 28200 4307 28203
rect 4982 28200 4988 28212
rect 4295 28172 4988 28200
rect 4295 28169 4307 28172
rect 4249 28163 4307 28169
rect 4982 28160 4988 28172
rect 5040 28160 5046 28212
rect 5350 28160 5356 28212
rect 5408 28200 5414 28212
rect 5408 28172 5488 28200
rect 5408 28160 5414 28172
rect 5460 28144 5488 28172
rect 658 28092 664 28144
rect 716 28132 722 28144
rect 716 28104 2912 28132
rect 716 28092 722 28104
rect 1673 28067 1731 28073
rect 1673 28033 1685 28067
rect 1719 28064 1731 28067
rect 1946 28064 1952 28076
rect 1719 28036 1952 28064
rect 1719 28033 1731 28036
rect 1673 28027 1731 28033
rect 1946 28024 1952 28036
rect 2004 28024 2010 28076
rect 1394 27996 1400 28008
rect 1355 27968 1400 27996
rect 1394 27956 1400 27968
rect 1452 27956 1458 28008
rect 1946 27888 1952 27940
rect 2004 27928 2010 27940
rect 2056 27928 2084 28104
rect 2884 28073 2912 28104
rect 5442 28092 5448 28144
rect 5500 28092 5506 28144
rect 2869 28067 2927 28073
rect 2869 28033 2881 28067
rect 2915 28033 2927 28067
rect 3602 28064 3608 28076
rect 3563 28036 3608 28064
rect 2869 28027 2927 28033
rect 3602 28024 3608 28036
rect 3660 28024 3666 28076
rect 3878 28024 3884 28076
rect 3936 28064 3942 28076
rect 4433 28067 4491 28073
rect 4433 28064 4445 28067
rect 3936 28036 4445 28064
rect 3936 28024 3942 28036
rect 4433 28033 4445 28036
rect 4479 28033 4491 28067
rect 4433 28027 4491 28033
rect 5166 28024 5172 28076
rect 5224 28064 5230 28076
rect 5350 28064 5356 28076
rect 5224 28036 5356 28064
rect 5224 28024 5230 28036
rect 5350 28024 5356 28036
rect 5408 28024 5414 28076
rect 2498 27956 2504 28008
rect 2556 27996 2562 28008
rect 2685 27999 2743 28005
rect 2685 27996 2697 27999
rect 2556 27968 2697 27996
rect 2556 27956 2562 27968
rect 2685 27965 2697 27968
rect 2731 27965 2743 27999
rect 2685 27959 2743 27965
rect 3789 27999 3847 28005
rect 3789 27965 3801 27999
rect 3835 27996 3847 27999
rect 7190 27996 7196 28008
rect 3835 27968 7196 27996
rect 3835 27965 3847 27968
rect 3789 27959 3847 27965
rect 7190 27956 7196 27968
rect 7248 27956 7254 28008
rect 9950 27996 9956 28008
rect 9911 27968 9956 27996
rect 9950 27956 9956 27968
rect 10008 27956 10014 28008
rect 2004 27900 2084 27928
rect 2004 27888 2010 27900
rect 2866 27888 2872 27940
rect 2924 27928 2930 27940
rect 3142 27928 3148 27940
rect 2924 27900 3148 27928
rect 2924 27888 2930 27900
rect 3142 27888 3148 27900
rect 3200 27888 3206 27940
rect 4430 27888 4436 27940
rect 4488 27928 4494 27940
rect 5626 27928 5632 27940
rect 4488 27900 5632 27928
rect 4488 27888 4494 27900
rect 5626 27888 5632 27900
rect 5684 27888 5690 27940
rect 1104 27770 10856 27792
rect 1104 27718 2582 27770
rect 2634 27718 2646 27770
rect 2698 27718 2710 27770
rect 2762 27718 2774 27770
rect 2826 27718 2838 27770
rect 2890 27718 5846 27770
rect 5898 27718 5910 27770
rect 5962 27718 5974 27770
rect 6026 27718 6038 27770
rect 6090 27718 6102 27770
rect 6154 27718 9110 27770
rect 9162 27718 9174 27770
rect 9226 27718 9238 27770
rect 9290 27718 9302 27770
rect 9354 27718 9366 27770
rect 9418 27718 10856 27770
rect 1104 27696 10856 27718
rect 3050 27588 3056 27600
rect 3011 27560 3056 27588
rect 3050 27548 3056 27560
rect 3108 27548 3114 27600
rect 4433 27591 4491 27597
rect 4433 27557 4445 27591
rect 4479 27588 4491 27591
rect 4614 27588 4620 27600
rect 4479 27560 4620 27588
rect 4479 27557 4491 27560
rect 4433 27551 4491 27557
rect 4614 27548 4620 27560
rect 4672 27548 4678 27600
rect 1210 27480 1216 27532
rect 1268 27520 1274 27532
rect 1397 27523 1455 27529
rect 1397 27520 1409 27523
rect 1268 27492 1409 27520
rect 1268 27480 1274 27492
rect 1397 27489 1409 27492
rect 1443 27489 1455 27523
rect 1397 27483 1455 27489
rect 2685 27523 2743 27529
rect 2685 27489 2697 27523
rect 2731 27520 2743 27523
rect 4062 27520 4068 27532
rect 2731 27492 4068 27520
rect 2731 27489 2743 27492
rect 2685 27483 2743 27489
rect 4062 27480 4068 27492
rect 4120 27480 4126 27532
rect 1026 27412 1032 27464
rect 1084 27452 1090 27464
rect 1673 27455 1731 27461
rect 1673 27452 1685 27455
rect 1084 27424 1685 27452
rect 1084 27412 1090 27424
rect 1673 27421 1685 27424
rect 1719 27421 1731 27455
rect 1673 27415 1731 27421
rect 1946 27412 1952 27464
rect 2004 27452 2010 27464
rect 2869 27455 2927 27461
rect 2869 27452 2881 27455
rect 2004 27424 2881 27452
rect 2004 27412 2010 27424
rect 2869 27421 2881 27424
rect 2915 27421 2927 27455
rect 2869 27415 2927 27421
rect 4249 27387 4307 27393
rect 4249 27353 4261 27387
rect 4295 27384 4307 27387
rect 4614 27384 4620 27396
rect 4295 27356 4620 27384
rect 4295 27353 4307 27356
rect 4249 27347 4307 27353
rect 4614 27344 4620 27356
rect 4672 27344 4678 27396
rect 9950 27316 9956 27328
rect 9911 27288 9956 27316
rect 9950 27276 9956 27288
rect 10008 27276 10014 27328
rect 1104 27226 10856 27248
rect 1104 27174 4214 27226
rect 4266 27174 4278 27226
rect 4330 27174 4342 27226
rect 4394 27174 4406 27226
rect 4458 27174 4470 27226
rect 4522 27174 7478 27226
rect 7530 27174 7542 27226
rect 7594 27174 7606 27226
rect 7658 27174 7670 27226
rect 7722 27174 7734 27226
rect 7786 27174 10856 27226
rect 1104 27152 10856 27174
rect 2958 27072 2964 27124
rect 3016 27112 3022 27124
rect 3053 27115 3111 27121
rect 3053 27112 3065 27115
rect 3016 27084 3065 27112
rect 3016 27072 3022 27084
rect 3053 27081 3065 27084
rect 3099 27081 3111 27115
rect 3694 27112 3700 27124
rect 3655 27084 3700 27112
rect 3053 27075 3111 27081
rect 3694 27072 3700 27084
rect 3752 27072 3758 27124
rect 1946 26936 1952 26988
rect 2004 26976 2010 26988
rect 2041 26979 2099 26985
rect 2041 26976 2053 26979
rect 2004 26948 2053 26976
rect 2004 26936 2010 26948
rect 2041 26945 2053 26948
rect 2087 26976 2099 26979
rect 2869 26979 2927 26985
rect 2869 26976 2881 26979
rect 2087 26948 2881 26976
rect 2087 26945 2099 26948
rect 2041 26939 2099 26945
rect 2869 26945 2881 26948
rect 2915 26976 2927 26979
rect 3050 26976 3056 26988
rect 2915 26948 3056 26976
rect 2915 26945 2927 26948
rect 2869 26939 2927 26945
rect 3050 26936 3056 26948
rect 3108 26936 3114 26988
rect 3602 26976 3608 26988
rect 3563 26948 3608 26976
rect 3602 26936 3608 26948
rect 3660 26936 3666 26988
rect 1857 26911 1915 26917
rect 1857 26877 1869 26911
rect 1903 26908 1915 26911
rect 2314 26908 2320 26920
rect 1903 26880 2320 26908
rect 1903 26877 1915 26880
rect 1857 26871 1915 26877
rect 2314 26868 2320 26880
rect 2372 26868 2378 26920
rect 2406 26868 2412 26920
rect 2464 26908 2470 26920
rect 2685 26911 2743 26917
rect 2685 26908 2697 26911
rect 2464 26880 2697 26908
rect 2464 26868 2470 26880
rect 2685 26877 2697 26880
rect 2731 26877 2743 26911
rect 2685 26871 2743 26877
rect 4798 26868 4804 26920
rect 4856 26908 4862 26920
rect 4982 26908 4988 26920
rect 4856 26880 4988 26908
rect 4856 26868 4862 26880
rect 4982 26868 4988 26880
rect 5040 26868 5046 26920
rect 1946 26800 1952 26852
rect 2004 26840 2010 26852
rect 2130 26840 2136 26852
rect 2004 26812 2136 26840
rect 2004 26800 2010 26812
rect 2130 26800 2136 26812
rect 2188 26800 2194 26852
rect 1854 26732 1860 26784
rect 1912 26772 1918 26784
rect 2225 26775 2283 26781
rect 2225 26772 2237 26775
rect 1912 26744 2237 26772
rect 1912 26732 1918 26744
rect 2225 26741 2237 26744
rect 2271 26741 2283 26775
rect 2225 26735 2283 26741
rect 5074 26732 5080 26784
rect 5132 26772 5138 26784
rect 5442 26772 5448 26784
rect 5132 26744 5448 26772
rect 5132 26732 5138 26744
rect 5442 26732 5448 26744
rect 5500 26732 5506 26784
rect 10134 26772 10140 26784
rect 10095 26744 10140 26772
rect 10134 26732 10140 26744
rect 10192 26732 10198 26784
rect 1104 26682 10856 26704
rect 1104 26630 2582 26682
rect 2634 26630 2646 26682
rect 2698 26630 2710 26682
rect 2762 26630 2774 26682
rect 2826 26630 2838 26682
rect 2890 26630 5846 26682
rect 5898 26630 5910 26682
rect 5962 26630 5974 26682
rect 6026 26630 6038 26682
rect 6090 26630 6102 26682
rect 6154 26630 9110 26682
rect 9162 26630 9174 26682
rect 9226 26630 9238 26682
rect 9290 26630 9302 26682
rect 9354 26630 9366 26682
rect 9418 26630 10856 26682
rect 1104 26608 10856 26630
rect 1949 26571 2007 26577
rect 1949 26537 1961 26571
rect 1995 26568 2007 26571
rect 1995 26540 4384 26568
rect 1995 26537 2007 26540
rect 1949 26531 2007 26537
rect 2777 26503 2835 26509
rect 2777 26469 2789 26503
rect 2823 26500 2835 26503
rect 3326 26500 3332 26512
rect 2823 26472 3332 26500
rect 2823 26469 2835 26472
rect 2777 26463 2835 26469
rect 3326 26460 3332 26472
rect 3384 26460 3390 26512
rect 4356 26432 4384 26540
rect 5074 26528 5080 26580
rect 5132 26568 5138 26580
rect 5534 26568 5540 26580
rect 5132 26540 5540 26568
rect 5132 26528 5138 26540
rect 5534 26528 5540 26540
rect 5592 26528 5598 26580
rect 4433 26503 4491 26509
rect 4433 26469 4445 26503
rect 4479 26500 4491 26503
rect 4706 26500 4712 26512
rect 4479 26472 4712 26500
rect 4479 26469 4491 26472
rect 4433 26463 4491 26469
rect 4706 26460 4712 26472
rect 4764 26460 4770 26512
rect 4890 26460 4896 26512
rect 4948 26500 4954 26512
rect 5626 26500 5632 26512
rect 4948 26472 5632 26500
rect 4948 26460 4954 26472
rect 5626 26460 5632 26472
rect 5684 26460 5690 26512
rect 6270 26432 6276 26444
rect 4356 26404 6276 26432
rect 6270 26392 6276 26404
rect 6328 26392 6334 26444
rect 1854 26364 1860 26376
rect 1815 26336 1860 26364
rect 1854 26324 1860 26336
rect 1912 26324 1918 26376
rect 2314 26296 2320 26308
rect 1872 26268 2320 26296
rect 1872 26240 1900 26268
rect 2314 26256 2320 26268
rect 2372 26256 2378 26308
rect 2590 26296 2596 26308
rect 2551 26268 2596 26296
rect 2590 26256 2596 26268
rect 2648 26256 2654 26308
rect 3326 26256 3332 26308
rect 3384 26296 3390 26308
rect 3786 26296 3792 26308
rect 3384 26268 3792 26296
rect 3384 26256 3390 26268
rect 3786 26256 3792 26268
rect 3844 26256 3850 26308
rect 4249 26299 4307 26305
rect 4249 26265 4261 26299
rect 4295 26265 4307 26299
rect 4249 26259 4307 26265
rect 1854 26188 1860 26240
rect 1912 26188 1918 26240
rect 3510 26188 3516 26240
rect 3568 26228 3574 26240
rect 4264 26228 4292 26259
rect 3568 26200 4292 26228
rect 3568 26188 3574 26200
rect 1104 26138 10856 26160
rect 1104 26086 4214 26138
rect 4266 26086 4278 26138
rect 4330 26086 4342 26138
rect 4394 26086 4406 26138
rect 4458 26086 4470 26138
rect 4522 26086 7478 26138
rect 7530 26086 7542 26138
rect 7594 26086 7606 26138
rect 7658 26086 7670 26138
rect 7722 26086 7734 26138
rect 7786 26086 10856 26138
rect 1104 26064 10856 26086
rect 2314 25984 2320 26036
rect 2372 26024 2378 26036
rect 2498 26024 2504 26036
rect 2372 25996 2504 26024
rect 2372 25984 2378 25996
rect 2498 25984 2504 25996
rect 2556 25984 2562 26036
rect 3053 26027 3111 26033
rect 3053 25993 3065 26027
rect 3099 26024 3111 26027
rect 3878 26024 3884 26036
rect 3099 25996 3884 26024
rect 3099 25993 3111 25996
rect 3053 25987 3111 25993
rect 3878 25984 3884 25996
rect 3936 25984 3942 26036
rect 1673 25891 1731 25897
rect 1673 25857 1685 25891
rect 1719 25888 1731 25891
rect 1762 25888 1768 25900
rect 1719 25860 1768 25888
rect 1719 25857 1731 25860
rect 1673 25851 1731 25857
rect 1762 25848 1768 25860
rect 1820 25848 1826 25900
rect 2869 25891 2927 25897
rect 2869 25857 2881 25891
rect 2915 25888 2927 25891
rect 2958 25888 2964 25900
rect 2915 25860 2964 25888
rect 2915 25857 2927 25860
rect 2869 25851 2927 25857
rect 2958 25848 2964 25860
rect 3016 25848 3022 25900
rect 1394 25820 1400 25832
rect 1355 25792 1400 25820
rect 1394 25780 1400 25792
rect 1452 25780 1458 25832
rect 2685 25823 2743 25829
rect 2685 25789 2697 25823
rect 2731 25820 2743 25823
rect 3510 25820 3516 25832
rect 2731 25792 3516 25820
rect 2731 25789 2743 25792
rect 2685 25783 2743 25789
rect 3510 25780 3516 25792
rect 3568 25780 3574 25832
rect 290 25712 296 25764
rect 348 25752 354 25764
rect 1762 25752 1768 25764
rect 348 25724 1768 25752
rect 348 25712 354 25724
rect 1762 25712 1768 25724
rect 1820 25712 1826 25764
rect 10134 25684 10140 25696
rect 10095 25656 10140 25684
rect 10134 25644 10140 25656
rect 10192 25644 10198 25696
rect 1104 25594 10856 25616
rect 1104 25542 2582 25594
rect 2634 25542 2646 25594
rect 2698 25542 2710 25594
rect 2762 25542 2774 25594
rect 2826 25542 2838 25594
rect 2890 25542 5846 25594
rect 5898 25542 5910 25594
rect 5962 25542 5974 25594
rect 6026 25542 6038 25594
rect 6090 25542 6102 25594
rect 6154 25542 9110 25594
rect 9162 25542 9174 25594
rect 9226 25542 9238 25594
rect 9290 25542 9302 25594
rect 9354 25542 9366 25594
rect 9418 25542 10856 25594
rect 1104 25520 10856 25542
rect 3145 25483 3203 25489
rect 3145 25449 3157 25483
rect 3191 25480 3203 25483
rect 3326 25480 3332 25492
rect 3191 25452 3332 25480
rect 3191 25449 3203 25452
rect 3145 25443 3203 25449
rect 3326 25440 3332 25452
rect 3384 25440 3390 25492
rect 1673 25347 1731 25353
rect 1673 25313 1685 25347
rect 1719 25344 1731 25347
rect 4522 25344 4528 25356
rect 1719 25316 4528 25344
rect 1719 25313 1731 25316
rect 1673 25307 1731 25313
rect 4522 25304 4528 25316
rect 4580 25304 4586 25356
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 2777 25279 2835 25285
rect 2777 25245 2789 25279
rect 2823 25245 2835 25279
rect 2958 25276 2964 25288
rect 2919 25248 2964 25276
rect 2777 25239 2835 25245
rect 2498 25168 2504 25220
rect 2556 25208 2562 25220
rect 2792 25208 2820 25239
rect 2958 25236 2964 25248
rect 3016 25276 3022 25288
rect 3694 25276 3700 25288
rect 3016 25248 3700 25276
rect 3016 25236 3022 25248
rect 3694 25236 3700 25248
rect 3752 25236 3758 25288
rect 10134 25276 10140 25288
rect 10095 25248 10140 25276
rect 10134 25236 10140 25248
rect 10192 25236 10198 25288
rect 2556 25180 2820 25208
rect 2556 25168 2562 25180
rect 1104 25050 10856 25072
rect 1104 24998 4214 25050
rect 4266 24998 4278 25050
rect 4330 24998 4342 25050
rect 4394 24998 4406 25050
rect 4458 24998 4470 25050
rect 4522 24998 7478 25050
rect 7530 24998 7542 25050
rect 7594 24998 7606 25050
rect 7658 24998 7670 25050
rect 7722 24998 7734 25050
rect 7786 24998 10856 25050
rect 1104 24976 10856 24998
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24769 1915 24803
rect 1857 24763 1915 24769
rect 2593 24803 2651 24809
rect 2593 24769 2605 24803
rect 2639 24769 2651 24803
rect 2593 24763 2651 24769
rect 1872 24664 1900 24763
rect 2608 24732 2636 24763
rect 2774 24760 2780 24812
rect 2832 24800 2838 24812
rect 3326 24800 3332 24812
rect 2832 24772 2877 24800
rect 3287 24772 3332 24800
rect 2832 24760 2838 24772
rect 3326 24760 3332 24772
rect 3384 24760 3390 24812
rect 3418 24760 3424 24812
rect 3476 24800 3482 24812
rect 3513 24803 3571 24809
rect 3513 24800 3525 24803
rect 3476 24772 3525 24800
rect 3476 24760 3482 24772
rect 3513 24769 3525 24772
rect 3559 24769 3571 24803
rect 3513 24763 3571 24769
rect 4154 24760 4160 24812
rect 4212 24800 4218 24812
rect 4890 24800 4896 24812
rect 4212 24772 4896 24800
rect 4212 24760 4218 24772
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 2958 24732 2964 24744
rect 2608 24704 2964 24732
rect 2958 24692 2964 24704
rect 3016 24692 3022 24744
rect 3142 24692 3148 24744
rect 3200 24732 3206 24744
rect 3200 24704 3372 24732
rect 3200 24692 3206 24704
rect 1872 24636 2360 24664
rect 1118 24556 1124 24608
rect 1176 24596 1182 24608
rect 1949 24599 2007 24605
rect 1949 24596 1961 24599
rect 1176 24568 1961 24596
rect 1176 24556 1182 24568
rect 1949 24565 1961 24568
rect 1995 24565 2007 24599
rect 2332 24596 2360 24636
rect 3344 24608 3372 24704
rect 4614 24624 4620 24676
rect 4672 24664 4678 24676
rect 4890 24664 4896 24676
rect 4672 24636 4896 24664
rect 4672 24624 4678 24636
rect 4890 24624 4896 24636
rect 4948 24624 4954 24676
rect 3142 24596 3148 24608
rect 2332 24568 3148 24596
rect 1949 24559 2007 24565
rect 3142 24556 3148 24568
rect 3200 24556 3206 24608
rect 3326 24556 3332 24608
rect 3384 24556 3390 24608
rect 1104 24506 10856 24528
rect 1104 24454 2582 24506
rect 2634 24454 2646 24506
rect 2698 24454 2710 24506
rect 2762 24454 2774 24506
rect 2826 24454 2838 24506
rect 2890 24454 5846 24506
rect 5898 24454 5910 24506
rect 5962 24454 5974 24506
rect 6026 24454 6038 24506
rect 6090 24454 6102 24506
rect 6154 24454 9110 24506
rect 9162 24454 9174 24506
rect 9226 24454 9238 24506
rect 9290 24454 9302 24506
rect 9354 24454 9366 24506
rect 9418 24454 10856 24506
rect 1104 24432 10856 24454
rect 2866 24284 2872 24336
rect 2924 24324 2930 24336
rect 3050 24324 3056 24336
rect 2924 24296 3056 24324
rect 2924 24284 2930 24296
rect 3050 24284 3056 24296
rect 3108 24284 3114 24336
rect 1673 24259 1731 24265
rect 1673 24225 1685 24259
rect 1719 24256 1731 24259
rect 2038 24256 2044 24268
rect 1719 24228 2044 24256
rect 1719 24225 1731 24228
rect 1673 24219 1731 24225
rect 2038 24216 2044 24228
rect 2096 24216 2102 24268
rect 2961 24259 3019 24265
rect 2961 24225 2973 24259
rect 3007 24256 3019 24259
rect 4154 24256 4160 24268
rect 3007 24228 4160 24256
rect 3007 24225 3019 24228
rect 2961 24219 3019 24225
rect 4154 24216 4160 24228
rect 4212 24216 4218 24268
rect 1394 24188 1400 24200
rect 1355 24160 1400 24188
rect 1394 24148 1400 24160
rect 1452 24148 1458 24200
rect 10134 24188 10140 24200
rect 10095 24160 10140 24188
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 2777 24123 2835 24129
rect 2777 24089 2789 24123
rect 2823 24120 2835 24123
rect 3050 24120 3056 24132
rect 2823 24092 3056 24120
rect 2823 24089 2835 24092
rect 2777 24083 2835 24089
rect 3050 24080 3056 24092
rect 3108 24080 3114 24132
rect 1762 24012 1768 24064
rect 1820 24052 1826 24064
rect 2130 24052 2136 24064
rect 1820 24024 2136 24052
rect 1820 24012 1826 24024
rect 2130 24012 2136 24024
rect 2188 24012 2194 24064
rect 1104 23962 10856 23984
rect 1104 23910 4214 23962
rect 4266 23910 4278 23962
rect 4330 23910 4342 23962
rect 4394 23910 4406 23962
rect 4458 23910 4470 23962
rect 4522 23910 7478 23962
rect 7530 23910 7542 23962
rect 7594 23910 7606 23962
rect 7658 23910 7670 23962
rect 7722 23910 7734 23962
rect 7786 23910 10856 23962
rect 1104 23888 10856 23910
rect 1670 23712 1676 23724
rect 1631 23684 1676 23712
rect 1670 23672 1676 23684
rect 1728 23672 1734 23724
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3970 23712 3976 23724
rect 3007 23684 3976 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 3970 23672 3976 23684
rect 4028 23672 4034 23724
rect 1210 23604 1216 23656
rect 1268 23644 1274 23656
rect 1397 23647 1455 23653
rect 1397 23644 1409 23647
rect 1268 23616 1409 23644
rect 1268 23604 1274 23616
rect 1397 23613 1409 23616
rect 1443 23613 1455 23647
rect 1397 23607 1455 23613
rect 2685 23647 2743 23653
rect 2685 23613 2697 23647
rect 2731 23644 2743 23647
rect 2774 23644 2780 23656
rect 2731 23616 2780 23644
rect 2731 23613 2743 23616
rect 2685 23607 2743 23613
rect 2774 23604 2780 23616
rect 2832 23604 2838 23656
rect 10134 23508 10140 23520
rect 10095 23480 10140 23508
rect 10134 23468 10140 23480
rect 10192 23468 10198 23520
rect 1104 23418 10856 23440
rect 1104 23366 2582 23418
rect 2634 23366 2646 23418
rect 2698 23366 2710 23418
rect 2762 23366 2774 23418
rect 2826 23366 2838 23418
rect 2890 23366 5846 23418
rect 5898 23366 5910 23418
rect 5962 23366 5974 23418
rect 6026 23366 6038 23418
rect 6090 23366 6102 23418
rect 6154 23366 9110 23418
rect 9162 23366 9174 23418
rect 9226 23366 9238 23418
rect 9290 23366 9302 23418
rect 9354 23366 9366 23418
rect 9418 23366 10856 23418
rect 1104 23344 10856 23366
rect 3050 23304 3056 23316
rect 3011 23276 3056 23304
rect 3050 23264 3056 23276
rect 3108 23264 3114 23316
rect 1673 23171 1731 23177
rect 1673 23137 1685 23171
rect 1719 23168 1731 23171
rect 3602 23168 3608 23180
rect 1719 23140 3608 23168
rect 1719 23137 1731 23140
rect 1673 23131 1731 23137
rect 3602 23128 3608 23140
rect 3660 23128 3666 23180
rect 1394 23100 1400 23112
rect 1355 23072 1400 23100
rect 1394 23060 1400 23072
rect 1452 23060 1458 23112
rect 2498 23060 2504 23112
rect 2556 23100 2562 23112
rect 2685 23103 2743 23109
rect 2685 23100 2697 23103
rect 2556 23072 2697 23100
rect 2556 23060 2562 23072
rect 2685 23069 2697 23072
rect 2731 23069 2743 23103
rect 2685 23063 2743 23069
rect 2869 23103 2927 23109
rect 2869 23069 2881 23103
rect 2915 23100 2927 23103
rect 2958 23100 2964 23112
rect 2915 23072 2964 23100
rect 2915 23069 2927 23072
rect 2869 23063 2927 23069
rect 2958 23060 2964 23072
rect 3016 23060 3022 23112
rect 1104 22874 10856 22896
rect 1104 22822 4214 22874
rect 4266 22822 4278 22874
rect 4330 22822 4342 22874
rect 4394 22822 4406 22874
rect 4458 22822 4470 22874
rect 4522 22822 7478 22874
rect 7530 22822 7542 22874
rect 7594 22822 7606 22874
rect 7658 22822 7670 22874
rect 7722 22822 7734 22874
rect 7786 22822 10856 22874
rect 1104 22800 10856 22822
rect 3050 22760 3056 22772
rect 3011 22732 3056 22760
rect 3050 22720 3056 22732
rect 3108 22720 3114 22772
rect 3694 22692 3700 22704
rect 2884 22664 3700 22692
rect 2884 22633 2912 22664
rect 3694 22652 3700 22664
rect 3752 22692 3758 22704
rect 3970 22692 3976 22704
rect 3752 22664 3976 22692
rect 3752 22652 3758 22664
rect 3970 22652 3976 22664
rect 4028 22652 4034 22704
rect 4525 22695 4583 22701
rect 4525 22661 4537 22695
rect 4571 22692 4583 22695
rect 5074 22692 5080 22704
rect 4571 22664 5080 22692
rect 4571 22661 4583 22664
rect 4525 22655 4583 22661
rect 5074 22652 5080 22664
rect 5132 22652 5138 22704
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22624 1731 22627
rect 2869 22627 2927 22633
rect 1719 22596 2820 22624
rect 1719 22593 1731 22596
rect 1673 22587 1731 22593
rect 1210 22516 1216 22568
rect 1268 22556 1274 22568
rect 1397 22559 1455 22565
rect 1397 22556 1409 22559
rect 1268 22528 1409 22556
rect 1268 22516 1274 22528
rect 1397 22525 1409 22528
rect 1443 22525 1455 22559
rect 2685 22559 2743 22565
rect 2685 22556 2697 22559
rect 1397 22519 1455 22525
rect 1688 22528 2697 22556
rect 1688 22500 1716 22528
rect 2685 22525 2697 22528
rect 2731 22525 2743 22559
rect 2792 22556 2820 22596
rect 2869 22593 2881 22627
rect 2915 22593 2927 22627
rect 3602 22624 3608 22636
rect 3563 22596 3608 22624
rect 2869 22587 2927 22593
rect 3602 22584 3608 22596
rect 3660 22584 3666 22636
rect 4154 22584 4160 22636
rect 4212 22624 4218 22636
rect 4341 22627 4399 22633
rect 4341 22624 4353 22627
rect 4212 22596 4353 22624
rect 4212 22584 4218 22596
rect 4341 22593 4353 22596
rect 4387 22593 4399 22627
rect 4341 22587 4399 22593
rect 3418 22556 3424 22568
rect 2792 22528 3424 22556
rect 2685 22519 2743 22525
rect 3418 22516 3424 22528
rect 3476 22516 3482 22568
rect 1670 22448 1676 22500
rect 1728 22448 1734 22500
rect 10134 22488 10140 22500
rect 10095 22460 10140 22488
rect 10134 22448 10140 22460
rect 10192 22448 10198 22500
rect 3694 22420 3700 22432
rect 3655 22392 3700 22420
rect 3694 22380 3700 22392
rect 3752 22380 3758 22432
rect 1104 22330 10856 22352
rect 934 22244 940 22296
rect 992 22244 998 22296
rect 1104 22278 2582 22330
rect 2634 22278 2646 22330
rect 2698 22278 2710 22330
rect 2762 22278 2774 22330
rect 2826 22278 2838 22330
rect 2890 22278 5846 22330
rect 5898 22278 5910 22330
rect 5962 22278 5974 22330
rect 6026 22278 6038 22330
rect 6090 22278 6102 22330
rect 6154 22278 9110 22330
rect 9162 22278 9174 22330
rect 9226 22278 9238 22330
rect 9290 22278 9302 22330
rect 9354 22278 9366 22330
rect 9418 22278 10856 22330
rect 1104 22256 10856 22278
rect 952 22216 980 22244
rect 952 22188 2360 22216
rect 2332 22160 2360 22188
rect 2498 22176 2504 22228
rect 2556 22216 2562 22228
rect 2556 22188 2728 22216
rect 2556 22176 2562 22188
rect 2700 22160 2728 22188
rect 934 22108 940 22160
rect 992 22148 998 22160
rect 1762 22148 1768 22160
rect 992 22120 1768 22148
rect 992 22108 998 22120
rect 1762 22108 1768 22120
rect 1820 22108 1826 22160
rect 2314 22108 2320 22160
rect 2372 22108 2378 22160
rect 2682 22108 2688 22160
rect 2740 22108 2746 22160
rect 10134 22148 10140 22160
rect 10095 22120 10140 22148
rect 10134 22108 10140 22120
rect 10192 22108 10198 22160
rect 1486 22040 1492 22092
rect 1544 22080 1550 22092
rect 1673 22083 1731 22089
rect 1673 22080 1685 22083
rect 1544 22052 1685 22080
rect 1544 22040 1550 22052
rect 1673 22049 1685 22052
rect 1719 22049 1731 22083
rect 1673 22043 1731 22049
rect 2222 22040 2228 22092
rect 2280 22080 2286 22092
rect 2590 22080 2596 22092
rect 2280 22052 2596 22080
rect 2280 22040 2286 22052
rect 2590 22040 2596 22052
rect 2648 22040 2654 22092
rect 3053 22083 3111 22089
rect 3053 22049 3065 22083
rect 3099 22080 3111 22083
rect 3142 22080 3148 22092
rect 3099 22052 3148 22080
rect 3099 22049 3111 22052
rect 3053 22043 3111 22049
rect 3142 22040 3148 22052
rect 3200 22040 3206 22092
rect 4157 22083 4215 22089
rect 4157 22049 4169 22083
rect 4203 22080 4215 22083
rect 4614 22080 4620 22092
rect 4203 22052 4620 22080
rect 4203 22049 4215 22052
rect 4157 22043 4215 22049
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 1394 22012 1400 22024
rect 1355 21984 1400 22012
rect 1394 21972 1400 21984
rect 1452 21972 1458 22024
rect 2038 21972 2044 22024
rect 2096 22012 2102 22024
rect 2685 22015 2743 22021
rect 2685 22012 2697 22015
rect 2096 21984 2697 22012
rect 2096 21972 2102 21984
rect 2685 21981 2697 21984
rect 2731 21981 2743 22015
rect 2685 21975 2743 21981
rect 2869 22015 2927 22021
rect 2869 21981 2881 22015
rect 2915 22012 2927 22015
rect 2958 22012 2964 22024
rect 2915 21984 2964 22012
rect 2915 21981 2927 21984
rect 2869 21975 2927 21981
rect 2700 21944 2728 21975
rect 2958 21972 2964 21984
rect 3016 21972 3022 22024
rect 3789 22015 3847 22021
rect 3789 21981 3801 22015
rect 3835 21981 3847 22015
rect 3970 22012 3976 22024
rect 3931 21984 3976 22012
rect 3789 21975 3847 21981
rect 3804 21944 3832 21975
rect 3970 21972 3976 21984
rect 4028 21972 4034 22024
rect 2700 21916 3832 21944
rect 1104 21786 10856 21808
rect 1104 21734 4214 21786
rect 4266 21734 4278 21786
rect 4330 21734 4342 21786
rect 4394 21734 4406 21786
rect 4458 21734 4470 21786
rect 4522 21734 7478 21786
rect 7530 21734 7542 21786
rect 7594 21734 7606 21786
rect 7658 21734 7670 21786
rect 7722 21734 7734 21786
rect 7786 21734 10856 21786
rect 1104 21712 10856 21734
rect 3973 21675 4031 21681
rect 3973 21641 3985 21675
rect 4019 21672 4031 21675
rect 4062 21672 4068 21684
rect 4019 21644 4068 21672
rect 4019 21641 4031 21644
rect 3973 21635 4031 21641
rect 4062 21632 4068 21644
rect 4120 21632 4126 21684
rect 934 21564 940 21616
rect 992 21604 998 21616
rect 2777 21607 2835 21613
rect 2777 21604 2789 21607
rect 992 21576 2789 21604
rect 992 21564 998 21576
rect 2777 21573 2789 21576
rect 2823 21604 2835 21607
rect 4798 21604 4804 21616
rect 2823 21576 4804 21604
rect 2823 21573 2835 21576
rect 2777 21567 2835 21573
rect 4798 21564 4804 21576
rect 4856 21564 4862 21616
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 2314 21536 2320 21548
rect 1719 21508 2320 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 2314 21496 2320 21508
rect 2372 21496 2378 21548
rect 2958 21496 2964 21548
rect 3016 21536 3022 21548
rect 3789 21539 3847 21545
rect 3789 21536 3801 21539
rect 3016 21508 3801 21536
rect 3016 21496 3022 21508
rect 3789 21505 3801 21508
rect 3835 21505 3847 21539
rect 3789 21499 3847 21505
rect 1394 21468 1400 21480
rect 1355 21440 1400 21468
rect 1394 21428 1400 21440
rect 1452 21428 1458 21480
rect 1762 21428 1768 21480
rect 1820 21468 1826 21480
rect 2682 21468 2688 21480
rect 1820 21440 2688 21468
rect 1820 21428 1826 21440
rect 2682 21428 2688 21440
rect 2740 21428 2746 21480
rect 3418 21428 3424 21480
rect 3476 21468 3482 21480
rect 3605 21471 3663 21477
rect 3605 21468 3617 21471
rect 3476 21440 3617 21468
rect 3476 21428 3482 21440
rect 3605 21437 3617 21440
rect 3651 21437 3663 21471
rect 3605 21431 3663 21437
rect 2314 21360 2320 21412
rect 2372 21400 2378 21412
rect 2590 21400 2596 21412
rect 2372 21372 2596 21400
rect 2372 21360 2378 21372
rect 2590 21360 2596 21372
rect 2648 21360 2654 21412
rect 2958 21400 2964 21412
rect 2919 21372 2964 21400
rect 2958 21360 2964 21372
rect 3016 21360 3022 21412
rect 10134 21332 10140 21344
rect 10095 21304 10140 21332
rect 10134 21292 10140 21304
rect 10192 21292 10198 21344
rect 1104 21242 10856 21264
rect 1104 21190 2582 21242
rect 2634 21190 2646 21242
rect 2698 21190 2710 21242
rect 2762 21190 2774 21242
rect 2826 21190 2838 21242
rect 2890 21190 5846 21242
rect 5898 21190 5910 21242
rect 5962 21190 5974 21242
rect 6026 21190 6038 21242
rect 6090 21190 6102 21242
rect 6154 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 9238 21242
rect 9290 21190 9302 21242
rect 9354 21190 9366 21242
rect 9418 21190 10856 21242
rect 1104 21168 10856 21190
rect 3053 21131 3111 21137
rect 3053 21097 3065 21131
rect 3099 21128 3111 21131
rect 3602 21128 3608 21140
rect 3099 21100 3608 21128
rect 3099 21097 3111 21100
rect 3053 21091 3111 21097
rect 3602 21088 3608 21100
rect 3660 21088 3666 21140
rect 1673 20995 1731 21001
rect 1673 20961 1685 20995
rect 1719 20992 1731 20995
rect 2406 20992 2412 21004
rect 1719 20964 2412 20992
rect 1719 20961 1731 20964
rect 1673 20955 1731 20961
rect 2406 20952 2412 20964
rect 2464 20952 2470 21004
rect 1394 20924 1400 20936
rect 1355 20896 1400 20924
rect 1394 20884 1400 20896
rect 1452 20884 1458 20936
rect 1578 20884 1584 20936
rect 1636 20924 1642 20936
rect 2685 20927 2743 20933
rect 2685 20924 2697 20927
rect 1636 20896 2697 20924
rect 1636 20884 1642 20896
rect 2685 20893 2697 20896
rect 2731 20893 2743 20927
rect 2685 20887 2743 20893
rect 2869 20927 2927 20933
rect 2869 20893 2881 20927
rect 2915 20924 2927 20927
rect 2958 20924 2964 20936
rect 2915 20896 2964 20924
rect 2915 20893 2927 20896
rect 2869 20887 2927 20893
rect 2958 20884 2964 20896
rect 3016 20884 3022 20936
rect 1104 20698 10856 20720
rect 1104 20646 4214 20698
rect 4266 20646 4278 20698
rect 4330 20646 4342 20698
rect 4394 20646 4406 20698
rect 4458 20646 4470 20698
rect 4522 20646 7478 20698
rect 7530 20646 7542 20698
rect 7594 20646 7606 20698
rect 7658 20646 7670 20698
rect 7722 20646 7734 20698
rect 7786 20646 10856 20698
rect 1104 20624 10856 20646
rect 3053 20587 3111 20593
rect 3053 20553 3065 20587
rect 3099 20584 3111 20587
rect 7834 20584 7840 20596
rect 3099 20556 7840 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 7834 20544 7840 20556
rect 7892 20544 7898 20596
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20448 1731 20451
rect 2222 20448 2228 20460
rect 1719 20420 2228 20448
rect 1719 20417 1731 20420
rect 1673 20411 1731 20417
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 2869 20451 2927 20457
rect 2869 20417 2881 20451
rect 2915 20448 2927 20451
rect 3602 20448 3608 20460
rect 2915 20420 3608 20448
rect 2915 20417 2927 20420
rect 2869 20411 2927 20417
rect 3602 20408 3608 20420
rect 3660 20448 3666 20460
rect 3970 20448 3976 20460
rect 3660 20420 3976 20448
rect 3660 20408 3666 20420
rect 3970 20408 3976 20420
rect 4028 20408 4034 20460
rect 9766 20408 9772 20460
rect 9824 20448 9830 20460
rect 9861 20451 9919 20457
rect 9861 20448 9873 20451
rect 9824 20420 9873 20448
rect 9824 20408 9830 20420
rect 9861 20417 9873 20420
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 1762 20340 1768 20392
rect 1820 20380 1826 20392
rect 2685 20383 2743 20389
rect 2685 20380 2697 20383
rect 1820 20352 2697 20380
rect 1820 20340 1826 20352
rect 2685 20349 2697 20352
rect 2731 20349 2743 20383
rect 2685 20343 2743 20349
rect 10042 20312 10048 20324
rect 10003 20284 10048 20312
rect 10042 20272 10048 20284
rect 10100 20272 10106 20324
rect 1104 20154 10856 20176
rect 1104 20102 2582 20154
rect 2634 20102 2646 20154
rect 2698 20102 2710 20154
rect 2762 20102 2774 20154
rect 2826 20102 2838 20154
rect 2890 20102 5846 20154
rect 5898 20102 5910 20154
rect 5962 20102 5974 20154
rect 6026 20102 6038 20154
rect 6090 20102 6102 20154
rect 6154 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 9238 20154
rect 9290 20102 9302 20154
rect 9354 20102 9366 20154
rect 9418 20102 10856 20154
rect 1104 20080 10856 20102
rect 2498 20000 2504 20052
rect 2556 20040 2562 20052
rect 2593 20043 2651 20049
rect 2593 20040 2605 20043
rect 2556 20012 2605 20040
rect 2556 20000 2562 20012
rect 2593 20009 2605 20012
rect 2639 20009 2651 20043
rect 2593 20003 2651 20009
rect 3789 20043 3847 20049
rect 3789 20009 3801 20043
rect 3835 20040 3847 20043
rect 3878 20040 3884 20052
rect 3835 20012 3884 20040
rect 3835 20009 3847 20012
rect 3789 20003 3847 20009
rect 3878 20000 3884 20012
rect 3936 20000 3942 20052
rect 1854 19932 1860 19984
rect 1912 19972 1918 19984
rect 2406 19972 2412 19984
rect 1912 19944 2412 19972
rect 1912 19932 1918 19944
rect 2406 19932 2412 19944
rect 2464 19932 2470 19984
rect 2958 19904 2964 19916
rect 1964 19876 2964 19904
rect 1762 19836 1768 19848
rect 1723 19808 1768 19836
rect 1762 19796 1768 19808
rect 1820 19796 1826 19848
rect 1964 19845 1992 19876
rect 2958 19864 2964 19876
rect 3016 19864 3022 19916
rect 1949 19839 2007 19845
rect 1949 19805 1961 19839
rect 1995 19805 2007 19839
rect 1949 19799 2007 19805
rect 2777 19839 2835 19845
rect 2777 19805 2789 19839
rect 2823 19836 2835 19839
rect 2866 19836 2872 19848
rect 2823 19808 2872 19836
rect 2823 19805 2835 19808
rect 2777 19799 2835 19805
rect 2866 19796 2872 19808
rect 2924 19796 2930 19848
rect 3970 19836 3976 19848
rect 3931 19808 3976 19836
rect 3970 19796 3976 19808
rect 4028 19796 4034 19848
rect 9858 19836 9864 19848
rect 9819 19808 9864 19836
rect 9858 19796 9864 19808
rect 9916 19796 9922 19848
rect 1854 19660 1860 19712
rect 1912 19700 1918 19712
rect 2133 19703 2191 19709
rect 2133 19700 2145 19703
rect 1912 19672 2145 19700
rect 1912 19660 1918 19672
rect 2133 19669 2145 19672
rect 2179 19669 2191 19703
rect 10042 19700 10048 19712
rect 10003 19672 10048 19700
rect 2133 19663 2191 19669
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 1104 19610 10856 19632
rect 1104 19558 4214 19610
rect 4266 19558 4278 19610
rect 4330 19558 4342 19610
rect 4394 19558 4406 19610
rect 4458 19558 4470 19610
rect 4522 19558 7478 19610
rect 7530 19558 7542 19610
rect 7594 19558 7606 19610
rect 7658 19558 7670 19610
rect 7722 19558 7734 19610
rect 7786 19558 10856 19610
rect 1104 19536 10856 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 2406 19456 2412 19508
rect 2464 19496 2470 19508
rect 2501 19499 2559 19505
rect 2501 19496 2513 19499
rect 2464 19468 2513 19496
rect 2464 19456 2470 19468
rect 2501 19465 2513 19468
rect 2547 19465 2559 19499
rect 9858 19496 9864 19508
rect 9819 19468 9864 19496
rect 2501 19459 2559 19465
rect 9858 19456 9864 19468
rect 9916 19456 9922 19508
rect 1854 19428 1860 19440
rect 1815 19400 1860 19428
rect 1854 19388 1860 19400
rect 1912 19388 1918 19440
rect 2424 19400 10088 19428
rect 2424 19372 2452 19400
rect 2406 19320 2412 19372
rect 2464 19320 2470 19372
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19360 2743 19363
rect 2774 19360 2780 19372
rect 2731 19332 2780 19360
rect 2731 19329 2743 19332
rect 2685 19323 2743 19329
rect 2774 19320 2780 19332
rect 2832 19320 2838 19372
rect 3142 19320 3148 19372
rect 3200 19360 3206 19372
rect 5442 19360 5448 19372
rect 3200 19332 5448 19360
rect 3200 19320 3206 19332
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 10060 19369 10088 19400
rect 10045 19363 10103 19369
rect 10045 19329 10057 19363
rect 10091 19329 10103 19363
rect 10045 19323 10103 19329
rect 1394 19116 1400 19168
rect 1452 19156 1458 19168
rect 1670 19156 1676 19168
rect 1452 19128 1676 19156
rect 1452 19116 1458 19128
rect 1670 19116 1676 19128
rect 1728 19116 1734 19168
rect 1104 19066 10856 19088
rect 1104 19014 2582 19066
rect 2634 19014 2646 19066
rect 2698 19014 2710 19066
rect 2762 19014 2774 19066
rect 2826 19014 2838 19066
rect 2890 19014 5846 19066
rect 5898 19014 5910 19066
rect 5962 19014 5974 19066
rect 6026 19014 6038 19066
rect 6090 19014 6102 19066
rect 6154 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 9238 19066
rect 9290 19014 9302 19066
rect 9354 19014 9366 19066
rect 9418 19014 10856 19066
rect 1104 18992 10856 19014
rect 1397 18955 1455 18961
rect 1397 18921 1409 18955
rect 1443 18952 1455 18955
rect 1578 18952 1584 18964
rect 1443 18924 1584 18952
rect 1443 18921 1455 18924
rect 1397 18915 1455 18921
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 2038 18952 2044 18964
rect 1999 18924 2044 18952
rect 2038 18912 2044 18924
rect 2096 18912 2102 18964
rect 2685 18955 2743 18961
rect 2685 18921 2697 18955
rect 2731 18952 2743 18955
rect 3418 18952 3424 18964
rect 2731 18924 3424 18952
rect 2731 18921 2743 18924
rect 2685 18915 2743 18921
rect 3418 18912 3424 18924
rect 3476 18912 3482 18964
rect 1486 18708 1492 18760
rect 1544 18748 1550 18760
rect 1581 18751 1639 18757
rect 1581 18748 1593 18751
rect 1544 18720 1593 18748
rect 1544 18708 1550 18720
rect 1581 18717 1593 18720
rect 1627 18717 1639 18751
rect 2222 18748 2228 18760
rect 2183 18720 2228 18748
rect 1581 18711 1639 18717
rect 2222 18708 2228 18720
rect 2280 18708 2286 18760
rect 2866 18748 2872 18760
rect 2827 18720 2872 18748
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 9214 18708 9220 18760
rect 9272 18748 9278 18760
rect 9861 18751 9919 18757
rect 9861 18748 9873 18751
rect 9272 18720 9873 18748
rect 9272 18708 9278 18720
rect 9861 18717 9873 18720
rect 9907 18717 9919 18751
rect 9861 18711 9919 18717
rect 10042 18612 10048 18624
rect 10003 18584 10048 18612
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 1104 18522 10856 18544
rect 1104 18470 4214 18522
rect 4266 18470 4278 18522
rect 4330 18470 4342 18522
rect 4394 18470 4406 18522
rect 4458 18470 4470 18522
rect 4522 18470 7478 18522
rect 7530 18470 7542 18522
rect 7594 18470 7606 18522
rect 7658 18470 7670 18522
rect 7722 18470 7734 18522
rect 7786 18470 10856 18522
rect 1104 18448 10856 18470
rect 1394 18408 1400 18420
rect 1355 18380 1400 18408
rect 1394 18368 1400 18380
rect 1452 18368 1458 18420
rect 9214 18408 9220 18420
rect 9175 18380 9220 18408
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 1026 18300 1032 18352
rect 1084 18340 1090 18352
rect 2317 18343 2375 18349
rect 2317 18340 2329 18343
rect 1084 18312 2329 18340
rect 1084 18300 1090 18312
rect 2317 18309 2329 18312
rect 2363 18340 2375 18343
rect 2406 18340 2412 18352
rect 2363 18312 2412 18340
rect 2363 18309 2375 18312
rect 2317 18303 2375 18309
rect 2406 18300 2412 18312
rect 2464 18300 2470 18352
rect 2533 18343 2591 18349
rect 2533 18309 2545 18343
rect 2579 18340 2591 18343
rect 5442 18340 5448 18352
rect 2579 18312 5448 18340
rect 2579 18309 2591 18312
rect 2533 18303 2591 18309
rect 5442 18300 5448 18312
rect 5500 18300 5506 18352
rect 1394 18232 1400 18284
rect 1452 18272 1458 18284
rect 1581 18275 1639 18281
rect 1581 18272 1593 18275
rect 1452 18244 1593 18272
rect 1452 18232 1458 18244
rect 1581 18241 1593 18244
rect 1627 18241 1639 18275
rect 9401 18275 9459 18281
rect 9401 18272 9413 18275
rect 1581 18235 1639 18241
rect 2746 18244 9413 18272
rect 2746 18136 2774 18244
rect 9401 18241 9413 18244
rect 9447 18241 9459 18275
rect 9858 18272 9864 18284
rect 9819 18244 9864 18272
rect 9401 18235 9459 18241
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 2516 18108 2774 18136
rect 1854 18028 1860 18080
rect 1912 18068 1918 18080
rect 2516 18077 2544 18108
rect 2501 18071 2559 18077
rect 2501 18068 2513 18071
rect 1912 18040 2513 18068
rect 1912 18028 1918 18040
rect 2501 18037 2513 18040
rect 2547 18037 2559 18071
rect 2501 18031 2559 18037
rect 2685 18071 2743 18077
rect 2685 18037 2697 18071
rect 2731 18068 2743 18071
rect 2958 18068 2964 18080
rect 2731 18040 2964 18068
rect 2731 18037 2743 18040
rect 2685 18031 2743 18037
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 10042 18068 10048 18080
rect 10003 18040 10048 18068
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 1104 17978 10856 18000
rect 1104 17926 2582 17978
rect 2634 17926 2646 17978
rect 2698 17926 2710 17978
rect 2762 17926 2774 17978
rect 2826 17926 2838 17978
rect 2890 17926 5846 17978
rect 5898 17926 5910 17978
rect 5962 17926 5974 17978
rect 6026 17926 6038 17978
rect 6090 17926 6102 17978
rect 6154 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 9238 17978
rect 9290 17926 9302 17978
rect 9354 17926 9366 17978
rect 9418 17926 10856 17978
rect 1104 17904 10856 17926
rect 1397 17867 1455 17873
rect 1397 17833 1409 17867
rect 1443 17864 1455 17867
rect 1762 17864 1768 17876
rect 1443 17836 1768 17864
rect 1443 17833 1455 17836
rect 1397 17827 1455 17833
rect 1762 17824 1768 17836
rect 1820 17824 1826 17876
rect 2409 17799 2467 17805
rect 2409 17765 2421 17799
rect 2455 17796 2467 17799
rect 3786 17796 3792 17808
rect 2455 17768 3792 17796
rect 2455 17765 2467 17768
rect 2409 17759 2467 17765
rect 3786 17756 3792 17768
rect 3844 17756 3850 17808
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 4893 17731 4951 17737
rect 4893 17728 4905 17731
rect 4856 17700 4905 17728
rect 4856 17688 4862 17700
rect 4893 17697 4905 17700
rect 4939 17697 4951 17731
rect 4893 17691 4951 17697
rect 1578 17660 1584 17672
rect 1539 17632 1584 17660
rect 1578 17620 1584 17632
rect 1636 17620 1642 17672
rect 2222 17660 2228 17672
rect 2183 17632 2228 17660
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 2774 17620 2780 17672
rect 2832 17660 2838 17672
rect 2832 17632 2877 17660
rect 2832 17620 2838 17632
rect 2958 17620 2964 17672
rect 3016 17660 3022 17672
rect 3016 17632 3061 17660
rect 3016 17620 3022 17632
rect 9490 17620 9496 17672
rect 9548 17660 9554 17672
rect 9861 17663 9919 17669
rect 9861 17660 9873 17663
rect 9548 17632 9873 17660
rect 9548 17620 9554 17632
rect 9861 17629 9873 17632
rect 9907 17629 9919 17663
rect 9861 17623 9919 17629
rect 3050 17552 3056 17604
rect 3108 17592 3114 17604
rect 4157 17595 4215 17601
rect 4157 17592 4169 17595
rect 3108 17564 4169 17592
rect 3108 17552 3114 17564
rect 4157 17561 4169 17564
rect 4203 17561 4215 17595
rect 4157 17555 4215 17561
rect 10042 17524 10048 17536
rect 10003 17496 10048 17524
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 1104 17434 10856 17456
rect 1104 17382 4214 17434
rect 4266 17382 4278 17434
rect 4330 17382 4342 17434
rect 4394 17382 4406 17434
rect 4458 17382 4470 17434
rect 4522 17382 7478 17434
rect 7530 17382 7542 17434
rect 7594 17382 7606 17434
rect 7658 17382 7670 17434
rect 7722 17382 7734 17434
rect 7786 17382 10856 17434
rect 1104 17360 10856 17382
rect 3050 17320 3056 17332
rect 3011 17292 3056 17320
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 9953 17323 10011 17329
rect 9953 17320 9965 17323
rect 9916 17292 9965 17320
rect 9916 17280 9922 17292
rect 9953 17289 9965 17292
rect 9999 17289 10011 17323
rect 9953 17283 10011 17289
rect 2869 17255 2927 17261
rect 2869 17221 2881 17255
rect 2915 17252 2927 17255
rect 2958 17252 2964 17264
rect 2915 17224 2964 17252
rect 2915 17221 2927 17224
rect 2869 17215 2927 17221
rect 2958 17212 2964 17224
rect 3016 17212 3022 17264
rect 1486 17144 1492 17196
rect 1544 17184 1550 17196
rect 1581 17187 1639 17193
rect 1581 17184 1593 17187
rect 1544 17156 1593 17184
rect 1544 17144 1550 17156
rect 1581 17153 1593 17156
rect 1627 17153 1639 17187
rect 1581 17147 1639 17153
rect 4614 17144 4620 17196
rect 4672 17184 4678 17196
rect 5442 17184 5448 17196
rect 4672 17156 5448 17184
rect 4672 17144 4678 17156
rect 5442 17144 5448 17156
rect 5500 17184 5506 17196
rect 10137 17187 10195 17193
rect 10137 17184 10149 17187
rect 5500 17156 10149 17184
rect 5500 17144 5506 17156
rect 10137 17153 10149 17156
rect 10183 17153 10195 17187
rect 10137 17147 10195 17153
rect 2222 17008 2228 17060
rect 2280 17048 2286 17060
rect 2501 17051 2559 17057
rect 2501 17048 2513 17051
rect 2280 17020 2513 17048
rect 2280 17008 2286 17020
rect 2501 17017 2513 17020
rect 2547 17017 2559 17051
rect 2501 17011 2559 17017
rect 2774 17008 2780 17060
rect 2832 17048 2838 17060
rect 2832 17020 2912 17048
rect 2832 17008 2838 17020
rect 1394 16980 1400 16992
rect 1355 16952 1400 16980
rect 1394 16940 1400 16952
rect 1452 16940 1458 16992
rect 2884 16989 2912 17020
rect 2869 16983 2927 16989
rect 2869 16949 2881 16983
rect 2915 16949 2927 16983
rect 2869 16943 2927 16949
rect 1104 16890 10856 16912
rect 1104 16838 2582 16890
rect 2634 16838 2646 16890
rect 2698 16838 2710 16890
rect 2762 16838 2774 16890
rect 2826 16838 2838 16890
rect 2890 16838 5846 16890
rect 5898 16838 5910 16890
rect 5962 16838 5974 16890
rect 6026 16838 6038 16890
rect 6090 16838 6102 16890
rect 6154 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 9238 16890
rect 9290 16838 9302 16890
rect 9354 16838 9366 16890
rect 9418 16838 10856 16890
rect 1104 16816 10856 16838
rect 1949 16779 2007 16785
rect 1949 16745 1961 16779
rect 1995 16776 2007 16779
rect 5350 16776 5356 16788
rect 1995 16748 5356 16776
rect 1995 16745 2007 16748
rect 1949 16739 2007 16745
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 1578 16668 1584 16720
rect 1636 16708 1642 16720
rect 1854 16708 1860 16720
rect 1636 16680 1860 16708
rect 1636 16668 1642 16680
rect 1854 16668 1860 16680
rect 1912 16668 1918 16720
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 5166 16640 5172 16652
rect 2924 16612 5172 16640
rect 2924 16600 2930 16612
rect 5166 16600 5172 16612
rect 5224 16600 5230 16652
rect 2685 16575 2743 16581
rect 2685 16541 2697 16575
rect 2731 16572 2743 16575
rect 2774 16572 2780 16584
rect 2731 16544 2780 16572
rect 2731 16541 2743 16544
rect 2685 16535 2743 16541
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 3970 16572 3976 16584
rect 3931 16544 3976 16572
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 9861 16575 9919 16581
rect 9861 16541 9873 16575
rect 9907 16572 9919 16575
rect 9950 16572 9956 16584
rect 9907 16544 9956 16572
rect 9907 16541 9919 16544
rect 9861 16535 9919 16541
rect 9950 16532 9956 16544
rect 10008 16532 10014 16584
rect 1857 16507 1915 16513
rect 1857 16473 1869 16507
rect 1903 16504 1915 16507
rect 2038 16504 2044 16516
rect 1903 16476 2044 16504
rect 1903 16473 1915 16476
rect 1857 16467 1915 16473
rect 2038 16464 2044 16476
rect 2096 16464 2102 16516
rect 2498 16436 2504 16448
rect 2459 16408 2504 16436
rect 2498 16396 2504 16408
rect 2556 16396 2562 16448
rect 3786 16436 3792 16448
rect 3747 16408 3792 16436
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 10042 16436 10048 16448
rect 10003 16408 10048 16436
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 1104 16346 10856 16368
rect 1104 16294 4214 16346
rect 4266 16294 4278 16346
rect 4330 16294 4342 16346
rect 4394 16294 4406 16346
rect 4458 16294 4470 16346
rect 4522 16294 7478 16346
rect 7530 16294 7542 16346
rect 7594 16294 7606 16346
rect 7658 16294 7670 16346
rect 7722 16294 7734 16346
rect 7786 16294 10856 16346
rect 1104 16272 10856 16294
rect 2777 16235 2835 16241
rect 2777 16201 2789 16235
rect 2823 16232 2835 16235
rect 2866 16232 2872 16244
rect 2823 16204 2872 16232
rect 2823 16201 2835 16204
rect 2777 16195 2835 16201
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 9217 16235 9275 16241
rect 9217 16201 9229 16235
rect 9263 16232 9275 16235
rect 9490 16232 9496 16244
rect 9263 16204 9496 16232
rect 9263 16201 9275 16204
rect 9217 16195 9275 16201
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 3786 16164 3792 16176
rect 1964 16136 3792 16164
rect 1394 16056 1400 16108
rect 1452 16096 1458 16108
rect 1964 16105 1992 16136
rect 3786 16124 3792 16136
rect 3844 16124 3850 16176
rect 1489 16099 1547 16105
rect 1489 16096 1501 16099
rect 1452 16068 1501 16096
rect 1452 16056 1458 16068
rect 1489 16065 1501 16068
rect 1535 16065 1547 16099
rect 1489 16059 1547 16065
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16065 1639 16099
rect 1581 16059 1639 16065
rect 1949 16099 2007 16105
rect 1949 16065 1961 16099
rect 1995 16065 2007 16099
rect 1949 16059 2007 16065
rect 2593 16099 2651 16105
rect 2593 16065 2605 16099
rect 2639 16096 2651 16099
rect 4062 16096 4068 16108
rect 2639 16068 4068 16096
rect 2639 16065 2651 16068
rect 2593 16059 2651 16065
rect 1596 16028 1624 16059
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 6178 16056 6184 16108
rect 6236 16096 6242 16108
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 6236 16068 9413 16096
rect 6236 16056 6242 16068
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 9674 16056 9680 16108
rect 9732 16096 9738 16108
rect 9861 16099 9919 16105
rect 9861 16096 9873 16099
rect 9732 16068 9873 16096
rect 9732 16056 9738 16068
rect 9861 16065 9873 16068
rect 9907 16065 9919 16099
rect 9861 16059 9919 16065
rect 3786 16028 3792 16040
rect 1596 16000 3792 16028
rect 3786 15988 3792 16000
rect 3844 15988 3850 16040
rect 2498 15960 2504 15972
rect 1872 15932 2504 15960
rect 1872 15901 1900 15932
rect 2498 15920 2504 15932
rect 2556 15920 2562 15972
rect 1857 15895 1915 15901
rect 1857 15861 1869 15895
rect 1903 15861 1915 15895
rect 1857 15855 1915 15861
rect 1946 15852 1952 15904
rect 2004 15892 2010 15904
rect 2133 15895 2191 15901
rect 2133 15892 2145 15895
rect 2004 15864 2145 15892
rect 2004 15852 2010 15864
rect 2133 15861 2145 15864
rect 2179 15861 2191 15895
rect 10042 15892 10048 15904
rect 10003 15864 10048 15892
rect 2133 15855 2191 15861
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 1104 15802 10856 15824
rect 1104 15750 2582 15802
rect 2634 15750 2646 15802
rect 2698 15750 2710 15802
rect 2762 15750 2774 15802
rect 2826 15750 2838 15802
rect 2890 15750 5846 15802
rect 5898 15750 5910 15802
rect 5962 15750 5974 15802
rect 6026 15750 6038 15802
rect 6090 15750 6102 15802
rect 6154 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 9238 15802
rect 9290 15750 9302 15802
rect 9354 15750 9366 15802
rect 9418 15750 10856 15802
rect 1104 15728 10856 15750
rect 1854 15688 1860 15700
rect 1815 15660 1860 15688
rect 1854 15648 1860 15660
rect 1912 15648 1918 15700
rect 2222 15688 2228 15700
rect 2183 15660 2228 15688
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 3786 15688 3792 15700
rect 3747 15660 3792 15688
rect 3786 15648 3792 15660
rect 3844 15648 3850 15700
rect 9950 15688 9956 15700
rect 9911 15660 9956 15688
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 1946 15552 1952 15564
rect 1907 15524 1952 15552
rect 1946 15512 1952 15524
rect 2004 15512 2010 15564
rect 2222 15512 2228 15564
rect 2280 15552 2286 15564
rect 6178 15552 6184 15564
rect 2280 15524 6184 15552
rect 2280 15512 2286 15524
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 1857 15487 1915 15493
rect 1857 15484 1869 15487
rect 1820 15456 1869 15484
rect 1820 15444 1826 15456
rect 1857 15453 1869 15456
rect 1903 15453 1915 15487
rect 2866 15484 2872 15496
rect 2827 15456 2872 15484
rect 1857 15447 1915 15453
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 3970 15484 3976 15496
rect 3931 15456 3976 15484
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 4890 15444 4896 15496
rect 4948 15484 4954 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 4948 15456 10149 15484
rect 4948 15444 4954 15456
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 2314 15308 2320 15360
rect 2372 15348 2378 15360
rect 2685 15351 2743 15357
rect 2685 15348 2697 15351
rect 2372 15320 2697 15348
rect 2372 15308 2378 15320
rect 2685 15317 2697 15320
rect 2731 15317 2743 15351
rect 2685 15311 2743 15317
rect 1104 15258 10856 15280
rect 1104 15206 4214 15258
rect 4266 15206 4278 15258
rect 4330 15206 4342 15258
rect 4394 15206 4406 15258
rect 4458 15206 4470 15258
rect 4522 15206 7478 15258
rect 7530 15206 7542 15258
rect 7594 15206 7606 15258
rect 7658 15206 7670 15258
rect 7722 15206 7734 15258
rect 7786 15206 10856 15258
rect 1104 15184 10856 15206
rect 2130 15144 2136 15156
rect 2091 15116 2136 15144
rect 2130 15104 2136 15116
rect 2188 15104 2194 15156
rect 2961 15079 3019 15085
rect 2961 15045 2973 15079
rect 3007 15076 3019 15079
rect 3142 15076 3148 15088
rect 3007 15048 3148 15076
rect 3007 15045 3019 15048
rect 2961 15039 3019 15045
rect 3142 15036 3148 15048
rect 3200 15036 3206 15088
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 15008 2099 15011
rect 2406 15008 2412 15020
rect 2087 14980 2412 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 2406 14968 2412 14980
rect 2464 14968 2470 15020
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 15008 2835 15011
rect 3418 15008 3424 15020
rect 2823 14980 3424 15008
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 3418 14968 3424 14980
rect 3476 14968 3482 15020
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 15008 9919 15011
rect 9950 15008 9956 15020
rect 9907 14980 9956 15008
rect 9907 14977 9919 14980
rect 9861 14971 9919 14977
rect 9950 14968 9956 14980
rect 10008 14968 10014 15020
rect 10042 14872 10048 14884
rect 10003 14844 10048 14872
rect 10042 14832 10048 14844
rect 10100 14832 10106 14884
rect 2222 14764 2228 14816
rect 2280 14804 2286 14816
rect 4798 14804 4804 14816
rect 2280 14776 4804 14804
rect 2280 14764 2286 14776
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 1104 14714 10856 14736
rect 1104 14662 2582 14714
rect 2634 14662 2646 14714
rect 2698 14662 2710 14714
rect 2762 14662 2774 14714
rect 2826 14662 2838 14714
rect 2890 14662 5846 14714
rect 5898 14662 5910 14714
rect 5962 14662 5974 14714
rect 6026 14662 6038 14714
rect 6090 14662 6102 14714
rect 6154 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 9238 14714
rect 9290 14662 9302 14714
rect 9354 14662 9366 14714
rect 9418 14662 10856 14714
rect 1104 14640 10856 14662
rect 1670 14600 1676 14612
rect 1631 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 2777 14603 2835 14609
rect 2777 14600 2789 14603
rect 2004 14572 2789 14600
rect 2004 14560 2010 14572
rect 2777 14569 2789 14572
rect 2823 14569 2835 14603
rect 2958 14600 2964 14612
rect 2919 14572 2964 14600
rect 2777 14563 2835 14569
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14464 1639 14467
rect 2314 14464 2320 14476
rect 1627 14436 2320 14464
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 2314 14424 2320 14436
rect 2372 14424 2378 14476
rect 2792 14464 2820 14563
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 2866 14492 2872 14544
rect 2924 14532 2930 14544
rect 3789 14535 3847 14541
rect 3789 14532 3801 14535
rect 2924 14504 3801 14532
rect 2924 14492 2930 14504
rect 3789 14501 3801 14504
rect 3835 14501 3847 14535
rect 3789 14495 3847 14501
rect 4890 14464 4896 14476
rect 2792 14436 4896 14464
rect 4890 14424 4896 14436
rect 4948 14424 4954 14476
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 3786 14396 3792 14408
rect 1719 14368 3792 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 3970 14396 3976 14408
rect 3931 14368 3976 14396
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 9858 14396 9864 14408
rect 9819 14368 9864 14396
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 1397 14331 1455 14337
rect 1397 14297 1409 14331
rect 1443 14297 1455 14331
rect 1397 14291 1455 14297
rect 1412 14260 1440 14291
rect 2130 14288 2136 14340
rect 2188 14328 2194 14340
rect 2593 14331 2651 14337
rect 2593 14328 2605 14331
rect 2188 14300 2605 14328
rect 2188 14288 2194 14300
rect 2593 14297 2605 14300
rect 2639 14297 2651 14331
rect 2593 14291 2651 14297
rect 2809 14331 2867 14337
rect 2809 14297 2821 14331
rect 2855 14328 2867 14331
rect 3050 14328 3056 14340
rect 2855 14300 3056 14328
rect 2855 14297 2867 14300
rect 2809 14291 2867 14297
rect 3050 14288 3056 14300
rect 3108 14288 3114 14340
rect 2682 14260 2688 14272
rect 1412 14232 2688 14260
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 10042 14260 10048 14272
rect 10003 14232 10048 14260
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 1104 14170 10856 14192
rect 1104 14118 4214 14170
rect 4266 14118 4278 14170
rect 4330 14118 4342 14170
rect 4394 14118 4406 14170
rect 4458 14118 4470 14170
rect 4522 14118 7478 14170
rect 7530 14118 7542 14170
rect 7594 14118 7606 14170
rect 7658 14118 7670 14170
rect 7722 14118 7734 14170
rect 7786 14118 10856 14170
rect 1104 14096 10856 14118
rect 1397 14059 1455 14065
rect 1397 14025 1409 14059
rect 1443 14056 1455 14059
rect 1486 14056 1492 14068
rect 1443 14028 1492 14056
rect 1443 14025 1455 14028
rect 1397 14019 1455 14025
rect 1486 14016 1492 14028
rect 1544 14016 1550 14068
rect 1670 14016 1676 14068
rect 1728 14016 1734 14068
rect 2406 14056 2412 14068
rect 2367 14028 2412 14056
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 3053 14059 3111 14065
rect 3053 14025 3065 14059
rect 3099 14025 3111 14059
rect 3053 14019 3111 14025
rect 1688 13988 1716 14016
rect 3068 13988 3096 14019
rect 9582 14016 9588 14068
rect 9640 14056 9646 14068
rect 10045 14059 10103 14065
rect 10045 14056 10057 14059
rect 9640 14028 10057 14056
rect 9640 14016 9646 14028
rect 10045 14025 10057 14028
rect 10091 14025 10103 14059
rect 10045 14019 10103 14025
rect 1688 13960 3004 13988
rect 3068 13960 9904 13988
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13889 1639 13923
rect 2222 13920 2228 13932
rect 2183 13892 2228 13920
rect 1581 13883 1639 13889
rect 1596 13796 1624 13883
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13852 2099 13855
rect 2976 13852 3004 13960
rect 3234 13920 3240 13932
rect 3195 13892 3240 13920
rect 3234 13880 3240 13892
rect 3292 13920 3298 13932
rect 3510 13920 3516 13932
rect 3292 13892 3516 13920
rect 3292 13880 3298 13892
rect 3510 13880 3516 13892
rect 3568 13880 3574 13932
rect 3878 13920 3884 13932
rect 3839 13892 3884 13920
rect 3878 13880 3884 13892
rect 3936 13880 3942 13932
rect 9876 13929 9904 13960
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 2087 13824 2912 13852
rect 2976 13824 3740 13852
rect 2087 13821 2099 13824
rect 2041 13815 2099 13821
rect 1578 13744 1584 13796
rect 1636 13744 1642 13796
rect 2884 13784 2912 13824
rect 3602 13784 3608 13796
rect 2884 13756 3608 13784
rect 3602 13744 3608 13756
rect 3660 13744 3666 13796
rect 3712 13793 3740 13824
rect 3697 13787 3755 13793
rect 3697 13753 3709 13787
rect 3743 13753 3755 13787
rect 3697 13747 3755 13753
rect 1104 13626 10856 13648
rect 1104 13574 2582 13626
rect 2634 13574 2646 13626
rect 2698 13574 2710 13626
rect 2762 13574 2774 13626
rect 2826 13574 2838 13626
rect 2890 13574 5846 13626
rect 5898 13574 5910 13626
rect 5962 13574 5974 13626
rect 6026 13574 6038 13626
rect 6090 13574 6102 13626
rect 6154 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 9238 13626
rect 9290 13574 9302 13626
rect 9354 13574 9366 13626
rect 9418 13574 10856 13626
rect 1104 13552 10856 13574
rect 2406 13472 2412 13524
rect 2464 13512 2470 13524
rect 2464 13484 9536 13512
rect 2464 13472 2470 13484
rect 3786 13444 3792 13456
rect 3747 13416 3792 13444
rect 3786 13404 3792 13416
rect 3844 13404 3850 13456
rect 2314 13336 2320 13388
rect 2372 13376 2378 13388
rect 2866 13376 2872 13388
rect 2372 13348 2872 13376
rect 2372 13336 2378 13348
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 1302 13268 1308 13320
rect 1360 13308 1366 13320
rect 1581 13311 1639 13317
rect 1581 13308 1593 13311
rect 1360 13280 1593 13308
rect 1360 13268 1366 13280
rect 1581 13277 1593 13280
rect 1627 13277 1639 13311
rect 1581 13271 1639 13277
rect 2498 13268 2504 13320
rect 2556 13308 2562 13320
rect 2593 13311 2651 13317
rect 2593 13308 2605 13311
rect 2556 13280 2605 13308
rect 2556 13268 2562 13280
rect 2593 13277 2605 13280
rect 2639 13277 2651 13311
rect 3234 13308 3240 13320
rect 3195 13280 3240 13308
rect 2593 13271 2651 13277
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 3970 13308 3976 13320
rect 3931 13280 3976 13308
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 9508 13317 9536 13484
rect 9858 13472 9864 13524
rect 9916 13512 9922 13524
rect 9953 13515 10011 13521
rect 9953 13512 9965 13515
rect 9916 13484 9965 13512
rect 9916 13472 9922 13484
rect 9953 13481 9965 13484
rect 9999 13481 10011 13515
rect 9953 13475 10011 13481
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13277 9551 13311
rect 10134 13308 10140 13320
rect 10095 13280 10140 13308
rect 9493 13271 9551 13277
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 9858 13240 9864 13252
rect 2746 13212 9864 13240
rect 1394 13172 1400 13184
rect 1355 13144 1400 13172
rect 1394 13132 1400 13144
rect 1452 13132 1458 13184
rect 2409 13175 2467 13181
rect 2409 13141 2421 13175
rect 2455 13172 2467 13175
rect 2746 13172 2774 13212
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 2455 13144 2774 13172
rect 2455 13141 2467 13144
rect 2409 13135 2467 13141
rect 2958 13132 2964 13184
rect 3016 13172 3022 13184
rect 3053 13175 3111 13181
rect 3053 13172 3065 13175
rect 3016 13144 3065 13172
rect 3016 13132 3022 13144
rect 3053 13141 3065 13144
rect 3099 13141 3111 13175
rect 3053 13135 3111 13141
rect 9309 13175 9367 13181
rect 9309 13141 9321 13175
rect 9355 13172 9367 13175
rect 9674 13172 9680 13184
rect 9355 13144 9680 13172
rect 9355 13141 9367 13144
rect 9309 13135 9367 13141
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 1104 13082 10856 13104
rect 1104 13030 4214 13082
rect 4266 13030 4278 13082
rect 4330 13030 4342 13082
rect 4394 13030 4406 13082
rect 4458 13030 4470 13082
rect 4522 13030 7478 13082
rect 7530 13030 7542 13082
rect 7594 13030 7606 13082
rect 7658 13030 7670 13082
rect 7722 13030 7734 13082
rect 7786 13030 10856 13082
rect 1104 13008 10856 13030
rect 1397 12971 1455 12977
rect 1397 12937 1409 12971
rect 1443 12968 1455 12971
rect 2777 12971 2835 12977
rect 2777 12968 2789 12971
rect 1443 12940 2789 12968
rect 1443 12937 1455 12940
rect 1397 12931 1455 12937
rect 2777 12937 2789 12940
rect 2823 12968 2835 12971
rect 2961 12971 3019 12977
rect 2823 12940 2925 12968
rect 2823 12937 2835 12940
rect 2777 12931 2835 12937
rect 2884 12900 2912 12940
rect 2961 12937 2973 12971
rect 3007 12968 3019 12971
rect 3050 12968 3056 12980
rect 3007 12940 3056 12968
rect 3007 12937 3019 12940
rect 2961 12931 3019 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 9217 12971 9275 12977
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 9766 12968 9772 12980
rect 9263 12940 9772 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 2884 12872 9444 12900
rect 1210 12792 1216 12844
rect 1268 12832 1274 12844
rect 1581 12835 1639 12841
rect 1581 12832 1593 12835
rect 1268 12804 1593 12832
rect 1268 12792 1274 12804
rect 1581 12801 1593 12804
rect 1627 12801 1639 12835
rect 2590 12832 2596 12844
rect 2551 12804 2596 12832
rect 1581 12795 1639 12801
rect 2590 12792 2596 12804
rect 2648 12792 2654 12844
rect 9416 12841 9444 12872
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12832 2743 12835
rect 9401 12835 9459 12841
rect 2731 12804 2765 12832
rect 2731 12801 2743 12804
rect 2685 12795 2743 12801
rect 9401 12801 9413 12835
rect 9447 12801 9459 12835
rect 9858 12832 9864 12844
rect 9819 12804 9864 12832
rect 9401 12795 9459 12801
rect 1946 12724 1952 12776
rect 2004 12764 2010 12776
rect 2700 12764 2728 12795
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 10134 12764 10140 12776
rect 2004 12736 10140 12764
rect 2004 12724 2010 12736
rect 10134 12724 10140 12736
rect 10192 12724 10198 12776
rect 2406 12696 2412 12708
rect 2367 12668 2412 12696
rect 2406 12656 2412 12668
rect 2464 12656 2470 12708
rect 2590 12656 2596 12708
rect 2648 12656 2654 12708
rect 2866 12656 2872 12708
rect 2924 12696 2930 12708
rect 3050 12696 3056 12708
rect 2924 12668 3056 12696
rect 2924 12656 2930 12668
rect 3050 12656 3056 12668
rect 3108 12656 3114 12708
rect 2222 12588 2228 12640
rect 2280 12628 2286 12640
rect 2608 12628 2636 12656
rect 10042 12628 10048 12640
rect 2280 12600 2636 12628
rect 10003 12600 10048 12628
rect 2280 12588 2286 12600
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 1104 12538 10856 12560
rect 1104 12486 2582 12538
rect 2634 12486 2646 12538
rect 2698 12486 2710 12538
rect 2762 12486 2774 12538
rect 2826 12486 2838 12538
rect 2890 12486 5846 12538
rect 5898 12486 5910 12538
rect 5962 12486 5974 12538
rect 6026 12486 6038 12538
rect 6090 12486 6102 12538
rect 6154 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 9238 12538
rect 9290 12486 9302 12538
rect 9354 12486 9366 12538
rect 9418 12486 10856 12538
rect 1104 12464 10856 12486
rect 1394 12424 1400 12436
rect 1355 12396 1400 12424
rect 1394 12384 1400 12396
rect 1452 12384 1458 12436
rect 1762 12384 1768 12436
rect 1820 12424 1826 12436
rect 1857 12427 1915 12433
rect 1857 12424 1869 12427
rect 1820 12396 1869 12424
rect 1820 12384 1826 12396
rect 1857 12393 1869 12396
rect 1903 12393 1915 12427
rect 1857 12387 1915 12393
rect 2222 12384 2228 12436
rect 2280 12424 2286 12436
rect 9217 12427 9275 12433
rect 2280 12396 6132 12424
rect 2280 12384 2286 12396
rect 2958 12356 2964 12368
rect 1596 12328 2964 12356
rect 1596 12297 1624 12328
rect 2958 12316 2964 12328
rect 3016 12316 3022 12368
rect 3053 12359 3111 12365
rect 3053 12325 3065 12359
rect 3099 12325 3111 12359
rect 6104 12356 6132 12396
rect 9217 12393 9229 12427
rect 9263 12424 9275 12427
rect 9950 12424 9956 12436
rect 9263 12396 9956 12424
rect 9263 12393 9275 12396
rect 9217 12387 9275 12393
rect 9950 12384 9956 12396
rect 10008 12384 10014 12436
rect 6104 12328 9444 12356
rect 3053 12319 3111 12325
rect 1581 12291 1639 12297
rect 1581 12257 1593 12291
rect 1627 12257 1639 12291
rect 3068 12288 3096 12319
rect 1581 12251 1639 12257
rect 1688 12260 3096 12288
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12220 1455 12223
rect 1486 12220 1492 12232
rect 1443 12192 1492 12220
rect 1443 12189 1455 12192
rect 1397 12183 1455 12189
rect 1486 12180 1492 12192
rect 1544 12180 1550 12232
rect 1688 12229 1716 12260
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12189 1731 12223
rect 1673 12183 1731 12189
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 3234 12220 3240 12232
rect 2363 12192 2774 12220
rect 3195 12192 3240 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 2746 12152 2774 12192
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 9416 12229 9444 12328
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12189 9459 12223
rect 9858 12220 9864 12232
rect 9819 12192 9864 12220
rect 9401 12183 9459 12189
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 3602 12152 3608 12164
rect 2746 12124 3608 12152
rect 3602 12112 3608 12124
rect 3660 12112 3666 12164
rect 1118 12044 1124 12096
rect 1176 12084 1182 12096
rect 2501 12087 2559 12093
rect 2501 12084 2513 12087
rect 1176 12056 2513 12084
rect 1176 12044 1182 12056
rect 2501 12053 2513 12056
rect 2547 12053 2559 12087
rect 10042 12084 10048 12096
rect 10003 12056 10048 12084
rect 2501 12047 2559 12053
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 1104 11994 10856 12016
rect 1104 11942 4214 11994
rect 4266 11942 4278 11994
rect 4330 11942 4342 11994
rect 4394 11942 4406 11994
rect 4458 11942 4470 11994
rect 4522 11942 7478 11994
rect 7530 11942 7542 11994
rect 7594 11942 7606 11994
rect 7658 11942 7670 11994
rect 7722 11942 7734 11994
rect 7786 11942 10856 11994
rect 1104 11920 10856 11942
rect 2869 11883 2927 11889
rect 2869 11849 2881 11883
rect 2915 11880 2927 11883
rect 3142 11880 3148 11892
rect 2915 11852 3148 11880
rect 2915 11849 2927 11852
rect 2869 11843 2927 11849
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 9858 11880 9864 11892
rect 3467 11852 9864 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 1026 11704 1032 11756
rect 1084 11744 1090 11756
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1084 11716 1685 11744
rect 1084 11704 1090 11716
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 2685 11747 2743 11753
rect 2685 11744 2697 11747
rect 1673 11707 1731 11713
rect 2608 11716 2697 11744
rect 1302 11636 1308 11688
rect 1360 11676 1366 11688
rect 1397 11679 1455 11685
rect 1397 11676 1409 11679
rect 1360 11648 1409 11676
rect 1360 11636 1366 11648
rect 1397 11645 1409 11648
rect 1443 11645 1455 11679
rect 1397 11639 1455 11645
rect 2314 11568 2320 11620
rect 2372 11608 2378 11620
rect 2608 11608 2636 11716
rect 2685 11713 2697 11716
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 3605 11747 3663 11753
rect 3605 11744 3617 11747
rect 3384 11716 3617 11744
rect 3384 11704 3390 11716
rect 3605 11713 3617 11716
rect 3651 11713 3663 11747
rect 3605 11707 3663 11713
rect 2372 11580 2636 11608
rect 2372 11568 2378 11580
rect 1762 11500 1768 11552
rect 1820 11540 1826 11552
rect 2222 11540 2228 11552
rect 1820 11512 2228 11540
rect 1820 11500 1826 11512
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 1104 11450 10856 11472
rect 1104 11398 2582 11450
rect 2634 11398 2646 11450
rect 2698 11398 2710 11450
rect 2762 11398 2774 11450
rect 2826 11398 2838 11450
rect 2890 11398 5846 11450
rect 5898 11398 5910 11450
rect 5962 11398 5974 11450
rect 6026 11398 6038 11450
rect 6090 11398 6102 11450
rect 6154 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 9238 11450
rect 9290 11398 9302 11450
rect 9354 11398 9366 11450
rect 9418 11398 10856 11450
rect 1104 11376 10856 11398
rect 2038 11296 2044 11348
rect 2096 11336 2102 11348
rect 2222 11336 2228 11348
rect 2096 11308 2228 11336
rect 2096 11296 2102 11308
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 4798 11336 4804 11348
rect 2915 11308 4804 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 3789 11271 3847 11277
rect 3789 11237 3801 11271
rect 3835 11237 3847 11271
rect 10042 11268 10048 11280
rect 10003 11240 10048 11268
rect 3789 11231 3847 11237
rect 1670 11200 1676 11212
rect 1631 11172 1676 11200
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 2038 11160 2044 11212
rect 2096 11200 2102 11212
rect 3804 11200 3832 11231
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 2096 11172 3740 11200
rect 3804 11172 9904 11200
rect 2096 11160 2102 11172
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 3712 11132 3740 11172
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 2731 11104 3648 11132
rect 3712 11104 3985 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 3620 11064 3648 11104
rect 3973 11101 3985 11104
rect 4019 11132 4031 11135
rect 4706 11132 4712 11144
rect 4019 11104 4712 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 9876 11141 9904 11172
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11101 9919 11135
rect 9861 11095 9919 11101
rect 4062 11064 4068 11076
rect 3620 11036 4068 11064
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 1104 10906 10856 10928
rect 1104 10854 4214 10906
rect 4266 10854 4278 10906
rect 4330 10854 4342 10906
rect 4394 10854 4406 10906
rect 4458 10854 4470 10906
rect 4522 10854 7478 10906
rect 7530 10854 7542 10906
rect 7594 10854 7606 10906
rect 7658 10854 7670 10906
rect 7722 10854 7734 10906
rect 7786 10854 10856 10906
rect 1104 10832 10856 10854
rect 3421 10795 3479 10801
rect 3421 10761 3433 10795
rect 3467 10761 3479 10795
rect 3421 10755 3479 10761
rect 3436 10724 3464 10755
rect 3436 10696 9904 10724
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 3142 10656 3148 10668
rect 2731 10628 3148 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10656 3663 10659
rect 3970 10656 3976 10668
rect 3651 10628 3976 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 9876 10665 9904 10696
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 1302 10548 1308 10600
rect 1360 10588 1366 10600
rect 1397 10591 1455 10597
rect 1397 10588 1409 10591
rect 1360 10560 1409 10588
rect 1360 10548 1366 10560
rect 1397 10557 1409 10560
rect 1443 10557 1455 10591
rect 1397 10551 1455 10557
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 4614 10588 4620 10600
rect 1719 10560 4620 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 2869 10523 2927 10529
rect 2869 10489 2881 10523
rect 2915 10520 2927 10523
rect 5258 10520 5264 10532
rect 2915 10492 5264 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 1104 10362 10856 10384
rect 1104 10310 2582 10362
rect 2634 10310 2646 10362
rect 2698 10310 2710 10362
rect 2762 10310 2774 10362
rect 2826 10310 2838 10362
rect 2890 10310 5846 10362
rect 5898 10310 5910 10362
rect 5962 10310 5974 10362
rect 6026 10310 6038 10362
rect 6090 10310 6102 10362
rect 6154 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 9238 10362
rect 9290 10310 9302 10362
rect 9354 10310 9366 10362
rect 9418 10310 10856 10362
rect 1104 10288 10856 10310
rect 3053 10251 3111 10257
rect 3053 10217 3065 10251
rect 3099 10248 3111 10251
rect 3418 10248 3424 10260
rect 3099 10220 3424 10248
rect 3099 10217 3111 10220
rect 3053 10211 3111 10217
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 2130 10112 2136 10124
rect 1719 10084 2136 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 2130 10072 2136 10084
rect 2188 10072 2194 10124
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10044 2927 10047
rect 3050 10044 3056 10056
rect 2915 10016 3056 10044
rect 2915 10013 2927 10016
rect 2869 10007 2927 10013
rect 2792 9976 2820 10007
rect 3050 10004 3056 10016
rect 3108 10044 3114 10056
rect 3234 10044 3240 10056
rect 3108 10016 3240 10044
rect 3108 10004 3114 10016
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 3418 9976 3424 9988
rect 2792 9948 3424 9976
rect 3418 9936 3424 9948
rect 3476 9936 3482 9988
rect 1104 9818 10856 9840
rect 1104 9766 4214 9818
rect 4266 9766 4278 9818
rect 4330 9766 4342 9818
rect 4394 9766 4406 9818
rect 4458 9766 4470 9818
rect 4522 9766 7478 9818
rect 7530 9766 7542 9818
rect 7594 9766 7606 9818
rect 7658 9766 7670 9818
rect 7722 9766 7734 9818
rect 7786 9766 10856 9818
rect 1104 9744 10856 9766
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 1854 9568 1860 9580
rect 1719 9540 1860 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 1854 9528 1860 9540
rect 1912 9528 1918 9580
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9568 2743 9571
rect 3050 9568 3056 9580
rect 2731 9540 3056 9568
rect 2731 9537 2743 9540
rect 2685 9531 2743 9537
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 3602 9568 3608 9580
rect 3563 9540 3608 9568
rect 3602 9528 3608 9540
rect 3660 9528 3666 9580
rect 3694 9528 3700 9580
rect 3752 9568 3758 9580
rect 9861 9571 9919 9577
rect 9861 9568 9873 9571
rect 3752 9540 9873 9568
rect 3752 9528 3758 9540
rect 9861 9537 9873 9540
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 2866 9432 2872 9444
rect 2827 9404 2872 9432
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 10042 9432 10048 9444
rect 10003 9404 10048 9432
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 3421 9367 3479 9373
rect 3421 9333 3433 9367
rect 3467 9364 3479 9367
rect 9858 9364 9864 9376
rect 3467 9336 9864 9364
rect 3467 9333 3479 9336
rect 3421 9327 3479 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 1104 9274 10856 9296
rect 1104 9222 2582 9274
rect 2634 9222 2646 9274
rect 2698 9222 2710 9274
rect 2762 9222 2774 9274
rect 2826 9222 2838 9274
rect 2890 9222 5846 9274
rect 5898 9222 5910 9274
rect 5962 9222 5974 9274
rect 6026 9222 6038 9274
rect 6090 9222 6102 9274
rect 6154 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 9238 9274
rect 9290 9222 9302 9274
rect 9354 9222 9366 9274
rect 9418 9222 10856 9274
rect 1104 9200 10856 9222
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 2958 9160 2964 9172
rect 2915 9132 2964 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 9024 1731 9027
rect 2406 9024 2412 9036
rect 1719 8996 2412 9024
rect 1719 8993 1731 8996
rect 1673 8987 1731 8993
rect 2406 8984 2412 8996
rect 2464 8984 2470 9036
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 3050 8956 3056 8968
rect 2731 8928 3056 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 3142 8916 3148 8968
rect 3200 8956 3206 8968
rect 3970 8956 3976 8968
rect 3200 8928 3976 8956
rect 3200 8916 3206 8928
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 9858 8956 9864 8968
rect 9819 8928 9864 8956
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8820 3847 8823
rect 9858 8820 9864 8832
rect 3835 8792 9864 8820
rect 3835 8789 3847 8792
rect 3789 8783 3847 8789
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 10042 8820 10048 8832
rect 10003 8792 10048 8820
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 1104 8730 10856 8752
rect 1104 8678 4214 8730
rect 4266 8678 4278 8730
rect 4330 8678 4342 8730
rect 4394 8678 4406 8730
rect 4458 8678 4470 8730
rect 4522 8678 7478 8730
rect 7530 8678 7542 8730
rect 7594 8678 7606 8730
rect 7658 8678 7670 8730
rect 7722 8678 7734 8730
rect 7786 8678 10856 8730
rect 1104 8656 10856 8678
rect 3050 8616 3056 8628
rect 3011 8588 3056 8616
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 3513 8619 3571 8625
rect 3513 8585 3525 8619
rect 3559 8616 3571 8619
rect 3694 8616 3700 8628
rect 3559 8588 3700 8616
rect 3559 8585 3571 8588
rect 3513 8579 3571 8585
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 1578 8508 1584 8560
rect 1636 8548 1642 8560
rect 1636 8520 3740 8548
rect 1636 8508 1642 8520
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 1762 8480 1768 8492
rect 1719 8452 1768 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 1762 8440 1768 8452
rect 1820 8440 1826 8492
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8480 2927 8483
rect 3234 8480 3240 8492
rect 2915 8452 3240 8480
rect 2915 8449 2927 8452
rect 2869 8443 2927 8449
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 3712 8489 3740 8520
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8449 3755 8483
rect 9858 8480 9864 8492
rect 9819 8452 9864 8480
rect 3697 8443 3755 8449
rect 9858 8440 9864 8452
rect 9916 8440 9922 8492
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 2406 8372 2412 8424
rect 2464 8412 2470 8424
rect 2685 8415 2743 8421
rect 2685 8412 2697 8415
rect 2464 8384 2697 8412
rect 2464 8372 2470 8384
rect 2685 8381 2697 8384
rect 2731 8381 2743 8415
rect 2685 8375 2743 8381
rect 10042 8344 10048 8356
rect 10003 8316 10048 8344
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 1104 8186 10856 8208
rect 1104 8134 2582 8186
rect 2634 8134 2646 8186
rect 2698 8134 2710 8186
rect 2762 8134 2774 8186
rect 2826 8134 2838 8186
rect 2890 8134 5846 8186
rect 5898 8134 5910 8186
rect 5962 8134 5974 8186
rect 6026 8134 6038 8186
rect 6090 8134 6102 8186
rect 6154 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 9238 8186
rect 9290 8134 9302 8186
rect 9354 8134 9366 8186
rect 9418 8134 10856 8186
rect 1104 8112 10856 8134
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 1946 7936 1952 7948
rect 1719 7908 1952 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7868 2927 7871
rect 3050 7868 3056 7880
rect 2915 7840 3056 7868
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 2685 7735 2743 7741
rect 2685 7701 2697 7735
rect 2731 7732 2743 7735
rect 9858 7732 9864 7744
rect 2731 7704 9864 7732
rect 2731 7701 2743 7704
rect 2685 7695 2743 7701
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 1104 7642 10856 7664
rect 1104 7590 4214 7642
rect 4266 7590 4278 7642
rect 4330 7590 4342 7642
rect 4394 7590 4406 7642
rect 4458 7590 4470 7642
rect 4522 7590 7478 7642
rect 7530 7590 7542 7642
rect 7594 7590 7606 7642
rect 7658 7590 7670 7642
rect 7722 7590 7734 7642
rect 7786 7590 10856 7642
rect 1104 7568 10856 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 3510 7528 3516 7540
rect 1627 7500 3516 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 2409 7463 2467 7469
rect 2409 7429 2421 7463
rect 2455 7460 2467 7463
rect 2498 7460 2504 7472
rect 2455 7432 2504 7460
rect 2455 7429 2467 7432
rect 2409 7423 2467 7429
rect 2498 7420 2504 7432
rect 2556 7420 2562 7472
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 2222 7392 2228 7404
rect 2183 7364 2228 7392
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 4062 7392 4068 7404
rect 4023 7364 4068 7392
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 9876 7324 9904 7355
rect 3896 7296 9904 7324
rect 3896 7265 3924 7296
rect 3881 7259 3939 7265
rect 3881 7225 3893 7259
rect 3927 7225 3939 7259
rect 3881 7219 3939 7225
rect 10042 7188 10048 7200
rect 10003 7160 10048 7188
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 1104 7098 10856 7120
rect 1104 7046 2582 7098
rect 2634 7046 2646 7098
rect 2698 7046 2710 7098
rect 2762 7046 2774 7098
rect 2826 7046 2838 7098
rect 2890 7046 5846 7098
rect 5898 7046 5910 7098
rect 5962 7046 5974 7098
rect 6026 7046 6038 7098
rect 6090 7046 6102 7098
rect 6154 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 9238 7098
rect 9290 7046 9302 7098
rect 9354 7046 9366 7098
rect 9418 7046 10856 7098
rect 1104 7024 10856 7046
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 3326 6848 3332 6860
rect 2455 6820 3332 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 3326 6808 3332 6820
rect 3384 6808 3390 6860
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6780 1455 6783
rect 1670 6780 1676 6792
rect 1443 6752 1676 6780
rect 1443 6749 1455 6752
rect 1397 6743 1455 6749
rect 1670 6740 1676 6752
rect 1728 6780 1734 6792
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 1728 6752 3065 6780
rect 1728 6740 1734 6752
rect 3053 6749 3065 6752
rect 3099 6749 3111 6783
rect 9858 6780 9864 6792
rect 9819 6752 9864 6780
rect 3053 6743 3111 6749
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 2222 6712 2228 6724
rect 2183 6684 2228 6712
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 9858 6644 9864 6656
rect 2915 6616 9864 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 10042 6644 10048 6656
rect 10003 6616 10048 6644
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 1104 6554 10856 6576
rect 1104 6502 4214 6554
rect 4266 6502 4278 6554
rect 4330 6502 4342 6554
rect 4394 6502 4406 6554
rect 4458 6502 4470 6554
rect 4522 6502 7478 6554
rect 7530 6502 7542 6554
rect 7594 6502 7606 6554
rect 7658 6502 7670 6554
rect 7722 6502 7734 6554
rect 7786 6502 10856 6554
rect 1104 6480 10856 6502
rect 2501 6443 2559 6449
rect 2501 6409 2513 6443
rect 2547 6440 2559 6443
rect 3970 6440 3976 6452
rect 2547 6412 3976 6440
rect 2547 6409 2559 6412
rect 2501 6403 2559 6409
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 2038 6372 2044 6384
rect 1999 6344 2044 6372
rect 2038 6332 2044 6344
rect 2096 6332 2102 6384
rect 1854 6304 1860 6316
rect 1815 6276 1860 6304
rect 1854 6264 1860 6276
rect 1912 6264 1918 6316
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 2958 6304 2964 6316
rect 2731 6276 2964 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3326 6304 3332 6316
rect 3287 6276 3332 6304
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 3145 6171 3203 6177
rect 3145 6137 3157 6171
rect 3191 6168 3203 6171
rect 3602 6168 3608 6180
rect 3191 6140 3608 6168
rect 3191 6137 3203 6140
rect 3145 6131 3203 6137
rect 3602 6128 3608 6140
rect 3660 6128 3666 6180
rect 1104 6010 10856 6032
rect 1104 5958 2582 6010
rect 2634 5958 2646 6010
rect 2698 5958 2710 6010
rect 2762 5958 2774 6010
rect 2826 5958 2838 6010
rect 2890 5958 5846 6010
rect 5898 5958 5910 6010
rect 5962 5958 5974 6010
rect 6026 5958 6038 6010
rect 6090 5958 6102 6010
rect 6154 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 9238 6010
rect 9290 5958 9302 6010
rect 9354 5958 9366 6010
rect 9418 5958 10856 6010
rect 1104 5936 10856 5958
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 3053 5899 3111 5905
rect 3053 5896 3065 5899
rect 2372 5868 3065 5896
rect 2372 5856 2378 5868
rect 3053 5865 3065 5868
rect 3099 5865 3111 5899
rect 3053 5859 3111 5865
rect 1486 5720 1492 5772
rect 1544 5760 1550 5772
rect 1673 5763 1731 5769
rect 1673 5760 1685 5763
rect 1544 5732 1685 5760
rect 1544 5720 1550 5732
rect 1673 5729 1685 5732
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 3418 5720 3424 5772
rect 3476 5760 3482 5772
rect 3789 5763 3847 5769
rect 3789 5760 3801 5763
rect 3476 5732 3801 5760
rect 3476 5720 3482 5732
rect 3789 5729 3801 5732
rect 3835 5729 3847 5763
rect 3789 5723 3847 5729
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 3234 5692 3240 5704
rect 2915 5664 3240 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 2792 5624 2820 5655
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 3878 5652 3884 5704
rect 3936 5692 3942 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3936 5664 3985 5692
rect 3936 5652 3942 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 9858 5692 9864 5704
rect 9819 5664 9864 5692
rect 3973 5655 4031 5661
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 3602 5624 3608 5636
rect 2792 5596 3608 5624
rect 3602 5584 3608 5596
rect 3660 5584 3666 5636
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5556 4215 5559
rect 6822 5556 6828 5568
rect 4203 5528 6828 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 10042 5556 10048 5568
rect 10003 5528 10048 5556
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 1104 5466 10856 5488
rect 1104 5414 4214 5466
rect 4266 5414 4278 5466
rect 4330 5414 4342 5466
rect 4394 5414 4406 5466
rect 4458 5414 4470 5466
rect 4522 5414 7478 5466
rect 7530 5414 7542 5466
rect 7594 5414 7606 5466
rect 7658 5414 7670 5466
rect 7722 5414 7734 5466
rect 7786 5414 10856 5466
rect 1104 5392 10856 5414
rect 3510 5352 3516 5364
rect 2746 5324 3516 5352
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 1360 5188 1409 5216
rect 1360 5176 1366 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 2746 5216 2774 5324
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 3694 5352 3700 5364
rect 3655 5324 3700 5352
rect 3694 5312 3700 5324
rect 3752 5312 3758 5364
rect 9217 5355 9275 5361
rect 9217 5321 9229 5355
rect 9263 5321 9275 5355
rect 9217 5315 9275 5321
rect 3142 5284 3148 5296
rect 2884 5256 3148 5284
rect 2884 5225 2912 5256
rect 3142 5244 3148 5256
rect 3200 5284 3206 5296
rect 3878 5284 3884 5296
rect 3200 5256 3884 5284
rect 3200 5244 3206 5256
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 9232 5284 9260 5315
rect 9232 5256 9904 5284
rect 1719 5188 2774 5216
rect 2869 5219 2927 5225
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 2869 5185 2881 5219
rect 2915 5185 2927 5219
rect 3510 5216 3516 5228
rect 3471 5188 3516 5216
rect 2869 5179 2927 5185
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 6822 5176 6828 5228
rect 6880 5216 6886 5228
rect 9876 5225 9904 5256
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 6880 5188 9413 5216
rect 6880 5176 6886 5188
rect 9401 5185 9413 5188
rect 9447 5185 9459 5219
rect 9401 5179 9459 5185
rect 9861 5219 9919 5225
rect 9861 5185 9873 5219
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 2222 5108 2228 5160
rect 2280 5148 2286 5160
rect 2406 5148 2412 5160
rect 2280 5120 2412 5148
rect 2280 5108 2286 5120
rect 2406 5108 2412 5120
rect 2464 5148 2470 5160
rect 2685 5151 2743 5157
rect 2685 5148 2697 5151
rect 2464 5120 2697 5148
rect 2464 5108 2470 5120
rect 2685 5117 2697 5120
rect 2731 5117 2743 5151
rect 2685 5111 2743 5117
rect 3053 5083 3111 5089
rect 3053 5049 3065 5083
rect 3099 5080 3111 5083
rect 5166 5080 5172 5092
rect 3099 5052 5172 5080
rect 3099 5049 3111 5052
rect 3053 5043 3111 5049
rect 5166 5040 5172 5052
rect 5224 5040 5230 5092
rect 10042 5012 10048 5024
rect 10003 4984 10048 5012
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 1104 4922 10856 4944
rect 1104 4870 2582 4922
rect 2634 4870 2646 4922
rect 2698 4870 2710 4922
rect 2762 4870 2774 4922
rect 2826 4870 2838 4922
rect 2890 4870 5846 4922
rect 5898 4870 5910 4922
rect 5962 4870 5974 4922
rect 6026 4870 6038 4922
rect 6090 4870 6102 4922
rect 6154 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 9238 4922
rect 9290 4870 9302 4922
rect 9354 4870 9366 4922
rect 9418 4870 10856 4922
rect 1104 4848 10856 4870
rect 3970 4808 3976 4820
rect 3931 4780 3976 4808
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 3234 4740 3240 4752
rect 1872 4712 3240 4740
rect 1762 4604 1768 4616
rect 1723 4576 1768 4604
rect 1762 4564 1768 4576
rect 1820 4564 1826 4616
rect 1872 4613 1900 4712
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 2041 4675 2099 4681
rect 2041 4641 2053 4675
rect 2087 4672 2099 4675
rect 2087 4644 3832 4672
rect 2087 4641 2099 4644
rect 2041 4635 2099 4641
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4604 1915 4607
rect 1946 4604 1952 4616
rect 1903 4576 1952 4604
rect 1903 4573 1915 4576
rect 1857 4567 1915 4573
rect 1946 4564 1952 4576
rect 2004 4564 2010 4616
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4604 3019 4607
rect 3234 4604 3240 4616
rect 3007 4576 3240 4604
rect 3007 4573 3019 4576
rect 2961 4567 3019 4573
rect 2884 4536 2912 4567
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 3804 4613 3832 4644
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4573 3847 4607
rect 4706 4604 4712 4616
rect 4667 4576 4712 4604
rect 3789 4567 3847 4573
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 9858 4604 9864 4616
rect 9819 4576 9864 4604
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 3145 4539 3203 4545
rect 2884 4508 3004 4536
rect 2976 4468 3004 4508
rect 3145 4505 3157 4539
rect 3191 4536 3203 4539
rect 4614 4536 4620 4548
rect 3191 4508 4620 4536
rect 3191 4505 3203 4508
rect 3145 4499 3203 4505
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 3326 4468 3332 4480
rect 2976 4440 3332 4468
rect 3326 4428 3332 4440
rect 3384 4468 3390 4480
rect 3786 4468 3792 4480
rect 3384 4440 3792 4468
rect 3384 4428 3390 4440
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 4525 4471 4583 4477
rect 4525 4437 4537 4471
rect 4571 4468 4583 4471
rect 9766 4468 9772 4480
rect 4571 4440 9772 4468
rect 4571 4437 4583 4440
rect 4525 4431 4583 4437
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 10042 4468 10048 4480
rect 10003 4440 10048 4468
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 1104 4378 10856 4400
rect 1104 4326 4214 4378
rect 4266 4326 4278 4378
rect 4330 4326 4342 4378
rect 4394 4326 4406 4378
rect 4458 4326 4470 4378
rect 4522 4326 7478 4378
rect 7530 4326 7542 4378
rect 7594 4326 7606 4378
rect 7658 4326 7670 4378
rect 7722 4326 7734 4378
rect 7786 4326 10856 4378
rect 1104 4304 10856 4326
rect 9858 4224 9864 4276
rect 9916 4264 9922 4276
rect 9953 4267 10011 4273
rect 9953 4264 9965 4267
rect 9916 4236 9965 4264
rect 9916 4224 9922 4236
rect 9953 4233 9965 4236
rect 9999 4233 10011 4267
rect 9953 4227 10011 4233
rect 2792 4168 4108 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 2792 4128 2820 4168
rect 4080 4140 4108 4168
rect 1719 4100 2820 4128
rect 2869 4131 2927 4137
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3142 4128 3148 4140
rect 2915 4100 3148 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3142 4088 3148 4100
rect 3200 4128 3206 4140
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 3200 4100 3709 4128
rect 3200 4088 3206 4100
rect 3697 4097 3709 4100
rect 3743 4128 3755 4131
rect 3970 4128 3976 4140
rect 3743 4100 3976 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4062 4088 4068 4140
rect 4120 4088 4126 4140
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 4614 4128 4620 4140
rect 4571 4100 4620 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 5166 4128 5172 4140
rect 5127 4100 5172 4128
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 10134 4128 10140 4140
rect 10095 4100 10140 4128
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 1394 4060 1400 4072
rect 1355 4032 1400 4060
rect 1394 4020 1400 4032
rect 1452 4020 1458 4072
rect 1762 4020 1768 4072
rect 1820 4060 1826 4072
rect 2406 4060 2412 4072
rect 1820 4032 2412 4060
rect 1820 4020 1826 4032
rect 2406 4020 2412 4032
rect 2464 4060 2470 4072
rect 2685 4063 2743 4069
rect 2685 4060 2697 4063
rect 2464 4032 2697 4060
rect 2464 4020 2470 4032
rect 2685 4029 2697 4032
rect 2731 4029 2743 4063
rect 2685 4023 2743 4029
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4029 3571 4063
rect 3513 4023 3571 4029
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4060 3939 4063
rect 4706 4060 4712 4072
rect 3927 4032 4712 4060
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 3528 3992 3556 4023
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 4154 3992 4160 4004
rect 3528 3964 4160 3992
rect 4154 3952 4160 3964
rect 4212 3952 4218 4004
rect 4341 3995 4399 4001
rect 4341 3961 4353 3995
rect 4387 3992 4399 3995
rect 5626 3992 5632 4004
rect 4387 3964 5632 3992
rect 4387 3961 4399 3964
rect 4341 3955 4399 3961
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 3053 3927 3111 3933
rect 3053 3893 3065 3927
rect 3099 3924 3111 3927
rect 3786 3924 3792 3936
rect 3099 3896 3792 3924
rect 3099 3893 3111 3896
rect 3053 3887 3111 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3924 5043 3927
rect 9030 3924 9036 3936
rect 5031 3896 9036 3924
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 1104 3834 10856 3856
rect 1104 3782 2582 3834
rect 2634 3782 2646 3834
rect 2698 3782 2710 3834
rect 2762 3782 2774 3834
rect 2826 3782 2838 3834
rect 2890 3782 5846 3834
rect 5898 3782 5910 3834
rect 5962 3782 5974 3834
rect 6026 3782 6038 3834
rect 6090 3782 6102 3834
rect 6154 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 9238 3834
rect 9290 3782 9302 3834
rect 9354 3782 9366 3834
rect 9418 3782 10856 3834
rect 1104 3760 10856 3782
rect 2225 3723 2283 3729
rect 2225 3689 2237 3723
rect 2271 3720 2283 3723
rect 3510 3720 3516 3732
rect 2271 3692 3516 3720
rect 2271 3689 2283 3692
rect 2225 3683 2283 3689
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 4157 3723 4215 3729
rect 4157 3689 4169 3723
rect 4203 3720 4215 3723
rect 10134 3720 10140 3732
rect 4203 3692 10140 3720
rect 4203 3689 4215 3692
rect 4157 3683 4215 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 4154 3584 4160 3596
rect 1903 3556 4160 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 4154 3544 4160 3556
rect 4212 3584 4218 3596
rect 4614 3584 4620 3596
rect 4212 3556 4620 3584
rect 4212 3544 4218 3556
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 1946 3476 1952 3528
rect 2004 3516 2010 3528
rect 2041 3519 2099 3525
rect 2041 3516 2053 3519
rect 2004 3488 2053 3516
rect 2004 3476 2010 3488
rect 2041 3485 2053 3488
rect 2087 3485 2099 3519
rect 2041 3479 2099 3485
rect 2498 3476 2504 3528
rect 2556 3516 2562 3528
rect 2869 3519 2927 3525
rect 2869 3516 2881 3519
rect 2556 3488 2881 3516
rect 2556 3476 2562 3488
rect 2869 3485 2881 3488
rect 2915 3485 2927 3519
rect 2869 3479 2927 3485
rect 3602 3476 3608 3528
rect 3660 3516 3666 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3660 3488 3801 3516
rect 3660 3476 3666 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3970 3516 3976 3528
rect 3931 3488 3976 3516
rect 3789 3479 3847 3485
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9824 3488 9873 3516
rect 9824 3476 9830 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 2682 3380 2688 3392
rect 2643 3352 2688 3380
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 10042 3380 10048 3392
rect 10003 3352 10048 3380
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 1104 3290 10856 3312
rect 1104 3238 4214 3290
rect 4266 3238 4278 3290
rect 4330 3238 4342 3290
rect 4394 3238 4406 3290
rect 4458 3238 4470 3290
rect 4522 3238 7478 3290
rect 7530 3238 7542 3290
rect 7594 3238 7606 3290
rect 7658 3238 7670 3290
rect 7722 3238 7734 3290
rect 7786 3238 10856 3290
rect 1104 3216 10856 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 2130 3176 2136 3188
rect 1627 3148 2136 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 2130 3136 2136 3148
rect 2188 3136 2194 3188
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 3050 3176 3056 3188
rect 2823 3148 3056 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 3602 3136 3608 3188
rect 3660 3176 3666 3188
rect 4249 3179 4307 3185
rect 4249 3176 4261 3179
rect 3660 3148 4261 3176
rect 3660 3136 3666 3148
rect 4249 3145 4261 3148
rect 4295 3145 4307 3179
rect 4249 3139 4307 3145
rect 2682 3068 2688 3120
rect 2740 3108 2746 3120
rect 9674 3108 9680 3120
rect 2740 3080 9680 3108
rect 2740 3068 2746 3080
rect 9674 3068 9680 3080
rect 9732 3068 9738 3120
rect 1397 3043 1455 3049
rect 1397 3009 1409 3043
rect 1443 3009 1455 3043
rect 2314 3040 2320 3052
rect 2275 3012 2320 3040
rect 1397 3003 1455 3009
rect 1412 2972 1440 3003
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 2958 3040 2964 3052
rect 2919 3012 2964 3040
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 3786 3040 3792 3052
rect 3747 3012 3792 3040
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 4430 3040 4436 3052
rect 4391 3012 4436 3040
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 2498 2972 2504 2984
rect 1412 2944 2504 2972
rect 2498 2932 2504 2944
rect 2556 2932 2562 2984
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 5092 2972 5120 3003
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 9125 3043 9183 3049
rect 9125 3040 9137 3043
rect 9088 3012 9137 3040
rect 9088 3000 9094 3012
rect 9125 3009 9137 3012
rect 9171 3009 9183 3043
rect 9125 3003 9183 3009
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 4212 2944 5120 2972
rect 4212 2932 4218 2944
rect 1670 2864 1676 2916
rect 1728 2904 1734 2916
rect 2133 2907 2191 2913
rect 2133 2904 2145 2907
rect 1728 2876 2145 2904
rect 1728 2864 1734 2876
rect 2133 2873 2145 2876
rect 2179 2873 2191 2907
rect 2133 2867 2191 2873
rect 3605 2907 3663 2913
rect 3605 2873 3617 2907
rect 3651 2904 3663 2907
rect 9876 2904 9904 3003
rect 3651 2876 9904 2904
rect 3651 2873 3663 2876
rect 3605 2867 3663 2873
rect 3418 2796 3424 2848
rect 3476 2836 3482 2848
rect 4893 2839 4951 2845
rect 4893 2836 4905 2839
rect 3476 2808 4905 2836
rect 3476 2796 3482 2808
rect 4893 2805 4905 2808
rect 4939 2805 4951 2839
rect 4893 2799 4951 2805
rect 9309 2839 9367 2845
rect 9309 2805 9321 2839
rect 9355 2836 9367 2839
rect 9490 2836 9496 2848
rect 9355 2808 9496 2836
rect 9355 2805 9367 2808
rect 9309 2799 9367 2805
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 10042 2836 10048 2848
rect 10003 2808 10048 2836
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 1104 2746 10856 2768
rect 1104 2694 2582 2746
rect 2634 2694 2646 2746
rect 2698 2694 2710 2746
rect 2762 2694 2774 2746
rect 2826 2694 2838 2746
rect 2890 2694 5846 2746
rect 5898 2694 5910 2746
rect 5962 2694 5974 2746
rect 6026 2694 6038 2746
rect 6090 2694 6102 2746
rect 6154 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 9238 2746
rect 9290 2694 9302 2746
rect 9354 2694 9366 2746
rect 9418 2694 10856 2746
rect 1104 2672 10856 2694
rect 2498 2592 2504 2644
rect 2556 2632 2562 2644
rect 2685 2635 2743 2641
rect 2685 2632 2697 2635
rect 2556 2604 2697 2632
rect 2556 2592 2562 2604
rect 2685 2601 2697 2604
rect 2731 2601 2743 2635
rect 2685 2595 2743 2601
rect 4433 2635 4491 2641
rect 4433 2601 4445 2635
rect 4479 2632 4491 2635
rect 4614 2632 4620 2644
rect 4479 2604 4620 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 2406 2524 2412 2576
rect 2464 2564 2470 2576
rect 3789 2567 3847 2573
rect 3789 2564 3801 2567
rect 2464 2536 3801 2564
rect 2464 2524 2470 2536
rect 3789 2533 3801 2536
rect 3835 2533 3847 2567
rect 3789 2527 3847 2533
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 4430 2496 4436 2508
rect 2832 2468 4436 2496
rect 2832 2456 2838 2468
rect 4430 2456 4436 2468
rect 4488 2456 4494 2508
rect 1394 2428 1400 2440
rect 1355 2400 1400 2428
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2397 1731 2431
rect 2866 2428 2872 2440
rect 2827 2400 2872 2428
rect 1673 2391 1731 2397
rect 1688 2360 1716 2391
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3970 2428 3976 2440
rect 3931 2400 3976 2428
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4120 2400 4629 2428
rect 4120 2388 4126 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 5258 2428 5264 2440
rect 5219 2400 5264 2428
rect 4617 2391 4675 2397
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 5684 2400 9137 2428
rect 5684 2388 5690 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9732 2400 9873 2428
rect 9732 2388 9738 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 3326 2360 3332 2372
rect 1688 2332 3332 2360
rect 3326 2320 3332 2332
rect 3384 2320 3390 2372
rect 2222 2252 2228 2304
rect 2280 2292 2286 2304
rect 5077 2295 5135 2301
rect 5077 2292 5089 2295
rect 2280 2264 5089 2292
rect 2280 2252 2286 2264
rect 5077 2261 5089 2264
rect 5123 2261 5135 2295
rect 9306 2292 9312 2304
rect 9267 2264 9312 2292
rect 5077 2255 5135 2261
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 9582 2252 9588 2304
rect 9640 2292 9646 2304
rect 10045 2295 10103 2301
rect 10045 2292 10057 2295
rect 9640 2264 10057 2292
rect 9640 2252 9646 2264
rect 10045 2261 10057 2264
rect 10091 2261 10103 2295
rect 10045 2255 10103 2261
rect 1104 2202 10856 2224
rect 1104 2150 4214 2202
rect 4266 2150 4278 2202
rect 4330 2150 4342 2202
rect 4394 2150 4406 2202
rect 4458 2150 4470 2202
rect 4522 2150 7478 2202
rect 7530 2150 7542 2202
rect 7594 2150 7606 2202
rect 7658 2150 7670 2202
rect 7722 2150 7734 2202
rect 7786 2150 10856 2202
rect 1104 2128 10856 2150
rect 2774 1028 2780 1080
rect 2832 1068 2838 1080
rect 5258 1068 5264 1080
rect 2832 1040 5264 1068
rect 2832 1028 2838 1040
rect 5258 1028 5264 1040
rect 5316 1028 5322 1080
<< via1 >>
rect 2582 77766 2634 77818
rect 2646 77766 2698 77818
rect 2710 77766 2762 77818
rect 2774 77766 2826 77818
rect 2838 77766 2890 77818
rect 5846 77766 5898 77818
rect 5910 77766 5962 77818
rect 5974 77766 6026 77818
rect 6038 77766 6090 77818
rect 6102 77766 6154 77818
rect 9110 77766 9162 77818
rect 9174 77766 9226 77818
rect 9238 77766 9290 77818
rect 9302 77766 9354 77818
rect 9366 77766 9418 77818
rect 3516 77664 3568 77716
rect 1400 77503 1452 77512
rect 1400 77469 1409 77503
rect 1409 77469 1443 77503
rect 1443 77469 1452 77503
rect 1400 77460 1452 77469
rect 2964 77596 3016 77648
rect 2964 77503 3016 77512
rect 2964 77469 2973 77503
rect 2973 77469 3007 77503
rect 3007 77469 3016 77503
rect 2964 77460 3016 77469
rect 3976 77503 4028 77512
rect 3976 77469 3985 77503
rect 3985 77469 4019 77503
rect 4019 77469 4028 77503
rect 3976 77460 4028 77469
rect 4068 77460 4120 77512
rect 9404 77503 9456 77512
rect 9404 77469 9413 77503
rect 9413 77469 9447 77503
rect 9447 77469 9456 77503
rect 9404 77460 9456 77469
rect 9956 77503 10008 77512
rect 9956 77469 9965 77503
rect 9965 77469 9999 77503
rect 9999 77469 10008 77503
rect 9956 77460 10008 77469
rect 7840 77392 7892 77444
rect 2044 77324 2096 77376
rect 2872 77324 2924 77376
rect 3148 77324 3200 77376
rect 3884 77324 3936 77376
rect 8300 77324 8352 77376
rect 4214 77222 4266 77274
rect 4278 77222 4330 77274
rect 4342 77222 4394 77274
rect 4406 77222 4458 77274
rect 4470 77222 4522 77274
rect 7478 77222 7530 77274
rect 7542 77222 7594 77274
rect 7606 77222 7658 77274
rect 7670 77222 7722 77274
rect 7734 77222 7786 77274
rect 3700 77052 3752 77104
rect 1492 76984 1544 77036
rect 2320 76984 2372 77036
rect 2504 76984 2556 77036
rect 3332 77027 3384 77036
rect 3332 76993 3341 77027
rect 3341 76993 3375 77027
rect 3375 76993 3384 77027
rect 3332 76984 3384 76993
rect 3424 76984 3476 77036
rect 9496 76984 9548 77036
rect 9588 76984 9640 77036
rect 3056 76916 3108 76968
rect 3608 76916 3660 76968
rect 1952 76823 2004 76832
rect 1952 76789 1961 76823
rect 1961 76789 1995 76823
rect 1995 76789 2004 76823
rect 1952 76780 2004 76789
rect 2412 76780 2464 76832
rect 3056 76780 3108 76832
rect 3240 76780 3292 76832
rect 9772 76780 9824 76832
rect 2582 76678 2634 76730
rect 2646 76678 2698 76730
rect 2710 76678 2762 76730
rect 2774 76678 2826 76730
rect 2838 76678 2890 76730
rect 5846 76678 5898 76730
rect 5910 76678 5962 76730
rect 5974 76678 6026 76730
rect 6038 76678 6090 76730
rect 6102 76678 6154 76730
rect 9110 76678 9162 76730
rect 9174 76678 9226 76730
rect 9238 76678 9290 76730
rect 9302 76678 9354 76730
rect 9366 76678 9418 76730
rect 3056 76508 3108 76560
rect 1400 76372 1452 76424
rect 2780 76372 2832 76424
rect 3976 76415 4028 76424
rect 3976 76381 3985 76415
rect 3985 76381 4019 76415
rect 4019 76381 4028 76415
rect 3976 76372 4028 76381
rect 10140 76415 10192 76424
rect 10140 76381 10149 76415
rect 10149 76381 10183 76415
rect 10183 76381 10192 76415
rect 10140 76372 10192 76381
rect 1676 76236 1728 76288
rect 3240 76304 3292 76356
rect 2596 76236 2648 76288
rect 3792 76279 3844 76288
rect 3792 76245 3801 76279
rect 3801 76245 3835 76279
rect 3835 76245 3844 76279
rect 3792 76236 3844 76245
rect 4214 76134 4266 76186
rect 4278 76134 4330 76186
rect 4342 76134 4394 76186
rect 4406 76134 4458 76186
rect 4470 76134 4522 76186
rect 7478 76134 7530 76186
rect 7542 76134 7594 76186
rect 7606 76134 7658 76186
rect 7670 76134 7722 76186
rect 7734 76134 7786 76186
rect 1768 76032 1820 76084
rect 1584 75939 1636 75948
rect 1584 75905 1593 75939
rect 1593 75905 1627 75939
rect 1627 75905 1636 75939
rect 1584 75896 1636 75905
rect 5264 75964 5316 76016
rect 2596 75939 2648 75948
rect 2596 75905 2605 75939
rect 2605 75905 2639 75939
rect 2639 75905 2648 75939
rect 2596 75896 2648 75905
rect 2044 75828 2096 75880
rect 2780 75939 2832 75948
rect 2780 75905 2794 75939
rect 2794 75905 2828 75939
rect 2828 75905 2832 75939
rect 2780 75896 2832 75905
rect 3148 75896 3200 75948
rect 3700 75939 3752 75948
rect 3700 75905 3709 75939
rect 3709 75905 3743 75939
rect 3743 75905 3752 75939
rect 3700 75896 3752 75905
rect 10140 75939 10192 75948
rect 10140 75905 10149 75939
rect 10149 75905 10183 75939
rect 10183 75905 10192 75939
rect 10140 75896 10192 75905
rect 2320 75760 2372 75812
rect 2780 75760 2832 75812
rect 3516 75735 3568 75744
rect 3516 75701 3525 75735
rect 3525 75701 3559 75735
rect 3559 75701 3568 75735
rect 3516 75692 3568 75701
rect 2582 75590 2634 75642
rect 2646 75590 2698 75642
rect 2710 75590 2762 75642
rect 2774 75590 2826 75642
rect 2838 75590 2890 75642
rect 5846 75590 5898 75642
rect 5910 75590 5962 75642
rect 5974 75590 6026 75642
rect 6038 75590 6090 75642
rect 6102 75590 6154 75642
rect 9110 75590 9162 75642
rect 9174 75590 9226 75642
rect 9238 75590 9290 75642
rect 9302 75590 9354 75642
rect 9366 75590 9418 75642
rect 2504 75463 2556 75472
rect 2504 75429 2513 75463
rect 2513 75429 2547 75463
rect 2547 75429 2556 75463
rect 2504 75420 2556 75429
rect 2320 75327 2372 75336
rect 1860 75216 1912 75268
rect 2320 75293 2334 75327
rect 2334 75293 2368 75327
rect 2368 75293 2372 75327
rect 2320 75284 2372 75293
rect 10140 75327 10192 75336
rect 10140 75293 10149 75327
rect 10149 75293 10183 75327
rect 10183 75293 10192 75327
rect 10140 75284 10192 75293
rect 1492 75148 1544 75200
rect 2044 75148 2096 75200
rect 2964 75216 3016 75268
rect 4214 75046 4266 75098
rect 4278 75046 4330 75098
rect 4342 75046 4394 75098
rect 4406 75046 4458 75098
rect 4470 75046 4522 75098
rect 7478 75046 7530 75098
rect 7542 75046 7594 75098
rect 7606 75046 7658 75098
rect 7670 75046 7722 75098
rect 7734 75046 7786 75098
rect 3884 74876 3936 74928
rect 1492 74808 1544 74860
rect 1860 74851 1912 74860
rect 1860 74817 1863 74851
rect 1863 74817 1912 74851
rect 1860 74808 1912 74817
rect 2964 74808 3016 74860
rect 8300 74740 8352 74792
rect 2044 74672 2096 74724
rect 2320 74604 2372 74656
rect 2582 74502 2634 74554
rect 2646 74502 2698 74554
rect 2710 74502 2762 74554
rect 2774 74502 2826 74554
rect 2838 74502 2890 74554
rect 5846 74502 5898 74554
rect 5910 74502 5962 74554
rect 5974 74502 6026 74554
rect 6038 74502 6090 74554
rect 6102 74502 6154 74554
rect 9110 74502 9162 74554
rect 9174 74502 9226 74554
rect 9238 74502 9290 74554
rect 9302 74502 9354 74554
rect 9366 74502 9418 74554
rect 940 74332 992 74384
rect 1860 74128 1912 74180
rect 10140 74239 10192 74248
rect 10140 74205 10149 74239
rect 10149 74205 10183 74239
rect 10183 74205 10192 74239
rect 10140 74196 10192 74205
rect 1124 74060 1176 74112
rect 1492 74060 1544 74112
rect 3608 74128 3660 74180
rect 4214 73958 4266 74010
rect 4278 73958 4330 74010
rect 4342 73958 4394 74010
rect 4406 73958 4458 74010
rect 4470 73958 4522 74010
rect 7478 73958 7530 74010
rect 7542 73958 7594 74010
rect 7606 73958 7658 74010
rect 7670 73958 7722 74010
rect 7734 73958 7786 74010
rect 1400 73720 1452 73772
rect 2228 73763 2280 73772
rect 2228 73729 2237 73763
rect 2237 73729 2271 73763
rect 2271 73729 2280 73763
rect 2228 73720 2280 73729
rect 2872 73763 2924 73772
rect 2872 73729 2881 73763
rect 2881 73729 2915 73763
rect 2915 73729 2924 73763
rect 2872 73720 2924 73729
rect 10140 73763 10192 73772
rect 10140 73729 10149 73763
rect 10149 73729 10183 73763
rect 10183 73729 10192 73763
rect 10140 73720 10192 73729
rect 1308 73516 1360 73568
rect 1492 73516 1544 73568
rect 3148 73516 3200 73568
rect 8300 73516 8352 73568
rect 2582 73414 2634 73466
rect 2646 73414 2698 73466
rect 2710 73414 2762 73466
rect 2774 73414 2826 73466
rect 2838 73414 2890 73466
rect 5846 73414 5898 73466
rect 5910 73414 5962 73466
rect 5974 73414 6026 73466
rect 6038 73414 6090 73466
rect 6102 73414 6154 73466
rect 9110 73414 9162 73466
rect 9174 73414 9226 73466
rect 9238 73414 9290 73466
rect 9302 73414 9354 73466
rect 9366 73414 9418 73466
rect 2320 73176 2372 73228
rect 3332 73176 3384 73228
rect 1584 73151 1636 73160
rect 1584 73117 1593 73151
rect 1593 73117 1627 73151
rect 1627 73117 1636 73151
rect 1584 73108 1636 73117
rect 2780 73040 2832 73092
rect 3792 73040 3844 73092
rect 1216 72972 1268 73024
rect 4214 72870 4266 72922
rect 4278 72870 4330 72922
rect 4342 72870 4394 72922
rect 4406 72870 4458 72922
rect 4470 72870 4522 72922
rect 7478 72870 7530 72922
rect 7542 72870 7594 72922
rect 7606 72870 7658 72922
rect 7670 72870 7722 72922
rect 7734 72870 7786 72922
rect 1124 72700 1176 72752
rect 3516 72768 3568 72820
rect 1860 72675 1912 72684
rect 1860 72641 1863 72675
rect 1863 72641 1912 72675
rect 1860 72632 1912 72641
rect 8300 72700 8352 72752
rect 2688 72675 2740 72684
rect 2688 72641 2697 72675
rect 2697 72641 2731 72675
rect 2731 72641 2740 72675
rect 2688 72632 2740 72641
rect 2780 72675 2832 72684
rect 2780 72641 2789 72675
rect 2789 72641 2823 72675
rect 2823 72641 2832 72675
rect 2964 72675 3016 72684
rect 2780 72632 2832 72641
rect 2964 72641 2967 72675
rect 2967 72641 3016 72675
rect 2964 72632 3016 72641
rect 10140 72675 10192 72684
rect 10140 72641 10149 72675
rect 10149 72641 10183 72675
rect 10183 72641 10192 72675
rect 10140 72632 10192 72641
rect 9956 72564 10008 72616
rect 5540 72496 5592 72548
rect 1860 72428 1912 72480
rect 2964 72428 3016 72480
rect 3884 72428 3936 72480
rect 4620 72428 4672 72480
rect 2582 72326 2634 72378
rect 2646 72326 2698 72378
rect 2710 72326 2762 72378
rect 2774 72326 2826 72378
rect 2838 72326 2890 72378
rect 5846 72326 5898 72378
rect 5910 72326 5962 72378
rect 5974 72326 6026 72378
rect 6038 72326 6090 72378
rect 6102 72326 6154 72378
rect 9110 72326 9162 72378
rect 9174 72326 9226 72378
rect 9238 72326 9290 72378
rect 9302 72326 9354 72378
rect 9366 72326 9418 72378
rect 9956 72267 10008 72276
rect 9956 72233 9965 72267
rect 9965 72233 9999 72267
rect 9999 72233 10008 72267
rect 9956 72224 10008 72233
rect 1860 72156 1912 72208
rect 1584 72063 1636 72072
rect 1584 72029 1593 72063
rect 1593 72029 1627 72063
rect 1627 72029 1636 72063
rect 1584 72020 1636 72029
rect 2228 72063 2280 72072
rect 2228 72029 2237 72063
rect 2237 72029 2271 72063
rect 2271 72029 2280 72063
rect 2228 72020 2280 72029
rect 2872 72063 2924 72072
rect 2872 72029 2881 72063
rect 2881 72029 2915 72063
rect 2915 72029 2924 72063
rect 2872 72020 2924 72029
rect 10140 72063 10192 72072
rect 10140 72029 10149 72063
rect 10149 72029 10183 72063
rect 10183 72029 10192 72063
rect 10140 72020 10192 72029
rect 1032 71884 1084 71936
rect 2320 71884 2372 71936
rect 2596 71884 2648 71936
rect 4620 71884 4672 71936
rect 4214 71782 4266 71834
rect 4278 71782 4330 71834
rect 4342 71782 4394 71834
rect 4406 71782 4458 71834
rect 4470 71782 4522 71834
rect 7478 71782 7530 71834
rect 7542 71782 7594 71834
rect 7606 71782 7658 71834
rect 7670 71782 7722 71834
rect 7734 71782 7786 71834
rect 1124 71612 1176 71664
rect 1676 71655 1728 71664
rect 1676 71621 1685 71655
rect 1685 71621 1719 71655
rect 1719 71621 1728 71655
rect 1676 71612 1728 71621
rect 2412 71680 2464 71732
rect 2412 71544 2464 71596
rect 2596 71544 2648 71596
rect 2964 71587 3016 71596
rect 2964 71553 2967 71587
rect 2967 71553 3016 71587
rect 2964 71544 3016 71553
rect 3700 71544 3752 71596
rect 10140 71587 10192 71596
rect 10140 71553 10149 71587
rect 10149 71553 10183 71587
rect 10183 71553 10192 71587
rect 10140 71544 10192 71553
rect 1676 71408 1728 71460
rect 2044 71408 2096 71460
rect 5632 71408 5684 71460
rect 2582 71238 2634 71290
rect 2646 71238 2698 71290
rect 2710 71238 2762 71290
rect 2774 71238 2826 71290
rect 2838 71238 2890 71290
rect 5846 71238 5898 71290
rect 5910 71238 5962 71290
rect 5974 71238 6026 71290
rect 6038 71238 6090 71290
rect 6102 71238 6154 71290
rect 9110 71238 9162 71290
rect 9174 71238 9226 71290
rect 9238 71238 9290 71290
rect 9302 71238 9354 71290
rect 9366 71238 9418 71290
rect 1584 70975 1636 70984
rect 1584 70941 1593 70975
rect 1593 70941 1627 70975
rect 1627 70941 1636 70975
rect 1584 70932 1636 70941
rect 1492 70796 1544 70848
rect 4214 70694 4266 70746
rect 4278 70694 4330 70746
rect 4342 70694 4394 70746
rect 4406 70694 4458 70746
rect 4470 70694 4522 70746
rect 7478 70694 7530 70746
rect 7542 70694 7594 70746
rect 7606 70694 7658 70746
rect 7670 70694 7722 70746
rect 7734 70694 7786 70746
rect 1768 70592 1820 70644
rect 3516 70592 3568 70644
rect 1124 70524 1176 70576
rect 2412 70524 2464 70576
rect 2964 70524 3016 70576
rect 2044 70456 2096 70508
rect 10140 70499 10192 70508
rect 10140 70465 10149 70499
rect 10149 70465 10183 70499
rect 10183 70465 10192 70499
rect 10140 70456 10192 70465
rect 1492 70252 1544 70304
rect 1860 70252 1912 70304
rect 2412 70252 2464 70304
rect 2582 70150 2634 70202
rect 2646 70150 2698 70202
rect 2710 70150 2762 70202
rect 2774 70150 2826 70202
rect 2838 70150 2890 70202
rect 5846 70150 5898 70202
rect 5910 70150 5962 70202
rect 5974 70150 6026 70202
rect 6038 70150 6090 70202
rect 6102 70150 6154 70202
rect 9110 70150 9162 70202
rect 9174 70150 9226 70202
rect 9238 70150 9290 70202
rect 9302 70150 9354 70202
rect 9366 70150 9418 70202
rect 1584 69887 1636 69896
rect 1584 69853 1593 69887
rect 1593 69853 1627 69887
rect 1627 69853 1636 69887
rect 1584 69844 1636 69853
rect 2228 69887 2280 69896
rect 2228 69853 2237 69887
rect 2237 69853 2271 69887
rect 2271 69853 2280 69887
rect 2228 69844 2280 69853
rect 2872 69887 2924 69896
rect 2872 69853 2881 69887
rect 2881 69853 2915 69887
rect 2915 69853 2924 69887
rect 2872 69844 2924 69853
rect 10140 69887 10192 69896
rect 10140 69853 10149 69887
rect 10149 69853 10183 69887
rect 10183 69853 10192 69887
rect 10140 69844 10192 69853
rect 1308 69776 1360 69828
rect 756 69708 808 69760
rect 1584 69708 1636 69760
rect 2044 69751 2096 69760
rect 2044 69717 2053 69751
rect 2053 69717 2087 69751
rect 2087 69717 2096 69751
rect 2044 69708 2096 69717
rect 2688 69751 2740 69760
rect 2688 69717 2697 69751
rect 2697 69717 2731 69751
rect 2731 69717 2740 69751
rect 2688 69708 2740 69717
rect 3056 69708 3108 69760
rect 3792 69708 3844 69760
rect 9956 69751 10008 69760
rect 9956 69717 9965 69751
rect 9965 69717 9999 69751
rect 9999 69717 10008 69751
rect 9956 69708 10008 69717
rect 4214 69606 4266 69658
rect 4278 69606 4330 69658
rect 4342 69606 4394 69658
rect 4406 69606 4458 69658
rect 4470 69606 4522 69658
rect 7478 69606 7530 69658
rect 7542 69606 7594 69658
rect 7606 69606 7658 69658
rect 7670 69606 7722 69658
rect 7734 69606 7786 69658
rect 1124 69436 1176 69488
rect 1676 69479 1728 69488
rect 1676 69445 1685 69479
rect 1685 69445 1719 69479
rect 1719 69445 1728 69479
rect 1676 69436 1728 69445
rect 1492 69368 1544 69420
rect 3056 69436 3108 69488
rect 2964 69368 3016 69420
rect 9956 69300 10008 69352
rect 5724 69232 5776 69284
rect 1124 69164 1176 69216
rect 2582 69062 2634 69114
rect 2646 69062 2698 69114
rect 2710 69062 2762 69114
rect 2774 69062 2826 69114
rect 2838 69062 2890 69114
rect 5846 69062 5898 69114
rect 5910 69062 5962 69114
rect 5974 69062 6026 69114
rect 6038 69062 6090 69114
rect 6102 69062 6154 69114
rect 9110 69062 9162 69114
rect 9174 69062 9226 69114
rect 9238 69062 9290 69114
rect 9302 69062 9354 69114
rect 9366 69062 9418 69114
rect 1584 68799 1636 68808
rect 1584 68765 1593 68799
rect 1593 68765 1627 68799
rect 1627 68765 1636 68799
rect 1584 68756 1636 68765
rect 4068 68892 4120 68944
rect 2872 68756 2924 68808
rect 3056 68756 3108 68808
rect 10140 68799 10192 68808
rect 10140 68765 10149 68799
rect 10149 68765 10183 68799
rect 10183 68765 10192 68799
rect 10140 68756 10192 68765
rect 1492 68688 1544 68740
rect 2504 68731 2556 68740
rect 2504 68697 2513 68731
rect 2513 68697 2547 68731
rect 2547 68697 2556 68731
rect 2504 68688 2556 68697
rect 3148 68688 3200 68740
rect 2228 68620 2280 68672
rect 4214 68518 4266 68570
rect 4278 68518 4330 68570
rect 4342 68518 4394 68570
rect 4406 68518 4458 68570
rect 4470 68518 4522 68570
rect 7478 68518 7530 68570
rect 7542 68518 7594 68570
rect 7606 68518 7658 68570
rect 7670 68518 7722 68570
rect 7734 68518 7786 68570
rect 664 68280 716 68332
rect 10140 68323 10192 68332
rect 10140 68289 10149 68323
rect 10149 68289 10183 68323
rect 10183 68289 10192 68323
rect 10140 68280 10192 68289
rect 1308 68212 1360 68264
rect 8300 68076 8352 68128
rect 2582 67974 2634 68026
rect 2646 67974 2698 68026
rect 2710 67974 2762 68026
rect 2774 67974 2826 68026
rect 2838 67974 2890 68026
rect 5846 67974 5898 68026
rect 5910 67974 5962 68026
rect 5974 67974 6026 68026
rect 6038 67974 6090 68026
rect 6102 67974 6154 68026
rect 9110 67974 9162 68026
rect 9174 67974 9226 68026
rect 9238 67974 9290 68026
rect 9302 67974 9354 68026
rect 9366 67974 9418 68026
rect 1400 67711 1452 67720
rect 1400 67677 1409 67711
rect 1409 67677 1443 67711
rect 1443 67677 1452 67711
rect 1400 67668 1452 67677
rect 1676 67711 1728 67720
rect 1676 67677 1685 67711
rect 1685 67677 1719 67711
rect 1719 67677 1728 67711
rect 1676 67668 1728 67677
rect 3516 67600 3568 67652
rect 4804 67600 4856 67652
rect 4214 67430 4266 67482
rect 4278 67430 4330 67482
rect 4342 67430 4394 67482
rect 4406 67430 4458 67482
rect 4470 67430 4522 67482
rect 7478 67430 7530 67482
rect 7542 67430 7594 67482
rect 7606 67430 7658 67482
rect 7670 67430 7722 67482
rect 7734 67430 7786 67482
rect 2228 67260 2280 67312
rect 2412 67260 2464 67312
rect 3056 67192 3108 67244
rect 10140 67235 10192 67244
rect 10140 67201 10149 67235
rect 10149 67201 10183 67235
rect 10183 67201 10192 67235
rect 10140 67192 10192 67201
rect 1400 67167 1452 67176
rect 1400 67133 1409 67167
rect 1409 67133 1443 67167
rect 1443 67133 1452 67167
rect 1400 67124 1452 67133
rect 2412 67124 2464 67176
rect 848 67056 900 67108
rect 1676 66988 1728 67040
rect 1860 66988 1912 67040
rect 5448 66988 5500 67040
rect 2582 66886 2634 66938
rect 2646 66886 2698 66938
rect 2710 66886 2762 66938
rect 2774 66886 2826 66938
rect 2838 66886 2890 66938
rect 5846 66886 5898 66938
rect 5910 66886 5962 66938
rect 5974 66886 6026 66938
rect 6038 66886 6090 66938
rect 6102 66886 6154 66938
rect 9110 66886 9162 66938
rect 9174 66886 9226 66938
rect 9238 66886 9290 66938
rect 9302 66886 9354 66938
rect 9366 66886 9418 66938
rect 8300 66784 8352 66836
rect 5172 66716 5224 66768
rect 1492 66648 1544 66700
rect 2964 66648 3016 66700
rect 3148 66648 3200 66700
rect 1308 66512 1360 66564
rect 2504 66623 2556 66632
rect 2504 66589 2513 66623
rect 2513 66589 2547 66623
rect 2547 66589 2556 66623
rect 2504 66580 2556 66589
rect 10140 66623 10192 66632
rect 10140 66589 10149 66623
rect 10149 66589 10183 66623
rect 10183 66589 10192 66623
rect 10140 66580 10192 66589
rect 2596 66444 2648 66496
rect 2964 66444 3016 66496
rect 8300 66444 8352 66496
rect 4214 66342 4266 66394
rect 4278 66342 4330 66394
rect 4342 66342 4394 66394
rect 4406 66342 4458 66394
rect 4470 66342 4522 66394
rect 7478 66342 7530 66394
rect 7542 66342 7594 66394
rect 7606 66342 7658 66394
rect 7670 66342 7722 66394
rect 7734 66342 7786 66394
rect 1124 66240 1176 66292
rect 1492 66240 1544 66292
rect 1584 66240 1636 66292
rect 1584 66104 1636 66156
rect 3148 66172 3200 66224
rect 10140 66147 10192 66156
rect 1308 65968 1360 66020
rect 10140 66113 10149 66147
rect 10149 66113 10183 66147
rect 10183 66113 10192 66147
rect 10140 66104 10192 66113
rect 1032 65900 1084 65952
rect 4988 65968 5040 66020
rect 3056 65900 3108 65952
rect 9956 65943 10008 65952
rect 9956 65909 9965 65943
rect 9965 65909 9999 65943
rect 9999 65909 10008 65943
rect 9956 65900 10008 65909
rect 2582 65798 2634 65850
rect 2646 65798 2698 65850
rect 2710 65798 2762 65850
rect 2774 65798 2826 65850
rect 2838 65798 2890 65850
rect 5846 65798 5898 65850
rect 5910 65798 5962 65850
rect 5974 65798 6026 65850
rect 6038 65798 6090 65850
rect 6102 65798 6154 65850
rect 9110 65798 9162 65850
rect 9174 65798 9226 65850
rect 9238 65798 9290 65850
rect 9302 65798 9354 65850
rect 9366 65798 9418 65850
rect 1768 65560 1820 65612
rect 1584 65535 1636 65544
rect 1584 65501 1593 65535
rect 1593 65501 1627 65535
rect 1627 65501 1636 65535
rect 1584 65492 1636 65501
rect 9956 65560 10008 65612
rect 2964 65492 3016 65544
rect 3608 65492 3660 65544
rect 388 65356 440 65408
rect 1860 65356 1912 65408
rect 2780 65424 2832 65476
rect 7840 65424 7892 65476
rect 3700 65356 3752 65408
rect 3976 65399 4028 65408
rect 3976 65365 3985 65399
rect 3985 65365 4019 65399
rect 4019 65365 4028 65399
rect 3976 65356 4028 65365
rect 4214 65254 4266 65306
rect 4278 65254 4330 65306
rect 4342 65254 4394 65306
rect 4406 65254 4458 65306
rect 4470 65254 4522 65306
rect 7478 65254 7530 65306
rect 7542 65254 7594 65306
rect 7606 65254 7658 65306
rect 7670 65254 7722 65306
rect 7734 65254 7786 65306
rect 8300 65152 8352 65204
rect 1492 65084 1544 65136
rect 3240 65084 3292 65136
rect 3700 65084 3752 65136
rect 4896 65084 4948 65136
rect 1308 64948 1360 65000
rect 1400 64880 1452 64932
rect 1860 64948 1912 65000
rect 2964 65016 3016 65068
rect 3148 65016 3200 65068
rect 3516 65059 3568 65068
rect 2780 64948 2832 65000
rect 3516 65025 3525 65059
rect 3525 65025 3559 65059
rect 3559 65025 3568 65059
rect 3516 65016 3568 65025
rect 10140 65059 10192 65068
rect 10140 65025 10149 65059
rect 10149 65025 10183 65059
rect 10183 65025 10192 65059
rect 10140 65016 10192 65025
rect 3148 64880 3200 64932
rect 8300 64880 8352 64932
rect 3240 64812 3292 64864
rect 3516 64812 3568 64864
rect 2582 64710 2634 64762
rect 2646 64710 2698 64762
rect 2710 64710 2762 64762
rect 2774 64710 2826 64762
rect 2838 64710 2890 64762
rect 5846 64710 5898 64762
rect 5910 64710 5962 64762
rect 5974 64710 6026 64762
rect 6038 64710 6090 64762
rect 6102 64710 6154 64762
rect 9110 64710 9162 64762
rect 9174 64710 9226 64762
rect 9238 64710 9290 64762
rect 9302 64710 9354 64762
rect 9366 64710 9418 64762
rect 1768 64540 1820 64592
rect 2228 64540 2280 64592
rect 3516 64540 3568 64592
rect 8300 64472 8352 64524
rect 2228 64447 2280 64456
rect 2228 64413 2237 64447
rect 2237 64413 2271 64447
rect 2271 64413 2280 64447
rect 2228 64404 2280 64413
rect 2964 64404 3016 64456
rect 4068 64404 4120 64456
rect 10140 64447 10192 64456
rect 10140 64413 10149 64447
rect 10149 64413 10183 64447
rect 10183 64413 10192 64447
rect 10140 64404 10192 64413
rect 1860 64336 1912 64388
rect 3056 64268 3108 64320
rect 8300 64268 8352 64320
rect 4214 64166 4266 64218
rect 4278 64166 4330 64218
rect 4342 64166 4394 64218
rect 4406 64166 4458 64218
rect 4470 64166 4522 64218
rect 7478 64166 7530 64218
rect 7542 64166 7594 64218
rect 7606 64166 7658 64218
rect 7670 64166 7722 64218
rect 7734 64166 7786 64218
rect 1308 63996 1360 64048
rect 296 63928 348 63980
rect 3240 63928 3292 63980
rect 3700 63928 3752 63980
rect 2964 63860 3016 63912
rect 1584 63767 1636 63776
rect 1584 63733 1593 63767
rect 1593 63733 1627 63767
rect 1627 63733 1636 63767
rect 1584 63724 1636 63733
rect 2582 63622 2634 63674
rect 2646 63622 2698 63674
rect 2710 63622 2762 63674
rect 2774 63622 2826 63674
rect 2838 63622 2890 63674
rect 5846 63622 5898 63674
rect 5910 63622 5962 63674
rect 5974 63622 6026 63674
rect 6038 63622 6090 63674
rect 6102 63622 6154 63674
rect 9110 63622 9162 63674
rect 9174 63622 9226 63674
rect 9238 63622 9290 63674
rect 9302 63622 9354 63674
rect 9366 63622 9418 63674
rect 1676 63452 1728 63504
rect 3056 63495 3108 63504
rect 3056 63461 3065 63495
rect 3065 63461 3099 63495
rect 3099 63461 3108 63495
rect 3056 63452 3108 63461
rect 1676 63316 1728 63368
rect 2872 63359 2924 63368
rect 2872 63325 2881 63359
rect 2881 63325 2915 63359
rect 2915 63325 2924 63359
rect 2872 63316 2924 63325
rect 10140 63359 10192 63368
rect 10140 63325 10149 63359
rect 10149 63325 10183 63359
rect 10183 63325 10192 63359
rect 10140 63316 10192 63325
rect 3240 63248 3292 63300
rect 1400 63180 1452 63232
rect 8484 63180 8536 63232
rect 572 63112 624 63164
rect 940 63112 992 63164
rect 4214 63078 4266 63130
rect 4278 63078 4330 63130
rect 4342 63078 4394 63130
rect 4406 63078 4458 63130
rect 4470 63078 4522 63130
rect 7478 63078 7530 63130
rect 7542 63078 7594 63130
rect 7606 63078 7658 63130
rect 7670 63078 7722 63130
rect 7734 63078 7786 63130
rect 1032 62840 1084 62892
rect 3056 62840 3108 62892
rect 10140 62883 10192 62892
rect 10140 62849 10149 62883
rect 10149 62849 10183 62883
rect 10183 62849 10192 62883
rect 10140 62840 10192 62849
rect 1584 62679 1636 62688
rect 1584 62645 1593 62679
rect 1593 62645 1627 62679
rect 1627 62645 1636 62679
rect 1584 62636 1636 62645
rect 2320 62679 2372 62688
rect 2320 62645 2329 62679
rect 2329 62645 2363 62679
rect 2363 62645 2372 62679
rect 2320 62636 2372 62645
rect 6184 62636 6236 62688
rect 2582 62534 2634 62586
rect 2646 62534 2698 62586
rect 2710 62534 2762 62586
rect 2774 62534 2826 62586
rect 2838 62534 2890 62586
rect 5846 62534 5898 62586
rect 5910 62534 5962 62586
rect 5974 62534 6026 62586
rect 6038 62534 6090 62586
rect 6102 62534 6154 62586
rect 9110 62534 9162 62586
rect 9174 62534 9226 62586
rect 9238 62534 9290 62586
rect 9302 62534 9354 62586
rect 9366 62534 9418 62586
rect 5356 62364 5408 62416
rect 8300 62296 8352 62348
rect 1124 62160 1176 62212
rect 2412 62271 2464 62280
rect 2412 62237 2415 62271
rect 2415 62237 2464 62271
rect 2412 62228 2464 62237
rect 2964 62228 3016 62280
rect 10140 62271 10192 62280
rect 10140 62237 10149 62271
rect 10149 62237 10183 62271
rect 10183 62237 10192 62271
rect 10140 62228 10192 62237
rect 1860 62092 1912 62144
rect 2596 62160 2648 62212
rect 2964 62092 3016 62144
rect 3516 62092 3568 62144
rect 8300 62092 8352 62144
rect 4214 61990 4266 62042
rect 4278 61990 4330 62042
rect 4342 61990 4394 62042
rect 4406 61990 4458 62042
rect 4470 61990 4522 62042
rect 7478 61990 7530 62042
rect 7542 61990 7594 62042
rect 7606 61990 7658 62042
rect 7670 61990 7722 62042
rect 7734 61990 7786 62042
rect 9956 61820 10008 61872
rect 1492 61752 1544 61804
rect 1768 61795 1820 61804
rect 1768 61761 1782 61795
rect 1782 61761 1816 61795
rect 1816 61761 1820 61795
rect 1768 61752 1820 61761
rect 2412 61752 2464 61804
rect 2688 61752 2740 61804
rect 3516 61795 3568 61804
rect 3516 61761 3525 61795
rect 3525 61761 3559 61795
rect 3559 61761 3568 61795
rect 3516 61752 3568 61761
rect 2228 61684 2280 61736
rect 2596 61616 2648 61668
rect 3700 61659 3752 61668
rect 3700 61625 3709 61659
rect 3709 61625 3743 61659
rect 3743 61625 3752 61659
rect 3700 61616 3752 61625
rect 1860 61548 1912 61600
rect 2136 61548 2188 61600
rect 2412 61548 2464 61600
rect 2582 61446 2634 61498
rect 2646 61446 2698 61498
rect 2710 61446 2762 61498
rect 2774 61446 2826 61498
rect 2838 61446 2890 61498
rect 5846 61446 5898 61498
rect 5910 61446 5962 61498
rect 5974 61446 6026 61498
rect 6038 61446 6090 61498
rect 6102 61446 6154 61498
rect 9110 61446 9162 61498
rect 9174 61446 9226 61498
rect 9238 61446 9290 61498
rect 9302 61446 9354 61498
rect 9366 61446 9418 61498
rect 9956 61387 10008 61396
rect 9956 61353 9965 61387
rect 9965 61353 9999 61387
rect 9999 61353 10008 61387
rect 9956 61344 10008 61353
rect 2228 61276 2280 61328
rect 8300 61208 8352 61260
rect 1768 61183 1820 61192
rect 1768 61149 1782 61183
rect 1782 61149 1816 61183
rect 1816 61149 1820 61183
rect 1768 61140 1820 61149
rect 10140 61183 10192 61192
rect 1124 61072 1176 61124
rect 1492 61072 1544 61124
rect 1676 61115 1728 61124
rect 1676 61081 1685 61115
rect 1685 61081 1719 61115
rect 1719 61081 1728 61115
rect 1676 61072 1728 61081
rect 20 61004 72 61056
rect 10140 61149 10149 61183
rect 10149 61149 10183 61183
rect 10183 61149 10192 61183
rect 10140 61140 10192 61149
rect 2780 61004 2832 61056
rect 4214 60902 4266 60954
rect 4278 60902 4330 60954
rect 4342 60902 4394 60954
rect 4406 60902 4458 60954
rect 4470 60902 4522 60954
rect 7478 60902 7530 60954
rect 7542 60902 7594 60954
rect 7606 60902 7658 60954
rect 7670 60902 7722 60954
rect 7734 60902 7786 60954
rect 848 60800 900 60852
rect 1216 60800 1268 60852
rect 1676 60800 1728 60852
rect 1952 60800 2004 60852
rect 2688 60800 2740 60852
rect 1492 60732 1544 60784
rect 1768 60664 1820 60716
rect 3240 60664 3292 60716
rect 3424 60664 3476 60716
rect 10140 60707 10192 60716
rect 10140 60673 10149 60707
rect 10149 60673 10183 60707
rect 10183 60673 10192 60707
rect 10140 60664 10192 60673
rect 3976 60596 4028 60648
rect 1216 60460 1268 60512
rect 2964 60528 3016 60580
rect 1584 60503 1636 60512
rect 1584 60469 1593 60503
rect 1593 60469 1627 60503
rect 1627 60469 1636 60503
rect 1584 60460 1636 60469
rect 2320 60503 2372 60512
rect 2320 60469 2329 60503
rect 2329 60469 2363 60503
rect 2363 60469 2372 60503
rect 2320 60460 2372 60469
rect 9956 60503 10008 60512
rect 9956 60469 9965 60503
rect 9965 60469 9999 60503
rect 9999 60469 10008 60503
rect 9956 60460 10008 60469
rect 2582 60358 2634 60410
rect 2646 60358 2698 60410
rect 2710 60358 2762 60410
rect 2774 60358 2826 60410
rect 2838 60358 2890 60410
rect 5846 60358 5898 60410
rect 5910 60358 5962 60410
rect 5974 60358 6026 60410
rect 6038 60358 6090 60410
rect 6102 60358 6154 60410
rect 9110 60358 9162 60410
rect 9174 60358 9226 60410
rect 9238 60358 9290 60410
rect 9302 60358 9354 60410
rect 9366 60358 9418 60410
rect 112 60256 164 60308
rect 1768 60256 1820 60308
rect 572 60188 624 60240
rect 1308 60188 1360 60240
rect 2228 60188 2280 60240
rect 2688 60188 2740 60240
rect 756 60120 808 60172
rect 2596 60120 2648 60172
rect 480 60052 532 60104
rect 1768 59984 1820 60036
rect 2504 59984 2556 60036
rect 2044 59916 2096 59968
rect 2780 59916 2832 59968
rect 4214 59814 4266 59866
rect 4278 59814 4330 59866
rect 4342 59814 4394 59866
rect 4406 59814 4458 59866
rect 4470 59814 4522 59866
rect 7478 59814 7530 59866
rect 7542 59814 7594 59866
rect 7606 59814 7658 59866
rect 7670 59814 7722 59866
rect 7734 59814 7786 59866
rect 1124 59712 1176 59764
rect 2044 59712 2096 59764
rect 2596 59712 2648 59764
rect 1124 59576 1176 59628
rect 2136 59619 2188 59628
rect 2136 59585 2145 59619
rect 2145 59585 2179 59619
rect 2179 59585 2188 59619
rect 2136 59576 2188 59585
rect 756 59372 808 59424
rect 2596 59619 2648 59628
rect 2596 59585 2599 59619
rect 2599 59585 2648 59619
rect 2596 59576 2648 59585
rect 10140 59619 10192 59628
rect 10140 59585 10149 59619
rect 10149 59585 10183 59619
rect 10183 59585 10192 59619
rect 10140 59576 10192 59585
rect 2688 59508 2740 59560
rect 5080 59508 5132 59560
rect 9956 59508 10008 59560
rect 2320 59440 2372 59492
rect 2412 59440 2464 59492
rect 2136 59372 2188 59424
rect 2228 59372 2280 59424
rect 3240 59372 3292 59424
rect 3700 59372 3752 59424
rect 3976 59372 4028 59424
rect 4620 59372 4672 59424
rect 8300 59372 8352 59424
rect 2582 59270 2634 59322
rect 2646 59270 2698 59322
rect 2710 59270 2762 59322
rect 2774 59270 2826 59322
rect 2838 59270 2890 59322
rect 5846 59270 5898 59322
rect 5910 59270 5962 59322
rect 5974 59270 6026 59322
rect 6038 59270 6090 59322
rect 6102 59270 6154 59322
rect 9110 59270 9162 59322
rect 9174 59270 9226 59322
rect 9238 59270 9290 59322
rect 9302 59270 9354 59322
rect 9366 59270 9418 59322
rect 1952 59168 2004 59220
rect 2044 59168 2096 59220
rect 2320 59168 2372 59220
rect 572 59100 624 59152
rect 1584 59007 1636 59016
rect 1584 58973 1593 59007
rect 1593 58973 1627 59007
rect 1627 58973 1636 59007
rect 1584 58964 1636 58973
rect 8484 59032 8536 59084
rect 1400 58896 1452 58948
rect 2596 58896 2648 58948
rect 388 58828 440 58880
rect 2044 58828 2096 58880
rect 2136 58828 2188 58880
rect 4712 58964 4764 59016
rect 10140 59007 10192 59016
rect 10140 58973 10149 59007
rect 10149 58973 10183 59007
rect 10183 58973 10192 59007
rect 10140 58964 10192 58973
rect 3976 58871 4028 58880
rect 3976 58837 3985 58871
rect 3985 58837 4019 58871
rect 4019 58837 4028 58871
rect 3976 58828 4028 58837
rect 9956 58871 10008 58880
rect 9956 58837 9965 58871
rect 9965 58837 9999 58871
rect 9999 58837 10008 58871
rect 9956 58828 10008 58837
rect 4214 58726 4266 58778
rect 4278 58726 4330 58778
rect 4342 58726 4394 58778
rect 4406 58726 4458 58778
rect 4470 58726 4522 58778
rect 7478 58726 7530 58778
rect 7542 58726 7594 58778
rect 7606 58726 7658 58778
rect 7670 58726 7722 58778
rect 7734 58726 7786 58778
rect 1584 58624 1636 58676
rect 756 58556 808 58608
rect 2228 58556 2280 58608
rect 2320 58556 2372 58608
rect 2596 58556 2648 58608
rect 3516 58556 3568 58608
rect 3976 58556 4028 58608
rect 204 58488 256 58540
rect 1952 58488 2004 58540
rect 2688 58531 2740 58540
rect 2688 58497 2697 58531
rect 2697 58497 2731 58531
rect 2731 58497 2740 58531
rect 2688 58488 2740 58497
rect 3700 58488 3752 58540
rect 5080 58488 5132 58540
rect 4160 58420 4212 58472
rect 9496 58420 9548 58472
rect 3516 58395 3568 58404
rect 3516 58361 3525 58395
rect 3525 58361 3559 58395
rect 3559 58361 3568 58395
rect 3516 58352 3568 58361
rect 1400 58284 1452 58336
rect 2582 58182 2634 58234
rect 2646 58182 2698 58234
rect 2710 58182 2762 58234
rect 2774 58182 2826 58234
rect 2838 58182 2890 58234
rect 5846 58182 5898 58234
rect 5910 58182 5962 58234
rect 5974 58182 6026 58234
rect 6038 58182 6090 58234
rect 6102 58182 6154 58234
rect 9110 58182 9162 58234
rect 9174 58182 9226 58234
rect 9238 58182 9290 58234
rect 9302 58182 9354 58234
rect 9366 58182 9418 58234
rect 3516 58080 3568 58132
rect 4160 58080 4212 58132
rect 2780 58012 2832 58064
rect 3240 58012 3292 58064
rect 756 57876 808 57928
rect 388 57808 440 57860
rect 1584 57783 1636 57792
rect 1584 57749 1593 57783
rect 1593 57749 1627 57783
rect 1627 57749 1636 57783
rect 1584 57740 1636 57749
rect 2596 57740 2648 57792
rect 4214 57638 4266 57690
rect 4278 57638 4330 57690
rect 4342 57638 4394 57690
rect 4406 57638 4458 57690
rect 4470 57638 4522 57690
rect 7478 57638 7530 57690
rect 7542 57638 7594 57690
rect 7606 57638 7658 57690
rect 7670 57638 7722 57690
rect 7734 57638 7786 57690
rect 1768 57536 1820 57588
rect 1768 57400 1820 57452
rect 2136 57400 2188 57452
rect 6552 57400 6604 57452
rect 2320 57332 2372 57384
rect 3056 57332 3108 57384
rect 3240 57332 3292 57384
rect 9496 57332 9548 57384
rect 9956 57264 10008 57316
rect 2136 57196 2188 57248
rect 2582 57094 2634 57146
rect 2646 57094 2698 57146
rect 2710 57094 2762 57146
rect 2774 57094 2826 57146
rect 2838 57094 2890 57146
rect 5846 57094 5898 57146
rect 5910 57094 5962 57146
rect 5974 57094 6026 57146
rect 6038 57094 6090 57146
rect 6102 57094 6154 57146
rect 9110 57094 9162 57146
rect 9174 57094 9226 57146
rect 9238 57094 9290 57146
rect 9302 57094 9354 57146
rect 9366 57094 9418 57146
rect 848 56992 900 57044
rect 1952 56967 2004 56976
rect 1952 56933 1961 56967
rect 1961 56933 1995 56967
rect 1995 56933 2004 56967
rect 1952 56924 2004 56933
rect 8300 56856 8352 56908
rect 8484 56856 8536 56908
rect 1676 56831 1728 56840
rect 1676 56797 1685 56831
rect 1685 56797 1719 56831
rect 1719 56797 1728 56831
rect 1676 56788 1728 56797
rect 1768 56831 1820 56840
rect 1768 56797 1782 56831
rect 1782 56797 1816 56831
rect 1816 56797 1820 56831
rect 1768 56788 1820 56797
rect 2320 56788 2372 56840
rect 3056 56788 3108 56840
rect 9312 56831 9364 56840
rect 9312 56797 9321 56831
rect 9321 56797 9355 56831
rect 9355 56797 9364 56831
rect 9312 56788 9364 56797
rect 1584 56763 1636 56772
rect 1584 56729 1593 56763
rect 1593 56729 1627 56763
rect 1627 56729 1636 56763
rect 1584 56720 1636 56729
rect 2412 56720 2464 56772
rect 4214 56550 4266 56602
rect 4278 56550 4330 56602
rect 4342 56550 4394 56602
rect 4406 56550 4458 56602
rect 4470 56550 4522 56602
rect 7478 56550 7530 56602
rect 7542 56550 7594 56602
rect 7606 56550 7658 56602
rect 7670 56550 7722 56602
rect 7734 56550 7786 56602
rect 1676 56448 1728 56500
rect 3608 56491 3660 56500
rect 3608 56457 3617 56491
rect 3617 56457 3651 56491
rect 3651 56457 3660 56491
rect 3608 56448 3660 56457
rect 1768 56380 1820 56432
rect 1492 56312 1544 56364
rect 1676 56312 1728 56364
rect 1216 56244 1268 56296
rect 3608 56312 3660 56364
rect 10140 56355 10192 56364
rect 10140 56321 10149 56355
rect 10149 56321 10183 56355
rect 10183 56321 10192 56355
rect 10140 56312 10192 56321
rect 6368 56244 6420 56296
rect 2688 56176 2740 56228
rect 2320 56151 2372 56160
rect 2320 56117 2329 56151
rect 2329 56117 2363 56151
rect 2363 56117 2372 56151
rect 2320 56108 2372 56117
rect 4988 56108 5040 56160
rect 5448 56108 5500 56160
rect 6184 56108 6236 56160
rect 2582 56006 2634 56058
rect 2646 56006 2698 56058
rect 2710 56006 2762 56058
rect 2774 56006 2826 56058
rect 2838 56006 2890 56058
rect 5846 56006 5898 56058
rect 5910 56006 5962 56058
rect 5974 56006 6026 56058
rect 6038 56006 6090 56058
rect 6102 56006 6154 56058
rect 9110 56006 9162 56058
rect 9174 56006 9226 56058
rect 9238 56006 9290 56058
rect 9302 56006 9354 56058
rect 9366 56006 9418 56058
rect 4988 55836 5040 55888
rect 5356 55836 5408 55888
rect 848 55700 900 55752
rect 2872 55743 2924 55752
rect 2872 55709 2881 55743
rect 2881 55709 2915 55743
rect 2915 55709 2924 55743
rect 3240 55768 3292 55820
rect 2872 55700 2924 55709
rect 3516 55700 3568 55752
rect 4160 55700 4212 55752
rect 9588 55700 9640 55752
rect 6460 55632 6512 55684
rect 1584 55607 1636 55616
rect 1584 55573 1593 55607
rect 1593 55573 1627 55607
rect 1627 55573 1636 55607
rect 1584 55564 1636 55573
rect 2320 55607 2372 55616
rect 2320 55573 2329 55607
rect 2329 55573 2363 55607
rect 2363 55573 2372 55607
rect 2320 55564 2372 55573
rect 3240 55607 3292 55616
rect 3240 55573 3249 55607
rect 3249 55573 3283 55607
rect 3283 55573 3292 55607
rect 3240 55564 3292 55573
rect 6828 55564 6880 55616
rect 8300 55564 8352 55616
rect 572 55496 624 55548
rect 4214 55462 4266 55514
rect 4278 55462 4330 55514
rect 4342 55462 4394 55514
rect 4406 55462 4458 55514
rect 4470 55462 4522 55514
rect 7478 55462 7530 55514
rect 7542 55462 7594 55514
rect 7606 55462 7658 55514
rect 7670 55462 7722 55514
rect 7734 55462 7786 55514
rect 3056 55360 3108 55412
rect 3240 55360 3292 55412
rect 3608 55403 3660 55412
rect 3608 55369 3617 55403
rect 3617 55369 3651 55403
rect 3651 55369 3660 55403
rect 3608 55360 3660 55369
rect 10140 55360 10192 55412
rect 1308 55292 1360 55344
rect 1768 55224 1820 55276
rect 3608 55224 3660 55276
rect 1308 55088 1360 55140
rect 664 55020 716 55072
rect 1124 55020 1176 55072
rect 1492 55020 1544 55072
rect 3516 55156 3568 55208
rect 3148 55088 3200 55140
rect 4344 55156 4396 55208
rect 9864 55020 9916 55072
rect 2582 54918 2634 54970
rect 2646 54918 2698 54970
rect 2710 54918 2762 54970
rect 2774 54918 2826 54970
rect 2838 54918 2890 54970
rect 5846 54918 5898 54970
rect 5910 54918 5962 54970
rect 5974 54918 6026 54970
rect 6038 54918 6090 54970
rect 6102 54918 6154 54970
rect 9110 54918 9162 54970
rect 9174 54918 9226 54970
rect 9238 54918 9290 54970
rect 9302 54918 9354 54970
rect 9366 54918 9418 54970
rect 3516 54816 3568 54868
rect 4068 54816 4120 54868
rect 1676 54748 1728 54800
rect 2412 54748 2464 54800
rect 2320 54612 2372 54664
rect 6276 54612 6328 54664
rect 6828 54612 6880 54664
rect 10140 54655 10192 54664
rect 10140 54621 10149 54655
rect 10149 54621 10183 54655
rect 10183 54621 10192 54655
rect 10140 54612 10192 54621
rect 1584 54587 1636 54596
rect 1584 54553 1593 54587
rect 1593 54553 1627 54587
rect 1627 54553 1636 54587
rect 1584 54544 1636 54553
rect 6184 54544 6236 54596
rect 2780 54476 2832 54528
rect 9680 54476 9732 54528
rect 9956 54519 10008 54528
rect 9956 54485 9965 54519
rect 9965 54485 9999 54519
rect 9999 54485 10008 54519
rect 9956 54476 10008 54485
rect 4214 54374 4266 54426
rect 4278 54374 4330 54426
rect 4342 54374 4394 54426
rect 4406 54374 4458 54426
rect 4470 54374 4522 54426
rect 7478 54374 7530 54426
rect 7542 54374 7594 54426
rect 7606 54374 7658 54426
rect 7670 54374 7722 54426
rect 7734 54374 7786 54426
rect 1400 54272 1452 54324
rect 1676 54272 1728 54324
rect 8300 54204 8352 54256
rect 1584 54179 1636 54188
rect 1584 54145 1593 54179
rect 1593 54145 1627 54179
rect 1627 54145 1636 54179
rect 1584 54136 1636 54145
rect 572 54068 624 54120
rect 2044 54068 2096 54120
rect 9864 54179 9916 54188
rect 2320 54068 2372 54120
rect 1308 54000 1360 54052
rect 9864 54145 9873 54179
rect 9873 54145 9907 54179
rect 9907 54145 9916 54179
rect 9864 54136 9916 54145
rect 10048 54043 10100 54052
rect 10048 54009 10057 54043
rect 10057 54009 10091 54043
rect 10091 54009 10100 54043
rect 10048 54000 10100 54009
rect 1768 53932 1820 53984
rect 2044 53932 2096 53984
rect 2582 53830 2634 53882
rect 2646 53830 2698 53882
rect 2710 53830 2762 53882
rect 2774 53830 2826 53882
rect 2838 53830 2890 53882
rect 5846 53830 5898 53882
rect 5910 53830 5962 53882
rect 5974 53830 6026 53882
rect 6038 53830 6090 53882
rect 6102 53830 6154 53882
rect 9110 53830 9162 53882
rect 9174 53830 9226 53882
rect 9238 53830 9290 53882
rect 9302 53830 9354 53882
rect 9366 53830 9418 53882
rect 2320 53592 2372 53644
rect 2596 53592 2648 53644
rect 4620 53524 4672 53576
rect 9680 53524 9732 53576
rect 5356 53456 5408 53508
rect 1400 53388 1452 53440
rect 2320 53431 2372 53440
rect 2320 53397 2329 53431
rect 2329 53397 2363 53431
rect 2363 53397 2372 53431
rect 2320 53388 2372 53397
rect 10048 53431 10100 53440
rect 10048 53397 10057 53431
rect 10057 53397 10091 53431
rect 10091 53397 10100 53431
rect 10048 53388 10100 53397
rect 4214 53286 4266 53338
rect 4278 53286 4330 53338
rect 4342 53286 4394 53338
rect 4406 53286 4458 53338
rect 4470 53286 4522 53338
rect 7478 53286 7530 53338
rect 7542 53286 7594 53338
rect 7606 53286 7658 53338
rect 7670 53286 7722 53338
rect 7734 53286 7786 53338
rect 2044 53184 2096 53236
rect 2228 53184 2280 53236
rect 4712 53116 4764 53168
rect 6828 53116 6880 53168
rect 664 53048 716 53100
rect 2228 53048 2280 53100
rect 2504 53048 2556 53100
rect 9956 53048 10008 53100
rect 1584 52887 1636 52896
rect 1584 52853 1593 52887
rect 1593 52853 1627 52887
rect 1627 52853 1636 52887
rect 1584 52844 1636 52853
rect 2136 52844 2188 52896
rect 2504 52844 2556 52896
rect 10048 52887 10100 52896
rect 10048 52853 10057 52887
rect 10057 52853 10091 52887
rect 10091 52853 10100 52887
rect 10048 52844 10100 52853
rect 2582 52742 2634 52794
rect 2646 52742 2698 52794
rect 2710 52742 2762 52794
rect 2774 52742 2826 52794
rect 2838 52742 2890 52794
rect 5846 52742 5898 52794
rect 5910 52742 5962 52794
rect 5974 52742 6026 52794
rect 6038 52742 6090 52794
rect 6102 52742 6154 52794
rect 9110 52742 9162 52794
rect 9174 52742 9226 52794
rect 9238 52742 9290 52794
rect 9302 52742 9354 52794
rect 9366 52742 9418 52794
rect 4160 52640 4212 52692
rect 480 52436 532 52488
rect 5356 52504 5408 52556
rect 2320 52479 2372 52488
rect 2320 52445 2329 52479
rect 2329 52445 2363 52479
rect 2363 52445 2372 52479
rect 2320 52436 2372 52445
rect 1492 52300 1544 52352
rect 4214 52198 4266 52250
rect 4278 52198 4330 52250
rect 4342 52198 4394 52250
rect 4406 52198 4458 52250
rect 4470 52198 4522 52250
rect 7478 52198 7530 52250
rect 7542 52198 7594 52250
rect 7606 52198 7658 52250
rect 7670 52198 7722 52250
rect 7734 52198 7786 52250
rect 1584 52096 1636 52148
rect 1400 52003 1452 52012
rect 1400 51969 1409 52003
rect 1409 51969 1443 52003
rect 1443 51969 1452 52003
rect 1400 51960 1452 51969
rect 2872 52096 2924 52148
rect 5356 51960 5408 52012
rect 9864 52003 9916 52012
rect 9864 51969 9873 52003
rect 9873 51969 9907 52003
rect 9907 51969 9916 52003
rect 9864 51960 9916 51969
rect 6920 51892 6972 51944
rect 1676 51756 1728 51808
rect 10048 51799 10100 51808
rect 10048 51765 10057 51799
rect 10057 51765 10091 51799
rect 10091 51765 10100 51799
rect 10048 51756 10100 51765
rect 2582 51654 2634 51706
rect 2646 51654 2698 51706
rect 2710 51654 2762 51706
rect 2774 51654 2826 51706
rect 2838 51654 2890 51706
rect 5846 51654 5898 51706
rect 5910 51654 5962 51706
rect 5974 51654 6026 51706
rect 6038 51654 6090 51706
rect 6102 51654 6154 51706
rect 9110 51654 9162 51706
rect 9174 51654 9226 51706
rect 9238 51654 9290 51706
rect 9302 51654 9354 51706
rect 9366 51654 9418 51706
rect 2320 51552 2372 51604
rect 2964 51595 3016 51604
rect 2964 51561 2973 51595
rect 2973 51561 3007 51595
rect 3007 51561 3016 51595
rect 2964 51552 3016 51561
rect 1308 51484 1360 51536
rect 1676 51484 1728 51536
rect 572 51212 624 51264
rect 1584 51255 1636 51264
rect 112 51076 164 51128
rect 572 51076 624 51128
rect 1584 51221 1593 51255
rect 1593 51221 1627 51255
rect 1627 51221 1636 51255
rect 1584 51212 1636 51221
rect 2596 51348 2648 51400
rect 3608 51416 3660 51468
rect 3148 51391 3200 51400
rect 3148 51357 3157 51391
rect 3157 51357 3191 51391
rect 3191 51357 3200 51391
rect 3148 51348 3200 51357
rect 9680 51348 9732 51400
rect 2780 51280 2832 51332
rect 6644 51212 6696 51264
rect 10048 51255 10100 51264
rect 10048 51221 10057 51255
rect 10057 51221 10091 51255
rect 10091 51221 10100 51255
rect 10048 51212 10100 51221
rect 4214 51110 4266 51162
rect 4278 51110 4330 51162
rect 4342 51110 4394 51162
rect 4406 51110 4458 51162
rect 4470 51110 4522 51162
rect 7478 51110 7530 51162
rect 7542 51110 7594 51162
rect 7606 51110 7658 51162
rect 7670 51110 7722 51162
rect 7734 51110 7786 51162
rect 1124 51008 1176 51060
rect 2136 51008 2188 51060
rect 2320 51008 2372 51060
rect 3148 51008 3200 51060
rect 388 50464 440 50516
rect 5080 51008 5132 51060
rect 5172 51008 5224 51060
rect 9864 51008 9916 51060
rect 1768 50915 1820 50924
rect 1768 50881 1777 50915
rect 1777 50881 1811 50915
rect 1811 50881 1820 50915
rect 1768 50872 1820 50881
rect 2136 50872 2188 50924
rect 1124 50736 1176 50788
rect 1492 50736 1544 50788
rect 4160 50872 4212 50924
rect 4804 50872 4856 50924
rect 5356 50872 5408 50924
rect 2596 50804 2648 50856
rect 2780 50804 2832 50856
rect 4068 50804 4120 50856
rect 4988 50804 5040 50856
rect 5172 50804 5224 50856
rect 5448 50804 5500 50856
rect 6644 50804 6696 50856
rect 1400 50668 1452 50720
rect 6184 50736 6236 50788
rect 2964 50668 3016 50720
rect 2582 50566 2634 50618
rect 2646 50566 2698 50618
rect 2710 50566 2762 50618
rect 2774 50566 2826 50618
rect 2838 50566 2890 50618
rect 5846 50566 5898 50618
rect 5910 50566 5962 50618
rect 5974 50566 6026 50618
rect 6038 50566 6090 50618
rect 6102 50566 6154 50618
rect 9110 50566 9162 50618
rect 9174 50566 9226 50618
rect 9238 50566 9290 50618
rect 9302 50566 9354 50618
rect 9366 50566 9418 50618
rect 1584 50464 1636 50516
rect 1032 50396 1084 50448
rect 2872 50396 2924 50448
rect 4160 50396 4212 50448
rect 112 50328 164 50380
rect 388 50328 440 50380
rect 8484 50328 8536 50380
rect 1584 50303 1636 50312
rect 1584 50269 1593 50303
rect 1593 50269 1627 50303
rect 1627 50269 1636 50303
rect 1584 50260 1636 50269
rect 1768 50303 1820 50312
rect 1768 50269 1777 50303
rect 1777 50269 1811 50303
rect 1811 50269 1820 50303
rect 1768 50260 1820 50269
rect 7104 50260 7156 50312
rect 9864 50303 9916 50312
rect 9864 50269 9873 50303
rect 9873 50269 9907 50303
rect 9907 50269 9916 50303
rect 9864 50260 9916 50269
rect 940 50192 992 50244
rect 1492 50124 1544 50176
rect 2780 50124 2832 50176
rect 10048 50167 10100 50176
rect 10048 50133 10057 50167
rect 10057 50133 10091 50167
rect 10091 50133 10100 50167
rect 10048 50124 10100 50133
rect 4214 50022 4266 50074
rect 4278 50022 4330 50074
rect 4342 50022 4394 50074
rect 4406 50022 4458 50074
rect 4470 50022 4522 50074
rect 7478 50022 7530 50074
rect 7542 50022 7594 50074
rect 7606 50022 7658 50074
rect 7670 50022 7722 50074
rect 7734 50022 7786 50074
rect 9588 49920 9640 49972
rect 1676 49895 1728 49904
rect 1676 49861 1685 49895
rect 1685 49861 1719 49895
rect 1719 49861 1728 49895
rect 1676 49852 1728 49861
rect 1124 49784 1176 49836
rect 1584 49827 1636 49836
rect 1584 49793 1593 49827
rect 1593 49793 1627 49827
rect 1627 49793 1636 49827
rect 1584 49784 1636 49793
rect 1768 49827 1820 49836
rect 1768 49793 1777 49827
rect 1777 49793 1811 49827
rect 1811 49793 1820 49827
rect 1768 49784 1820 49793
rect 2504 49784 2556 49836
rect 9956 49784 10008 49836
rect 1768 49648 1820 49700
rect 2596 49716 2648 49768
rect 3792 49716 3844 49768
rect 3976 49716 4028 49768
rect 1124 49580 1176 49632
rect 2504 49580 2556 49632
rect 3424 49580 3476 49632
rect 3976 49580 4028 49632
rect 2582 49478 2634 49530
rect 2646 49478 2698 49530
rect 2710 49478 2762 49530
rect 2774 49478 2826 49530
rect 2838 49478 2890 49530
rect 5846 49478 5898 49530
rect 5910 49478 5962 49530
rect 5974 49478 6026 49530
rect 6038 49478 6090 49530
rect 6102 49478 6154 49530
rect 9110 49478 9162 49530
rect 9174 49478 9226 49530
rect 9238 49478 9290 49530
rect 9302 49478 9354 49530
rect 9366 49478 9418 49530
rect 20 49376 72 49428
rect 2412 49376 2464 49428
rect 3516 49376 3568 49428
rect 3884 49376 3936 49428
rect 9680 49376 9732 49428
rect 1400 49308 1452 49360
rect 1676 49308 1728 49360
rect 2688 49308 2740 49360
rect 4528 49308 4580 49360
rect 2872 49240 2924 49292
rect 6552 49172 6604 49224
rect 9496 49172 9548 49224
rect 6736 49104 6788 49156
rect 1400 49036 1452 49088
rect 2320 49079 2372 49088
rect 2320 49045 2329 49079
rect 2329 49045 2363 49079
rect 2363 49045 2372 49079
rect 2320 49036 2372 49045
rect 10048 49079 10100 49088
rect 10048 49045 10057 49079
rect 10057 49045 10091 49079
rect 10091 49045 10100 49079
rect 10048 49036 10100 49045
rect 4214 48934 4266 48986
rect 4278 48934 4330 48986
rect 4342 48934 4394 48986
rect 4406 48934 4458 48986
rect 4470 48934 4522 48986
rect 7478 48934 7530 48986
rect 7542 48934 7594 48986
rect 7606 48934 7658 48986
rect 7670 48934 7722 48986
rect 7734 48934 7786 48986
rect 9864 48832 9916 48884
rect 2688 48764 2740 48816
rect 2964 48764 3016 48816
rect 2780 48696 2832 48748
rect 3148 48696 3200 48748
rect 2964 48628 3016 48680
rect 1124 48492 1176 48544
rect 1584 48535 1636 48544
rect 1584 48501 1593 48535
rect 1593 48501 1627 48535
rect 1627 48501 1636 48535
rect 1584 48492 1636 48501
rect 10140 48739 10192 48748
rect 10140 48705 10149 48739
rect 10149 48705 10183 48739
rect 10183 48705 10192 48739
rect 10140 48696 10192 48705
rect 3516 48492 3568 48544
rect 6552 48492 6604 48544
rect 2582 48390 2634 48442
rect 2646 48390 2698 48442
rect 2710 48390 2762 48442
rect 2774 48390 2826 48442
rect 2838 48390 2890 48442
rect 5846 48390 5898 48442
rect 5910 48390 5962 48442
rect 5974 48390 6026 48442
rect 6038 48390 6090 48442
rect 6102 48390 6154 48442
rect 9110 48390 9162 48442
rect 9174 48390 9226 48442
rect 9238 48390 9290 48442
rect 9302 48390 9354 48442
rect 9366 48390 9418 48442
rect 1768 48288 1820 48340
rect 2688 48274 2740 48326
rect 4528 48288 4580 48340
rect 2780 48263 2832 48272
rect 2780 48229 2789 48263
rect 2789 48229 2823 48263
rect 2823 48229 2832 48263
rect 2780 48220 2832 48229
rect 6184 48220 6236 48272
rect 7196 48220 7248 48272
rect 9496 48220 9548 48272
rect 1400 48127 1452 48136
rect 1400 48093 1409 48127
rect 1409 48093 1443 48127
rect 1443 48093 1452 48127
rect 1400 48084 1452 48093
rect 2412 48127 2464 48136
rect 2412 48093 2421 48127
rect 2421 48093 2455 48127
rect 2455 48093 2464 48127
rect 2412 48084 2464 48093
rect 2596 48127 2648 48136
rect 2596 48093 2605 48127
rect 2605 48093 2639 48127
rect 2639 48093 2648 48127
rect 2596 48084 2648 48093
rect 2964 48016 3016 48068
rect 1584 47991 1636 48000
rect 1584 47957 1593 47991
rect 1593 47957 1627 47991
rect 1627 47957 1636 47991
rect 1584 47948 1636 47957
rect 4528 48016 4580 48068
rect 6184 48016 6236 48068
rect 10048 47991 10100 48000
rect 10048 47957 10057 47991
rect 10057 47957 10091 47991
rect 10091 47957 10100 47991
rect 10048 47948 10100 47957
rect 4214 47846 4266 47898
rect 4278 47846 4330 47898
rect 4342 47846 4394 47898
rect 4406 47846 4458 47898
rect 4470 47846 4522 47898
rect 7478 47846 7530 47898
rect 7542 47846 7594 47898
rect 7606 47846 7658 47898
rect 7670 47846 7722 47898
rect 7734 47846 7786 47898
rect 3516 47744 3568 47796
rect 2596 47676 2648 47728
rect 3884 47676 3936 47728
rect 2412 47540 2464 47592
rect 3148 47540 3200 47592
rect 3424 47540 3476 47592
rect 7472 47608 7524 47660
rect 3884 47540 3936 47592
rect 1492 47404 1544 47456
rect 3700 47447 3752 47456
rect 3700 47413 3709 47447
rect 3709 47413 3743 47447
rect 3743 47413 3752 47447
rect 3700 47404 3752 47413
rect 10048 47447 10100 47456
rect 10048 47413 10057 47447
rect 10057 47413 10091 47447
rect 10091 47413 10100 47447
rect 10048 47404 10100 47413
rect 2582 47302 2634 47354
rect 2646 47302 2698 47354
rect 2710 47302 2762 47354
rect 2774 47302 2826 47354
rect 2838 47302 2890 47354
rect 5846 47302 5898 47354
rect 5910 47302 5962 47354
rect 5974 47302 6026 47354
rect 6038 47302 6090 47354
rect 6102 47302 6154 47354
rect 9110 47302 9162 47354
rect 9174 47302 9226 47354
rect 9238 47302 9290 47354
rect 9302 47302 9354 47354
rect 9366 47302 9418 47354
rect 2412 47200 2464 47252
rect 1492 47107 1544 47116
rect 1492 47073 1501 47107
rect 1501 47073 1535 47107
rect 1535 47073 1544 47107
rect 1492 47064 1544 47073
rect 1768 47107 1820 47116
rect 1768 47073 1777 47107
rect 1777 47073 1811 47107
rect 1811 47073 1820 47107
rect 1768 47064 1820 47073
rect 2412 47064 2464 47116
rect 7288 47200 7340 47252
rect 7472 47243 7524 47252
rect 7472 47209 7481 47243
rect 7481 47209 7515 47243
rect 7515 47209 7524 47243
rect 7472 47200 7524 47209
rect 9956 47243 10008 47252
rect 9956 47209 9965 47243
rect 9965 47209 9999 47243
rect 9999 47209 10008 47243
rect 9956 47200 10008 47209
rect 4620 47132 4672 47184
rect 5172 47132 5224 47184
rect 1492 46928 1544 46980
rect 1676 46928 1728 46980
rect 4528 46996 4580 47048
rect 5816 47064 5868 47116
rect 6184 47064 6236 47116
rect 3976 46903 4028 46912
rect 3976 46869 3985 46903
rect 3985 46869 4019 46903
rect 4019 46869 4028 46903
rect 3976 46860 4028 46869
rect 5172 46860 5224 46912
rect 4214 46758 4266 46810
rect 4278 46758 4330 46810
rect 4342 46758 4394 46810
rect 4406 46758 4458 46810
rect 4470 46758 4522 46810
rect 7478 46758 7530 46810
rect 7542 46758 7594 46810
rect 7606 46758 7658 46810
rect 7670 46758 7722 46810
rect 7734 46758 7786 46810
rect 112 46656 164 46708
rect 1400 46656 1452 46708
rect 1768 46656 1820 46708
rect 1952 46656 2004 46708
rect 10140 46656 10192 46708
rect 112 46520 164 46572
rect 2412 46520 2464 46572
rect 3700 46563 3752 46572
rect 3700 46529 3709 46563
rect 3709 46529 3743 46563
rect 3743 46529 3752 46563
rect 3700 46520 3752 46529
rect 5724 46520 5776 46572
rect 6552 46520 6604 46572
rect 7012 46520 7064 46572
rect 3332 46452 3384 46504
rect 4160 46452 4212 46504
rect 5632 46452 5684 46504
rect 6184 46452 6236 46504
rect 3884 46427 3936 46436
rect 3884 46393 3893 46427
rect 3893 46393 3927 46427
rect 3927 46393 3936 46427
rect 3884 46384 3936 46393
rect 10048 46427 10100 46436
rect 10048 46393 10057 46427
rect 10057 46393 10091 46427
rect 10091 46393 10100 46427
rect 10048 46384 10100 46393
rect 1400 46316 1452 46368
rect 4988 46316 5040 46368
rect 6644 46316 6696 46368
rect 2582 46214 2634 46266
rect 2646 46214 2698 46266
rect 2710 46214 2762 46266
rect 2774 46214 2826 46266
rect 2838 46214 2890 46266
rect 5846 46214 5898 46266
rect 5910 46214 5962 46266
rect 5974 46214 6026 46266
rect 6038 46214 6090 46266
rect 6102 46214 6154 46266
rect 9110 46214 9162 46266
rect 9174 46214 9226 46266
rect 9238 46214 9290 46266
rect 9302 46214 9354 46266
rect 9366 46214 9418 46266
rect 3056 46044 3108 46096
rect 3240 46044 3292 46096
rect 4528 46044 4580 46096
rect 4712 46044 4764 46096
rect 1400 46019 1452 46028
rect 1400 45985 1409 46019
rect 1409 45985 1443 46019
rect 1443 45985 1452 46019
rect 1400 45976 1452 45985
rect 1676 46019 1728 46028
rect 1676 45985 1685 46019
rect 1685 45985 1719 46019
rect 1719 45985 1728 46019
rect 1676 45976 1728 45985
rect 2688 45951 2740 45960
rect 2688 45917 2697 45951
rect 2697 45917 2731 45951
rect 2731 45917 2740 45951
rect 2688 45908 2740 45917
rect 3792 45951 3844 45960
rect 3792 45917 3801 45951
rect 3801 45917 3835 45951
rect 3835 45917 3844 45951
rect 3792 45908 3844 45917
rect 9864 45951 9916 45960
rect 9864 45917 9873 45951
rect 9873 45917 9907 45951
rect 9907 45917 9916 45951
rect 9864 45908 9916 45917
rect 3056 45840 3108 45892
rect 4160 45840 4212 45892
rect 2872 45815 2924 45824
rect 2872 45781 2881 45815
rect 2881 45781 2915 45815
rect 2915 45781 2924 45815
rect 2872 45772 2924 45781
rect 3976 45815 4028 45824
rect 3976 45781 3985 45815
rect 3985 45781 4019 45815
rect 4019 45781 4028 45815
rect 3976 45772 4028 45781
rect 5540 45772 5592 45824
rect 5724 45772 5776 45824
rect 10048 45815 10100 45824
rect 10048 45781 10057 45815
rect 10057 45781 10091 45815
rect 10091 45781 10100 45815
rect 10048 45772 10100 45781
rect 4214 45670 4266 45722
rect 4278 45670 4330 45722
rect 4342 45670 4394 45722
rect 4406 45670 4458 45722
rect 4470 45670 4522 45722
rect 7478 45670 7530 45722
rect 7542 45670 7594 45722
rect 7606 45670 7658 45722
rect 7670 45670 7722 45722
rect 7734 45670 7786 45722
rect 572 45568 624 45620
rect 1032 45568 1084 45620
rect 296 45432 348 45484
rect 1032 45432 1084 45484
rect 1492 45432 1544 45484
rect 2872 45500 2924 45552
rect 3792 45500 3844 45552
rect 572 45364 624 45416
rect 1860 45407 1912 45416
rect 1860 45373 1869 45407
rect 1869 45373 1903 45407
rect 1903 45373 1912 45407
rect 1860 45364 1912 45373
rect 20 45228 72 45280
rect 112 45228 164 45280
rect 296 45228 348 45280
rect 2582 45126 2634 45178
rect 2646 45126 2698 45178
rect 2710 45126 2762 45178
rect 2774 45126 2826 45178
rect 2838 45126 2890 45178
rect 5846 45126 5898 45178
rect 5910 45126 5962 45178
rect 5974 45126 6026 45178
rect 6038 45126 6090 45178
rect 6102 45126 6154 45178
rect 9110 45126 9162 45178
rect 9174 45126 9226 45178
rect 9238 45126 9290 45178
rect 9302 45126 9354 45178
rect 9366 45126 9418 45178
rect 112 45024 164 45076
rect 1308 45024 1360 45076
rect 1584 45067 1636 45076
rect 1584 45033 1593 45067
rect 1593 45033 1627 45067
rect 1627 45033 1636 45067
rect 1584 45024 1636 45033
rect 1860 45024 1912 45076
rect 7012 45024 7064 45076
rect 1400 44863 1452 44872
rect 1400 44829 1409 44863
rect 1409 44829 1443 44863
rect 1443 44829 1452 44863
rect 1400 44820 1452 44829
rect 2412 44820 2464 44872
rect 2596 44820 2648 44872
rect 4896 44820 4948 44872
rect 8300 44820 8352 44872
rect 3976 44752 4028 44804
rect 1860 44684 1912 44736
rect 3884 44684 3936 44736
rect 10048 44727 10100 44736
rect 10048 44693 10057 44727
rect 10057 44693 10091 44727
rect 10091 44693 10100 44727
rect 10048 44684 10100 44693
rect 4214 44582 4266 44634
rect 4278 44582 4330 44634
rect 4342 44582 4394 44634
rect 4406 44582 4458 44634
rect 4470 44582 4522 44634
rect 7478 44582 7530 44634
rect 7542 44582 7594 44634
rect 7606 44582 7658 44634
rect 7670 44582 7722 44634
rect 7734 44582 7786 44634
rect 1584 44523 1636 44532
rect 1584 44489 1593 44523
rect 1593 44489 1627 44523
rect 1627 44489 1636 44523
rect 1584 44480 1636 44489
rect 3056 44480 3108 44532
rect 4896 44523 4948 44532
rect 4896 44489 4905 44523
rect 4905 44489 4939 44523
rect 4939 44489 4948 44523
rect 4896 44480 4948 44489
rect 296 44276 348 44328
rect 3792 44344 3844 44396
rect 4252 44344 4304 44396
rect 4896 44344 4948 44396
rect 5632 44344 5684 44396
rect 9496 44344 9548 44396
rect 3884 44276 3936 44328
rect 3976 44276 4028 44328
rect 2964 44208 3016 44260
rect 5172 44208 5224 44260
rect 3792 44183 3844 44192
rect 3792 44149 3801 44183
rect 3801 44149 3835 44183
rect 3835 44149 3844 44183
rect 3792 44140 3844 44149
rect 10048 44183 10100 44192
rect 10048 44149 10057 44183
rect 10057 44149 10091 44183
rect 10091 44149 10100 44183
rect 10048 44140 10100 44149
rect 2582 44038 2634 44090
rect 2646 44038 2698 44090
rect 2710 44038 2762 44090
rect 2774 44038 2826 44090
rect 2838 44038 2890 44090
rect 5846 44038 5898 44090
rect 5910 44038 5962 44090
rect 5974 44038 6026 44090
rect 6038 44038 6090 44090
rect 6102 44038 6154 44090
rect 9110 44038 9162 44090
rect 9174 44038 9226 44090
rect 9238 44038 9290 44090
rect 9302 44038 9354 44090
rect 9366 44038 9418 44090
rect 2228 43868 2280 43920
rect 9496 43936 9548 43988
rect 1492 43664 1544 43716
rect 2136 43800 2188 43852
rect 2872 43800 2924 43852
rect 3148 43800 3200 43852
rect 2504 43732 2556 43784
rect 3424 43732 3476 43784
rect 3884 43775 3936 43784
rect 3884 43741 3893 43775
rect 3893 43741 3927 43775
rect 3927 43741 3936 43775
rect 3884 43732 3936 43741
rect 4252 43732 4304 43784
rect 9772 43868 9824 43920
rect 2780 43664 2832 43716
rect 9956 43732 10008 43784
rect 2228 43596 2280 43648
rect 2964 43596 3016 43648
rect 3148 43639 3200 43648
rect 3148 43605 3157 43639
rect 3157 43605 3191 43639
rect 3191 43605 3200 43639
rect 3148 43596 3200 43605
rect 3424 43596 3476 43648
rect 10048 43639 10100 43648
rect 10048 43605 10057 43639
rect 10057 43605 10091 43639
rect 10091 43605 10100 43639
rect 10048 43596 10100 43605
rect 4214 43494 4266 43546
rect 4278 43494 4330 43546
rect 4342 43494 4394 43546
rect 4406 43494 4458 43546
rect 4470 43494 4522 43546
rect 7478 43494 7530 43546
rect 7542 43494 7594 43546
rect 7606 43494 7658 43546
rect 7670 43494 7722 43546
rect 7734 43494 7786 43546
rect 1584 43435 1636 43444
rect 1584 43401 1593 43435
rect 1593 43401 1627 43435
rect 1627 43401 1636 43435
rect 1584 43392 1636 43401
rect 9956 43435 10008 43444
rect 9956 43401 9965 43435
rect 9965 43401 9999 43435
rect 9999 43401 10008 43435
rect 9956 43392 10008 43401
rect 1492 43256 1544 43308
rect 2504 43256 2556 43308
rect 2688 43256 2740 43308
rect 1308 43188 1360 43240
rect 1676 43188 1728 43240
rect 2412 43188 2464 43240
rect 2780 43188 2832 43240
rect 3424 43188 3476 43240
rect 10140 43299 10192 43308
rect 10140 43265 10149 43299
rect 10149 43265 10183 43299
rect 10183 43265 10192 43299
rect 10140 43256 10192 43265
rect 4160 43188 4212 43240
rect 1492 43120 1544 43172
rect 3792 43120 3844 43172
rect 3056 43052 3108 43104
rect 3976 43095 4028 43104
rect 3976 43061 3985 43095
rect 3985 43061 4019 43095
rect 4019 43061 4028 43095
rect 3976 43052 4028 43061
rect 2582 42950 2634 43002
rect 2646 42950 2698 43002
rect 2710 42950 2762 43002
rect 2774 42950 2826 43002
rect 2838 42950 2890 43002
rect 5846 42950 5898 43002
rect 5910 42950 5962 43002
rect 5974 42950 6026 43002
rect 6038 42950 6090 43002
rect 6102 42950 6154 43002
rect 9110 42950 9162 43002
rect 9174 42950 9226 43002
rect 9238 42950 9290 43002
rect 9302 42950 9354 43002
rect 9366 42950 9418 43002
rect 572 42780 624 42832
rect 3148 42712 3200 42764
rect 3516 42712 3568 42764
rect 1492 42687 1544 42696
rect 1492 42653 1501 42687
rect 1501 42653 1535 42687
rect 1535 42653 1544 42687
rect 1492 42644 1544 42653
rect 2964 42644 3016 42696
rect 3792 42687 3844 42696
rect 3792 42653 3801 42687
rect 3801 42653 3835 42687
rect 3835 42653 3844 42687
rect 3792 42644 3844 42653
rect 9772 42644 9824 42696
rect 2964 42551 3016 42560
rect 2964 42517 2973 42551
rect 2973 42517 3007 42551
rect 3007 42517 3016 42551
rect 2964 42508 3016 42517
rect 3424 42508 3476 42560
rect 10048 42551 10100 42560
rect 10048 42517 10057 42551
rect 10057 42517 10091 42551
rect 10091 42517 10100 42551
rect 10048 42508 10100 42517
rect 4214 42406 4266 42458
rect 4278 42406 4330 42458
rect 4342 42406 4394 42458
rect 4406 42406 4458 42458
rect 4470 42406 4522 42458
rect 7478 42406 7530 42458
rect 7542 42406 7594 42458
rect 7606 42406 7658 42458
rect 7670 42406 7722 42458
rect 7734 42406 7786 42458
rect 1492 42304 1544 42356
rect 10140 42304 10192 42356
rect 1308 42236 1360 42288
rect 1768 42236 1820 42288
rect 2688 42236 2740 42288
rect 2780 42168 2832 42220
rect 3976 42211 4028 42220
rect 1400 42143 1452 42152
rect 1400 42109 1409 42143
rect 1409 42109 1443 42143
rect 1443 42109 1452 42143
rect 1400 42100 1452 42109
rect 2228 42100 2280 42152
rect 572 42032 624 42084
rect 2228 41964 2280 42016
rect 3976 42177 3985 42211
rect 3985 42177 4019 42211
rect 4019 42177 4028 42211
rect 3976 42168 4028 42177
rect 4436 42236 4488 42288
rect 4896 42236 4948 42288
rect 5264 42168 5316 42220
rect 5632 42211 5684 42220
rect 5632 42177 5641 42211
rect 5641 42177 5675 42211
rect 5675 42177 5684 42211
rect 5632 42168 5684 42177
rect 9496 42168 9548 42220
rect 3792 42032 3844 42084
rect 8300 42032 8352 42084
rect 10048 42007 10100 42016
rect 10048 41973 10057 42007
rect 10057 41973 10091 42007
rect 10091 41973 10100 42007
rect 10048 41964 10100 41973
rect 2582 41862 2634 41914
rect 2646 41862 2698 41914
rect 2710 41862 2762 41914
rect 2774 41862 2826 41914
rect 2838 41862 2890 41914
rect 5846 41862 5898 41914
rect 5910 41862 5962 41914
rect 5974 41862 6026 41914
rect 6038 41862 6090 41914
rect 6102 41862 6154 41914
rect 9110 41862 9162 41914
rect 9174 41862 9226 41914
rect 9238 41862 9290 41914
rect 9302 41862 9354 41914
rect 9366 41862 9418 41914
rect 5632 41760 5684 41812
rect 2780 41692 2832 41744
rect 4160 41624 4212 41676
rect 5264 41624 5316 41676
rect 1308 41556 1360 41608
rect 3424 41556 3476 41608
rect 4068 41556 4120 41608
rect 4436 41599 4488 41608
rect 4436 41565 4445 41599
rect 4445 41565 4479 41599
rect 4479 41565 4488 41599
rect 4436 41556 4488 41565
rect 5080 41556 5132 41608
rect 1032 41488 1084 41540
rect 1952 41488 2004 41540
rect 2688 41488 2740 41540
rect 3792 41488 3844 41540
rect 1768 41420 1820 41472
rect 3516 41420 3568 41472
rect 4214 41318 4266 41370
rect 4278 41318 4330 41370
rect 4342 41318 4394 41370
rect 4406 41318 4458 41370
rect 4470 41318 4522 41370
rect 7478 41318 7530 41370
rect 7542 41318 7594 41370
rect 7606 41318 7658 41370
rect 7670 41318 7722 41370
rect 7734 41318 7786 41370
rect 1400 41216 1452 41268
rect 2412 41216 2464 41268
rect 2596 41216 2648 41268
rect 2780 41259 2832 41268
rect 2780 41225 2789 41259
rect 2789 41225 2823 41259
rect 2823 41225 2832 41259
rect 2780 41216 2832 41225
rect 3516 41216 3568 41268
rect 6184 41216 6236 41268
rect 1124 41148 1176 41200
rect 1676 41148 1728 41200
rect 3884 41148 3936 41200
rect 4344 41148 4396 41200
rect 1400 41080 1452 41132
rect 1952 41080 2004 41132
rect 2228 41080 2280 41132
rect 2688 41080 2740 41132
rect 4528 41123 4580 41132
rect 4528 41089 4537 41123
rect 4537 41089 4571 41123
rect 4571 41089 4580 41123
rect 4528 41080 4580 41089
rect 6184 41080 6236 41132
rect 5080 41012 5132 41064
rect 5356 41012 5408 41064
rect 5632 41012 5684 41064
rect 4068 40944 4120 40996
rect 9864 40944 9916 40996
rect 10048 40987 10100 40996
rect 10048 40953 10057 40987
rect 10057 40953 10091 40987
rect 10091 40953 10100 40987
rect 10048 40944 10100 40953
rect 3424 40919 3476 40928
rect 3424 40885 3433 40919
rect 3433 40885 3467 40919
rect 3467 40885 3476 40919
rect 3424 40876 3476 40885
rect 5080 40876 5132 40928
rect 7288 40876 7340 40928
rect 2582 40774 2634 40826
rect 2646 40774 2698 40826
rect 2710 40774 2762 40826
rect 2774 40774 2826 40826
rect 2838 40774 2890 40826
rect 5846 40774 5898 40826
rect 5910 40774 5962 40826
rect 5974 40774 6026 40826
rect 6038 40774 6090 40826
rect 6102 40774 6154 40826
rect 9110 40774 9162 40826
rect 9174 40774 9226 40826
rect 9238 40774 9290 40826
rect 9302 40774 9354 40826
rect 9366 40774 9418 40826
rect 3792 40672 3844 40724
rect 4068 40672 4120 40724
rect 9496 40672 9548 40724
rect 2228 40604 2280 40656
rect 3976 40604 4028 40656
rect 4712 40604 4764 40656
rect 5632 40604 5684 40656
rect 20 40536 72 40588
rect 20 40400 72 40452
rect 572 40400 624 40452
rect 4344 40468 4396 40520
rect 4988 40468 5040 40520
rect 9864 40511 9916 40520
rect 9864 40477 9873 40511
rect 9873 40477 9907 40511
rect 9907 40477 9916 40511
rect 9864 40468 9916 40477
rect 4528 40400 4580 40452
rect 4712 40400 4764 40452
rect 3148 40332 3200 40384
rect 3240 40332 3292 40384
rect 3424 40332 3476 40384
rect 3976 40375 4028 40384
rect 3976 40341 3985 40375
rect 3985 40341 4019 40375
rect 4019 40341 4028 40375
rect 3976 40332 4028 40341
rect 10048 40375 10100 40384
rect 10048 40341 10057 40375
rect 10057 40341 10091 40375
rect 10091 40341 10100 40375
rect 10048 40332 10100 40341
rect 4214 40230 4266 40282
rect 4278 40230 4330 40282
rect 4342 40230 4394 40282
rect 4406 40230 4458 40282
rect 4470 40230 4522 40282
rect 7478 40230 7530 40282
rect 7542 40230 7594 40282
rect 7606 40230 7658 40282
rect 7670 40230 7722 40282
rect 7734 40230 7786 40282
rect 2228 40128 2280 40180
rect 1952 40060 2004 40112
rect 2964 40060 3016 40112
rect 4344 40060 4396 40112
rect 4712 40060 4764 40112
rect 9864 40128 9916 40180
rect 6644 40060 6696 40112
rect 5724 39992 5776 40044
rect 6552 40035 6604 40044
rect 6552 40001 6561 40035
rect 6561 40001 6595 40035
rect 6595 40001 6604 40035
rect 6552 39992 6604 40001
rect 9864 40035 9916 40044
rect 9864 40001 9873 40035
rect 9873 40001 9907 40035
rect 9907 40001 9916 40035
rect 9864 39992 9916 40001
rect 2596 39924 2648 39976
rect 3332 39856 3384 39908
rect 4252 39788 4304 39840
rect 10048 39831 10100 39840
rect 10048 39797 10057 39831
rect 10057 39797 10091 39831
rect 10091 39797 10100 39831
rect 10048 39788 10100 39797
rect 2582 39686 2634 39738
rect 2646 39686 2698 39738
rect 2710 39686 2762 39738
rect 2774 39686 2826 39738
rect 2838 39686 2890 39738
rect 5846 39686 5898 39738
rect 5910 39686 5962 39738
rect 5974 39686 6026 39738
rect 6038 39686 6090 39738
rect 6102 39686 6154 39738
rect 9110 39686 9162 39738
rect 9174 39686 9226 39738
rect 9238 39686 9290 39738
rect 9302 39686 9354 39738
rect 9366 39686 9418 39738
rect 3148 39627 3200 39636
rect 3148 39593 3157 39627
rect 3157 39593 3191 39627
rect 3191 39593 3200 39627
rect 3148 39584 3200 39593
rect 6184 39584 6236 39636
rect 9772 39584 9824 39636
rect 2228 39516 2280 39568
rect 3332 39516 3384 39568
rect 3792 39516 3844 39568
rect 5724 39448 5776 39500
rect 1124 39380 1176 39432
rect 2780 39423 2832 39432
rect 2780 39389 2789 39423
rect 2789 39389 2823 39423
rect 2823 39389 2832 39423
rect 2780 39380 2832 39389
rect 2964 39423 3016 39432
rect 2964 39389 2973 39423
rect 2973 39389 3007 39423
rect 3007 39389 3016 39423
rect 2964 39380 3016 39389
rect 2504 39312 2556 39364
rect 4344 39380 4396 39432
rect 4620 39423 4672 39432
rect 4620 39389 4629 39423
rect 4629 39389 4663 39423
rect 4663 39389 4672 39423
rect 4620 39380 4672 39389
rect 5540 39423 5592 39432
rect 5540 39389 5549 39423
rect 5549 39389 5583 39423
rect 5583 39389 5592 39423
rect 5540 39380 5592 39389
rect 4214 39142 4266 39194
rect 4278 39142 4330 39194
rect 4342 39142 4394 39194
rect 4406 39142 4458 39194
rect 4470 39142 4522 39194
rect 7478 39142 7530 39194
rect 7542 39142 7594 39194
rect 7606 39142 7658 39194
rect 7670 39142 7722 39194
rect 7734 39142 7786 39194
rect 1124 39040 1176 39092
rect 1768 39040 1820 39092
rect 1952 39040 2004 39092
rect 6552 39040 6604 39092
rect 3240 38972 3292 39024
rect 3792 38972 3844 39024
rect 5632 38972 5684 39024
rect 940 38904 992 38956
rect 4436 38904 4488 38956
rect 5724 38904 5776 38956
rect 9680 38904 9732 38956
rect 1676 38836 1728 38888
rect 2964 38836 3016 38888
rect 3056 38768 3108 38820
rect 4160 38836 4212 38888
rect 4252 38768 4304 38820
rect 10048 38743 10100 38752
rect 10048 38709 10057 38743
rect 10057 38709 10091 38743
rect 10091 38709 10100 38743
rect 10048 38700 10100 38709
rect 2582 38598 2634 38650
rect 2646 38598 2698 38650
rect 2710 38598 2762 38650
rect 2774 38598 2826 38650
rect 2838 38598 2890 38650
rect 5846 38598 5898 38650
rect 5910 38598 5962 38650
rect 5974 38598 6026 38650
rect 6038 38598 6090 38650
rect 6102 38598 6154 38650
rect 9110 38598 9162 38650
rect 9174 38598 9226 38650
rect 9238 38598 9290 38650
rect 9302 38598 9354 38650
rect 9366 38598 9418 38650
rect 572 38496 624 38548
rect 1400 38496 1452 38548
rect 1492 38496 1544 38548
rect 1676 38496 1728 38548
rect 1768 38496 1820 38548
rect 940 38360 992 38412
rect 1308 38360 1360 38412
rect 1124 38292 1176 38344
rect 1676 38360 1728 38412
rect 1952 38496 2004 38548
rect 2044 38496 2096 38548
rect 2136 38496 2188 38548
rect 2228 38496 2280 38548
rect 2964 38496 3016 38548
rect 1952 38360 2004 38412
rect 1768 38292 1820 38344
rect 1860 38224 1912 38276
rect 2136 38224 2188 38276
rect 3148 38496 3200 38548
rect 5540 38496 5592 38548
rect 3056 38428 3108 38480
rect 4252 38428 4304 38480
rect 2504 38292 2556 38344
rect 4436 38335 4488 38344
rect 2320 38224 2372 38276
rect 2964 38224 3016 38276
rect 4160 38224 4212 38276
rect 940 38156 992 38208
rect 2044 38156 2096 38208
rect 2228 38156 2280 38208
rect 2688 38156 2740 38208
rect 4436 38301 4445 38335
rect 4445 38301 4479 38335
rect 4479 38301 4488 38335
rect 4436 38292 4488 38301
rect 5540 38292 5592 38344
rect 9956 38292 10008 38344
rect 10048 38199 10100 38208
rect 10048 38165 10057 38199
rect 10057 38165 10091 38199
rect 10091 38165 10100 38199
rect 10048 38156 10100 38165
rect 4214 38054 4266 38106
rect 4278 38054 4330 38106
rect 4342 38054 4394 38106
rect 4406 38054 4458 38106
rect 4470 38054 4522 38106
rect 7478 38054 7530 38106
rect 7542 38054 7594 38106
rect 7606 38054 7658 38106
rect 7670 38054 7722 38106
rect 7734 38054 7786 38106
rect 1124 37952 1176 38004
rect 1676 37952 1728 38004
rect 2780 37995 2832 38004
rect 2780 37961 2789 37995
rect 2789 37961 2823 37995
rect 2823 37961 2832 37995
rect 2780 37952 2832 37961
rect 9864 37952 9916 38004
rect 1216 37884 1268 37936
rect 2964 37884 3016 37936
rect 2596 37859 2648 37868
rect 1400 37748 1452 37800
rect 2596 37825 2605 37859
rect 2605 37825 2639 37859
rect 2639 37825 2648 37859
rect 2596 37816 2648 37825
rect 3792 37816 3844 37868
rect 6736 37816 6788 37868
rect 10232 37816 10284 37868
rect 1952 37748 2004 37800
rect 2320 37748 2372 37800
rect 1676 37680 1728 37732
rect 2688 37748 2740 37800
rect 3516 37680 3568 37732
rect 20 37612 72 37664
rect 1952 37612 2004 37664
rect 3424 37655 3476 37664
rect 3424 37621 3433 37655
rect 3433 37621 3467 37655
rect 3467 37621 3476 37655
rect 3424 37612 3476 37621
rect 2582 37510 2634 37562
rect 2646 37510 2698 37562
rect 2710 37510 2762 37562
rect 2774 37510 2826 37562
rect 2838 37510 2890 37562
rect 5846 37510 5898 37562
rect 5910 37510 5962 37562
rect 5974 37510 6026 37562
rect 6038 37510 6090 37562
rect 6102 37510 6154 37562
rect 9110 37510 9162 37562
rect 9174 37510 9226 37562
rect 9238 37510 9290 37562
rect 9302 37510 9354 37562
rect 9366 37510 9418 37562
rect 1492 37408 1544 37460
rect 2228 37408 2280 37460
rect 2504 37408 2556 37460
rect 572 37340 624 37392
rect 1676 37272 1728 37324
rect 1860 37340 1912 37392
rect 1492 37204 1544 37256
rect 5632 37272 5684 37324
rect 7104 37272 7156 37324
rect 3700 37204 3752 37256
rect 9864 37247 9916 37256
rect 9864 37213 9873 37247
rect 9873 37213 9907 37247
rect 9907 37213 9916 37247
rect 9864 37204 9916 37213
rect 2228 37136 2280 37188
rect 2320 37136 2372 37188
rect 2688 37179 2740 37188
rect 2688 37145 2697 37179
rect 2697 37145 2731 37179
rect 2731 37145 2740 37179
rect 2688 37136 2740 37145
rect 1584 37111 1636 37120
rect 1584 37077 1593 37111
rect 1593 37077 1627 37111
rect 1627 37077 1636 37111
rect 1584 37068 1636 37077
rect 2964 37068 3016 37120
rect 3700 37068 3752 37120
rect 10048 37111 10100 37120
rect 10048 37077 10057 37111
rect 10057 37077 10091 37111
rect 10091 37077 10100 37111
rect 10048 37068 10100 37077
rect 4214 36966 4266 37018
rect 4278 36966 4330 37018
rect 4342 36966 4394 37018
rect 4406 36966 4458 37018
rect 4470 36966 4522 37018
rect 7478 36966 7530 37018
rect 7542 36966 7594 37018
rect 7606 36966 7658 37018
rect 7670 36966 7722 37018
rect 7734 36966 7786 37018
rect 1124 36864 1176 36916
rect 2320 36864 2372 36916
rect 2688 36864 2740 36916
rect 2872 36796 2924 36848
rect 4988 36864 5040 36916
rect 2504 36728 2556 36780
rect 4528 36796 4580 36848
rect 5540 36728 5592 36780
rect 5724 36728 5776 36780
rect 10140 36728 10192 36780
rect 1124 36660 1176 36712
rect 1860 36660 1912 36712
rect 3424 36635 3476 36644
rect 3424 36601 3433 36635
rect 3433 36601 3467 36635
rect 3467 36601 3476 36635
rect 3424 36592 3476 36601
rect 2504 36524 2556 36576
rect 3056 36524 3108 36576
rect 3332 36524 3384 36576
rect 10048 36567 10100 36576
rect 10048 36533 10057 36567
rect 10057 36533 10091 36567
rect 10091 36533 10100 36567
rect 10048 36524 10100 36533
rect 2582 36422 2634 36474
rect 2646 36422 2698 36474
rect 2710 36422 2762 36474
rect 2774 36422 2826 36474
rect 2838 36422 2890 36474
rect 5846 36422 5898 36474
rect 5910 36422 5962 36474
rect 5974 36422 6026 36474
rect 6038 36422 6090 36474
rect 6102 36422 6154 36474
rect 9110 36422 9162 36474
rect 9174 36422 9226 36474
rect 9238 36422 9290 36474
rect 9302 36422 9354 36474
rect 9366 36422 9418 36474
rect 6828 36320 6880 36372
rect 9680 36320 9732 36372
rect 756 36184 808 36236
rect 1492 36159 1544 36168
rect 1492 36125 1501 36159
rect 1501 36125 1535 36159
rect 1535 36125 1544 36159
rect 1492 36116 1544 36125
rect 2504 36116 2556 36168
rect 5540 36116 5592 36168
rect 9772 36116 9824 36168
rect 10048 36023 10100 36032
rect 10048 35989 10057 36023
rect 10057 35989 10091 36023
rect 10091 35989 10100 36023
rect 10048 35980 10100 35989
rect 4214 35878 4266 35930
rect 4278 35878 4330 35930
rect 4342 35878 4394 35930
rect 4406 35878 4458 35930
rect 4470 35878 4522 35930
rect 7478 35878 7530 35930
rect 7542 35878 7594 35930
rect 7606 35878 7658 35930
rect 7670 35878 7722 35930
rect 7734 35878 7786 35930
rect 5540 35776 5592 35828
rect 9956 35819 10008 35828
rect 9956 35785 9965 35819
rect 9965 35785 9999 35819
rect 9999 35785 10008 35819
rect 9956 35776 10008 35785
rect 3516 35708 3568 35760
rect 4436 35708 4488 35760
rect 480 35640 532 35692
rect 3792 35640 3844 35692
rect 5724 35708 5776 35760
rect 4896 35640 4948 35692
rect 4620 35615 4672 35624
rect 4620 35581 4629 35615
rect 4629 35581 4663 35615
rect 4663 35581 4672 35615
rect 4620 35572 4672 35581
rect 2320 35547 2372 35556
rect 2320 35513 2329 35547
rect 2329 35513 2363 35547
rect 2363 35513 2372 35547
rect 2320 35504 2372 35513
rect 1584 35479 1636 35488
rect 1584 35445 1593 35479
rect 1593 35445 1627 35479
rect 1627 35445 1636 35479
rect 1584 35436 1636 35445
rect 2582 35334 2634 35386
rect 2646 35334 2698 35386
rect 2710 35334 2762 35386
rect 2774 35334 2826 35386
rect 2838 35334 2890 35386
rect 5846 35334 5898 35386
rect 5910 35334 5962 35386
rect 5974 35334 6026 35386
rect 6038 35334 6090 35386
rect 6102 35334 6154 35386
rect 9110 35334 9162 35386
rect 9174 35334 9226 35386
rect 9238 35334 9290 35386
rect 9302 35334 9354 35386
rect 9366 35334 9418 35386
rect 1492 35232 1544 35284
rect 4896 35275 4948 35284
rect 4896 35241 4905 35275
rect 4905 35241 4939 35275
rect 4939 35241 4948 35275
rect 4896 35232 4948 35241
rect 1492 35028 1544 35080
rect 4620 35164 4672 35216
rect 3976 35096 4028 35148
rect 4436 35096 4488 35148
rect 2412 35071 2464 35080
rect 1400 34960 1452 35012
rect 2412 35037 2421 35071
rect 2421 35037 2455 35071
rect 2455 35037 2464 35071
rect 2412 35028 2464 35037
rect 3700 35028 3752 35080
rect 5172 35164 5224 35216
rect 4988 35028 5040 35080
rect 5172 35028 5224 35080
rect 2504 34960 2556 35012
rect 2780 34892 2832 34944
rect 10048 34935 10100 34944
rect 10048 34901 10057 34935
rect 10057 34901 10091 34935
rect 10091 34901 10100 34935
rect 10048 34892 10100 34901
rect 4214 34790 4266 34842
rect 4278 34790 4330 34842
rect 4342 34790 4394 34842
rect 4406 34790 4458 34842
rect 4470 34790 4522 34842
rect 7478 34790 7530 34842
rect 7542 34790 7594 34842
rect 7606 34790 7658 34842
rect 7670 34790 7722 34842
rect 7734 34790 7786 34842
rect 1584 34731 1636 34740
rect 1584 34697 1593 34731
rect 1593 34697 1627 34731
rect 1627 34697 1636 34731
rect 1584 34688 1636 34697
rect 9588 34688 9640 34740
rect 3976 34620 4028 34672
rect 10232 34620 10284 34672
rect 388 34552 440 34604
rect 2044 34552 2096 34604
rect 2964 34552 3016 34604
rect 4160 34595 4212 34604
rect 4160 34561 4169 34595
rect 4169 34561 4203 34595
rect 4203 34561 4212 34595
rect 4160 34552 4212 34561
rect 9680 34552 9732 34604
rect 3976 34527 4028 34536
rect 3976 34493 3985 34527
rect 3985 34493 4019 34527
rect 4019 34493 4028 34527
rect 3976 34484 4028 34493
rect 2044 34416 2096 34468
rect 2228 34416 2280 34468
rect 1400 34348 1452 34400
rect 3056 34391 3108 34400
rect 3056 34357 3065 34391
rect 3065 34357 3099 34391
rect 3099 34357 3108 34391
rect 3056 34348 3108 34357
rect 2582 34246 2634 34298
rect 2646 34246 2698 34298
rect 2710 34246 2762 34298
rect 2774 34246 2826 34298
rect 2838 34246 2890 34298
rect 5846 34246 5898 34298
rect 5910 34246 5962 34298
rect 5974 34246 6026 34298
rect 6038 34246 6090 34298
rect 6102 34246 6154 34298
rect 9110 34246 9162 34298
rect 9174 34246 9226 34298
rect 9238 34246 9290 34298
rect 9302 34246 9354 34298
rect 9366 34246 9418 34298
rect 9864 34144 9916 34196
rect 204 34076 256 34128
rect 10140 34076 10192 34128
rect 2412 33940 2464 33992
rect 2872 33985 2924 33992
rect 2872 33951 2901 33985
rect 2901 33951 2924 33985
rect 2872 33940 2924 33951
rect 2228 33872 2280 33924
rect 2320 33872 2372 33924
rect 10140 33983 10192 33992
rect 10140 33949 10149 33983
rect 10149 33949 10183 33983
rect 10183 33949 10192 33983
rect 10140 33940 10192 33949
rect 3792 33872 3844 33924
rect 3976 33804 4028 33856
rect 4214 33702 4266 33754
rect 4278 33702 4330 33754
rect 4342 33702 4394 33754
rect 4406 33702 4458 33754
rect 4470 33702 4522 33754
rect 7478 33702 7530 33754
rect 7542 33702 7594 33754
rect 7606 33702 7658 33754
rect 7670 33702 7722 33754
rect 7734 33702 7786 33754
rect 2228 33643 2280 33652
rect 2228 33609 2237 33643
rect 2237 33609 2271 33643
rect 2271 33609 2280 33643
rect 2228 33600 2280 33609
rect 3240 33600 3292 33652
rect 10140 33600 10192 33652
rect 2320 33532 2372 33584
rect 2504 33532 2556 33584
rect 2228 33464 2280 33516
rect 2964 33464 3016 33516
rect 3056 33464 3108 33516
rect 3240 33464 3292 33516
rect 3792 33464 3844 33516
rect 5540 33464 5592 33516
rect 2504 33396 2556 33448
rect 2872 33328 2924 33380
rect 3056 33328 3108 33380
rect 10048 33371 10100 33380
rect 10048 33337 10057 33371
rect 10057 33337 10091 33371
rect 10091 33337 10100 33371
rect 10048 33328 10100 33337
rect 2582 33158 2634 33210
rect 2646 33158 2698 33210
rect 2710 33158 2762 33210
rect 2774 33158 2826 33210
rect 2838 33158 2890 33210
rect 5846 33158 5898 33210
rect 5910 33158 5962 33210
rect 5974 33158 6026 33210
rect 6038 33158 6090 33210
rect 6102 33158 6154 33210
rect 9110 33158 9162 33210
rect 9174 33158 9226 33210
rect 9238 33158 9290 33210
rect 9302 33158 9354 33210
rect 9366 33158 9418 33210
rect 9680 33056 9732 33108
rect 1492 32920 1544 32972
rect 1676 32852 1728 32904
rect 2136 32895 2188 32904
rect 2136 32861 2145 32895
rect 2145 32861 2179 32895
rect 2179 32861 2188 32895
rect 2136 32852 2188 32861
rect 3792 32852 3844 32904
rect 9864 32895 9916 32904
rect 9864 32861 9873 32895
rect 9873 32861 9907 32895
rect 9907 32861 9916 32895
rect 9864 32852 9916 32861
rect 2320 32759 2372 32768
rect 2320 32725 2329 32759
rect 2329 32725 2363 32759
rect 2363 32725 2372 32759
rect 2320 32716 2372 32725
rect 2780 32716 2832 32768
rect 4988 32716 5040 32768
rect 5724 32716 5776 32768
rect 10048 32759 10100 32768
rect 10048 32725 10057 32759
rect 10057 32725 10091 32759
rect 10091 32725 10100 32759
rect 10048 32716 10100 32725
rect 4214 32614 4266 32666
rect 4278 32614 4330 32666
rect 4342 32614 4394 32666
rect 4406 32614 4458 32666
rect 4470 32614 4522 32666
rect 7478 32614 7530 32666
rect 7542 32614 7594 32666
rect 7606 32614 7658 32666
rect 7670 32614 7722 32666
rect 7734 32614 7786 32666
rect 1584 32512 1636 32564
rect 2964 32512 3016 32564
rect 9864 32512 9916 32564
rect 2228 32419 2280 32428
rect 2228 32385 2237 32419
rect 2237 32385 2271 32419
rect 2271 32385 2280 32419
rect 2228 32376 2280 32385
rect 3884 32444 3936 32496
rect 940 32308 992 32360
rect 3700 32308 3752 32360
rect 3056 32283 3108 32292
rect 3056 32249 3065 32283
rect 3065 32249 3099 32283
rect 3099 32249 3108 32283
rect 3056 32240 3108 32249
rect 3424 32172 3476 32224
rect 3700 32172 3752 32224
rect 4988 32376 5040 32428
rect 5172 32240 5224 32292
rect 4712 32172 4764 32224
rect 2582 32070 2634 32122
rect 2646 32070 2698 32122
rect 2710 32070 2762 32122
rect 2774 32070 2826 32122
rect 2838 32070 2890 32122
rect 5846 32070 5898 32122
rect 5910 32070 5962 32122
rect 5974 32070 6026 32122
rect 6038 32070 6090 32122
rect 6102 32070 6154 32122
rect 9110 32070 9162 32122
rect 9174 32070 9226 32122
rect 9238 32070 9290 32122
rect 9302 32070 9354 32122
rect 9366 32070 9418 32122
rect 848 31968 900 32020
rect 2504 31968 2556 32020
rect 1860 31900 1912 31952
rect 2596 31900 2648 31952
rect 4252 31968 4304 32020
rect 9772 31968 9824 32020
rect 3976 31943 4028 31952
rect 3976 31909 3985 31943
rect 3985 31909 4019 31943
rect 4019 31909 4028 31943
rect 3976 31900 4028 31909
rect 10048 31943 10100 31952
rect 10048 31909 10057 31943
rect 10057 31909 10091 31943
rect 10091 31909 10100 31943
rect 10048 31900 10100 31909
rect 664 31832 716 31884
rect 2228 31832 2280 31884
rect 2504 31832 2556 31884
rect 4620 31832 4672 31884
rect 1124 31764 1176 31816
rect 1400 31764 1452 31816
rect 2136 31764 2188 31816
rect 5356 31832 5408 31884
rect 5632 31832 5684 31884
rect 1584 31696 1636 31748
rect 1860 31739 1912 31748
rect 1860 31705 1869 31739
rect 1869 31705 1903 31739
rect 1903 31705 1912 31739
rect 1860 31696 1912 31705
rect 2228 31696 2280 31748
rect 3056 31696 3108 31748
rect 1124 31628 1176 31680
rect 2320 31628 2372 31680
rect 2688 31628 2740 31680
rect 4214 31526 4266 31578
rect 4278 31526 4330 31578
rect 4342 31526 4394 31578
rect 4406 31526 4458 31578
rect 4470 31526 4522 31578
rect 7478 31526 7530 31578
rect 7542 31526 7594 31578
rect 7606 31526 7658 31578
rect 7670 31526 7722 31578
rect 7734 31526 7786 31578
rect 1860 31424 1912 31476
rect 2320 31424 2372 31476
rect 2504 31424 2556 31476
rect 3056 31424 3108 31476
rect 2688 31356 2740 31408
rect 664 31288 716 31340
rect 2964 31288 3016 31340
rect 5356 31288 5408 31340
rect 5632 31288 5684 31340
rect 9864 31331 9916 31340
rect 9864 31297 9873 31331
rect 9873 31297 9907 31331
rect 9907 31297 9916 31331
rect 9864 31288 9916 31297
rect 848 31220 900 31272
rect 3884 31220 3936 31272
rect 2412 31152 2464 31204
rect 2596 31152 2648 31204
rect 4896 31152 4948 31204
rect 10048 31127 10100 31136
rect 10048 31093 10057 31127
rect 10057 31093 10091 31127
rect 10091 31093 10100 31127
rect 10048 31084 10100 31093
rect 2582 30982 2634 31034
rect 2646 30982 2698 31034
rect 2710 30982 2762 31034
rect 2774 30982 2826 31034
rect 2838 30982 2890 31034
rect 5846 30982 5898 31034
rect 5910 30982 5962 31034
rect 5974 30982 6026 31034
rect 6038 30982 6090 31034
rect 6102 30982 6154 31034
rect 9110 30982 9162 31034
rect 9174 30982 9226 31034
rect 9238 30982 9290 31034
rect 9302 30982 9354 31034
rect 9366 30982 9418 31034
rect 3332 30880 3384 30932
rect 4712 30812 4764 30864
rect 4896 30812 4948 30864
rect 1768 30676 1820 30728
rect 4528 30676 4580 30728
rect 4712 30676 4764 30728
rect 8300 30676 8352 30728
rect 1860 30651 1912 30660
rect 1860 30617 1869 30651
rect 1869 30617 1903 30651
rect 1903 30617 1912 30651
rect 1860 30608 1912 30617
rect 2780 30540 2832 30592
rect 10048 30583 10100 30592
rect 10048 30549 10057 30583
rect 10057 30549 10091 30583
rect 10091 30549 10100 30583
rect 10048 30540 10100 30549
rect 4214 30438 4266 30490
rect 4278 30438 4330 30490
rect 4342 30438 4394 30490
rect 4406 30438 4458 30490
rect 4470 30438 4522 30490
rect 7478 30438 7530 30490
rect 7542 30438 7594 30490
rect 7606 30438 7658 30490
rect 7670 30438 7722 30490
rect 7734 30438 7786 30490
rect 3792 30336 3844 30388
rect 1124 30268 1176 30320
rect 2044 30268 2096 30320
rect 1676 30243 1728 30252
rect 1676 30209 1685 30243
rect 1685 30209 1719 30243
rect 1719 30209 1728 30243
rect 1676 30200 1728 30209
rect 4528 30268 4580 30320
rect 5724 30268 5776 30320
rect 2320 30175 2372 30184
rect 2320 30141 2329 30175
rect 2329 30141 2363 30175
rect 2363 30141 2372 30175
rect 2320 30132 2372 30141
rect 3792 30200 3844 30252
rect 5632 30200 5684 30252
rect 2964 30132 3016 30184
rect 3332 30107 3384 30116
rect 3332 30073 3341 30107
rect 3341 30073 3375 30107
rect 3375 30073 3384 30107
rect 3332 30064 3384 30073
rect 4620 30064 4672 30116
rect 848 29996 900 30048
rect 1860 29996 1912 30048
rect 9864 29996 9916 30048
rect 2582 29894 2634 29946
rect 2646 29894 2698 29946
rect 2710 29894 2762 29946
rect 2774 29894 2826 29946
rect 2838 29894 2890 29946
rect 5846 29894 5898 29946
rect 5910 29894 5962 29946
rect 5974 29894 6026 29946
rect 6038 29894 6090 29946
rect 6102 29894 6154 29946
rect 9110 29894 9162 29946
rect 9174 29894 9226 29946
rect 9238 29894 9290 29946
rect 9302 29894 9354 29946
rect 9366 29894 9418 29946
rect 756 29792 808 29844
rect 8300 29792 8352 29844
rect 6920 29588 6972 29640
rect 7840 29631 7892 29640
rect 7840 29597 7849 29631
rect 7849 29597 7883 29631
rect 7883 29597 7892 29631
rect 7840 29588 7892 29597
rect 10140 29631 10192 29640
rect 10140 29597 10149 29631
rect 10149 29597 10183 29631
rect 10183 29597 10192 29631
rect 10140 29588 10192 29597
rect 2780 29520 2832 29572
rect 3056 29452 3108 29504
rect 4214 29350 4266 29402
rect 4278 29350 4330 29402
rect 4342 29350 4394 29402
rect 4406 29350 4458 29402
rect 4470 29350 4522 29402
rect 7478 29350 7530 29402
rect 7542 29350 7594 29402
rect 7606 29350 7658 29402
rect 7670 29350 7722 29402
rect 7734 29350 7786 29402
rect 112 29248 164 29300
rect 3148 29248 3200 29300
rect 2964 29112 3016 29164
rect 3148 29112 3200 29164
rect 10140 29019 10192 29028
rect 10140 28985 10149 29019
rect 10149 28985 10183 29019
rect 10183 28985 10192 29019
rect 10140 28976 10192 28985
rect 2582 28806 2634 28858
rect 2646 28806 2698 28858
rect 2710 28806 2762 28858
rect 2774 28806 2826 28858
rect 2838 28806 2890 28858
rect 5846 28806 5898 28858
rect 5910 28806 5962 28858
rect 5974 28806 6026 28858
rect 6038 28806 6090 28858
rect 6102 28806 6154 28858
rect 9110 28806 9162 28858
rect 9174 28806 9226 28858
rect 9238 28806 9290 28858
rect 9302 28806 9354 28858
rect 9366 28806 9418 28858
rect 6460 28704 6512 28756
rect 2872 28636 2924 28688
rect 3056 28636 3108 28688
rect 4068 28679 4120 28688
rect 4068 28645 4077 28679
rect 4077 28645 4111 28679
rect 4111 28645 4120 28679
rect 4068 28636 4120 28645
rect 6368 28568 6420 28620
rect 3056 28500 3108 28552
rect 3332 28432 3384 28484
rect 2964 28364 3016 28416
rect 4214 28262 4266 28314
rect 4278 28262 4330 28314
rect 4342 28262 4394 28314
rect 4406 28262 4458 28314
rect 4470 28262 4522 28314
rect 7478 28262 7530 28314
rect 7542 28262 7594 28314
rect 7606 28262 7658 28314
rect 7670 28262 7722 28314
rect 7734 28262 7786 28314
rect 1400 28160 1452 28212
rect 1676 28160 1728 28212
rect 3148 28160 3200 28212
rect 3332 28160 3384 28212
rect 3608 28160 3660 28212
rect 4988 28160 5040 28212
rect 5356 28160 5408 28212
rect 664 28092 716 28144
rect 1952 28024 2004 28076
rect 1400 27999 1452 28008
rect 1400 27965 1409 27999
rect 1409 27965 1443 27999
rect 1443 27965 1452 27999
rect 1400 27956 1452 27965
rect 1952 27888 2004 27940
rect 5448 28092 5500 28144
rect 3608 28067 3660 28076
rect 3608 28033 3617 28067
rect 3617 28033 3651 28067
rect 3651 28033 3660 28067
rect 3608 28024 3660 28033
rect 3884 28024 3936 28076
rect 5172 28024 5224 28076
rect 5356 28024 5408 28076
rect 2504 27956 2556 28008
rect 7196 27956 7248 28008
rect 9956 27999 10008 28008
rect 9956 27965 9965 27999
rect 9965 27965 9999 27999
rect 9999 27965 10008 27999
rect 9956 27956 10008 27965
rect 2872 27888 2924 27940
rect 3148 27888 3200 27940
rect 4436 27888 4488 27940
rect 5632 27888 5684 27940
rect 2582 27718 2634 27770
rect 2646 27718 2698 27770
rect 2710 27718 2762 27770
rect 2774 27718 2826 27770
rect 2838 27718 2890 27770
rect 5846 27718 5898 27770
rect 5910 27718 5962 27770
rect 5974 27718 6026 27770
rect 6038 27718 6090 27770
rect 6102 27718 6154 27770
rect 9110 27718 9162 27770
rect 9174 27718 9226 27770
rect 9238 27718 9290 27770
rect 9302 27718 9354 27770
rect 9366 27718 9418 27770
rect 3056 27591 3108 27600
rect 3056 27557 3065 27591
rect 3065 27557 3099 27591
rect 3099 27557 3108 27591
rect 3056 27548 3108 27557
rect 4620 27548 4672 27600
rect 1216 27480 1268 27532
rect 4068 27480 4120 27532
rect 1032 27412 1084 27464
rect 1952 27412 2004 27464
rect 4620 27344 4672 27396
rect 9956 27319 10008 27328
rect 9956 27285 9965 27319
rect 9965 27285 9999 27319
rect 9999 27285 10008 27319
rect 9956 27276 10008 27285
rect 4214 27174 4266 27226
rect 4278 27174 4330 27226
rect 4342 27174 4394 27226
rect 4406 27174 4458 27226
rect 4470 27174 4522 27226
rect 7478 27174 7530 27226
rect 7542 27174 7594 27226
rect 7606 27174 7658 27226
rect 7670 27174 7722 27226
rect 7734 27174 7786 27226
rect 2964 27072 3016 27124
rect 3700 27115 3752 27124
rect 3700 27081 3709 27115
rect 3709 27081 3743 27115
rect 3743 27081 3752 27115
rect 3700 27072 3752 27081
rect 1952 26936 2004 26988
rect 3056 26936 3108 26988
rect 3608 26979 3660 26988
rect 3608 26945 3617 26979
rect 3617 26945 3651 26979
rect 3651 26945 3660 26979
rect 3608 26936 3660 26945
rect 2320 26868 2372 26920
rect 2412 26868 2464 26920
rect 4804 26868 4856 26920
rect 4988 26868 5040 26920
rect 1952 26800 2004 26852
rect 2136 26800 2188 26852
rect 1860 26732 1912 26784
rect 5080 26732 5132 26784
rect 5448 26732 5500 26784
rect 10140 26775 10192 26784
rect 10140 26741 10149 26775
rect 10149 26741 10183 26775
rect 10183 26741 10192 26775
rect 10140 26732 10192 26741
rect 2582 26630 2634 26682
rect 2646 26630 2698 26682
rect 2710 26630 2762 26682
rect 2774 26630 2826 26682
rect 2838 26630 2890 26682
rect 5846 26630 5898 26682
rect 5910 26630 5962 26682
rect 5974 26630 6026 26682
rect 6038 26630 6090 26682
rect 6102 26630 6154 26682
rect 9110 26630 9162 26682
rect 9174 26630 9226 26682
rect 9238 26630 9290 26682
rect 9302 26630 9354 26682
rect 9366 26630 9418 26682
rect 3332 26460 3384 26512
rect 5080 26528 5132 26580
rect 5540 26528 5592 26580
rect 4712 26460 4764 26512
rect 4896 26460 4948 26512
rect 5632 26460 5684 26512
rect 6276 26392 6328 26444
rect 1860 26367 1912 26376
rect 1860 26333 1869 26367
rect 1869 26333 1903 26367
rect 1903 26333 1912 26367
rect 1860 26324 1912 26333
rect 2320 26256 2372 26308
rect 2596 26299 2648 26308
rect 2596 26265 2605 26299
rect 2605 26265 2639 26299
rect 2639 26265 2648 26299
rect 2596 26256 2648 26265
rect 3332 26256 3384 26308
rect 3792 26256 3844 26308
rect 1860 26188 1912 26240
rect 3516 26188 3568 26240
rect 4214 26086 4266 26138
rect 4278 26086 4330 26138
rect 4342 26086 4394 26138
rect 4406 26086 4458 26138
rect 4470 26086 4522 26138
rect 7478 26086 7530 26138
rect 7542 26086 7594 26138
rect 7606 26086 7658 26138
rect 7670 26086 7722 26138
rect 7734 26086 7786 26138
rect 2320 25984 2372 26036
rect 2504 25984 2556 26036
rect 3884 25984 3936 26036
rect 1768 25848 1820 25900
rect 2964 25848 3016 25900
rect 1400 25823 1452 25832
rect 1400 25789 1409 25823
rect 1409 25789 1443 25823
rect 1443 25789 1452 25823
rect 1400 25780 1452 25789
rect 3516 25780 3568 25832
rect 296 25712 348 25764
rect 1768 25712 1820 25764
rect 10140 25687 10192 25696
rect 10140 25653 10149 25687
rect 10149 25653 10183 25687
rect 10183 25653 10192 25687
rect 10140 25644 10192 25653
rect 2582 25542 2634 25594
rect 2646 25542 2698 25594
rect 2710 25542 2762 25594
rect 2774 25542 2826 25594
rect 2838 25542 2890 25594
rect 5846 25542 5898 25594
rect 5910 25542 5962 25594
rect 5974 25542 6026 25594
rect 6038 25542 6090 25594
rect 6102 25542 6154 25594
rect 9110 25542 9162 25594
rect 9174 25542 9226 25594
rect 9238 25542 9290 25594
rect 9302 25542 9354 25594
rect 9366 25542 9418 25594
rect 3332 25440 3384 25492
rect 4528 25304 4580 25356
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 2964 25279 3016 25288
rect 2504 25168 2556 25220
rect 2964 25245 2973 25279
rect 2973 25245 3007 25279
rect 3007 25245 3016 25279
rect 2964 25236 3016 25245
rect 3700 25236 3752 25288
rect 10140 25279 10192 25288
rect 10140 25245 10149 25279
rect 10149 25245 10183 25279
rect 10183 25245 10192 25279
rect 10140 25236 10192 25245
rect 4214 24998 4266 25050
rect 4278 24998 4330 25050
rect 4342 24998 4394 25050
rect 4406 24998 4458 25050
rect 4470 24998 4522 25050
rect 7478 24998 7530 25050
rect 7542 24998 7594 25050
rect 7606 24998 7658 25050
rect 7670 24998 7722 25050
rect 7734 24998 7786 25050
rect 2780 24803 2832 24812
rect 2780 24769 2789 24803
rect 2789 24769 2823 24803
rect 2823 24769 2832 24803
rect 3332 24803 3384 24812
rect 2780 24760 2832 24769
rect 3332 24769 3341 24803
rect 3341 24769 3375 24803
rect 3375 24769 3384 24803
rect 3332 24760 3384 24769
rect 3424 24760 3476 24812
rect 4160 24760 4212 24812
rect 4896 24760 4948 24812
rect 2964 24692 3016 24744
rect 3148 24692 3200 24744
rect 1124 24556 1176 24608
rect 4620 24624 4672 24676
rect 4896 24624 4948 24676
rect 3148 24556 3200 24608
rect 3332 24556 3384 24608
rect 2582 24454 2634 24506
rect 2646 24454 2698 24506
rect 2710 24454 2762 24506
rect 2774 24454 2826 24506
rect 2838 24454 2890 24506
rect 5846 24454 5898 24506
rect 5910 24454 5962 24506
rect 5974 24454 6026 24506
rect 6038 24454 6090 24506
rect 6102 24454 6154 24506
rect 9110 24454 9162 24506
rect 9174 24454 9226 24506
rect 9238 24454 9290 24506
rect 9302 24454 9354 24506
rect 9366 24454 9418 24506
rect 2872 24284 2924 24336
rect 3056 24284 3108 24336
rect 2044 24216 2096 24268
rect 4160 24216 4212 24268
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 10140 24191 10192 24200
rect 10140 24157 10149 24191
rect 10149 24157 10183 24191
rect 10183 24157 10192 24191
rect 10140 24148 10192 24157
rect 3056 24080 3108 24132
rect 1768 24012 1820 24064
rect 2136 24012 2188 24064
rect 4214 23910 4266 23962
rect 4278 23910 4330 23962
rect 4342 23910 4394 23962
rect 4406 23910 4458 23962
rect 4470 23910 4522 23962
rect 7478 23910 7530 23962
rect 7542 23910 7594 23962
rect 7606 23910 7658 23962
rect 7670 23910 7722 23962
rect 7734 23910 7786 23962
rect 1676 23715 1728 23724
rect 1676 23681 1685 23715
rect 1685 23681 1719 23715
rect 1719 23681 1728 23715
rect 1676 23672 1728 23681
rect 3976 23672 4028 23724
rect 1216 23604 1268 23656
rect 2780 23604 2832 23656
rect 10140 23511 10192 23520
rect 10140 23477 10149 23511
rect 10149 23477 10183 23511
rect 10183 23477 10192 23511
rect 10140 23468 10192 23477
rect 2582 23366 2634 23418
rect 2646 23366 2698 23418
rect 2710 23366 2762 23418
rect 2774 23366 2826 23418
rect 2838 23366 2890 23418
rect 5846 23366 5898 23418
rect 5910 23366 5962 23418
rect 5974 23366 6026 23418
rect 6038 23366 6090 23418
rect 6102 23366 6154 23418
rect 9110 23366 9162 23418
rect 9174 23366 9226 23418
rect 9238 23366 9290 23418
rect 9302 23366 9354 23418
rect 9366 23366 9418 23418
rect 3056 23307 3108 23316
rect 3056 23273 3065 23307
rect 3065 23273 3099 23307
rect 3099 23273 3108 23307
rect 3056 23264 3108 23273
rect 3608 23128 3660 23180
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2504 23060 2556 23112
rect 2964 23060 3016 23112
rect 4214 22822 4266 22874
rect 4278 22822 4330 22874
rect 4342 22822 4394 22874
rect 4406 22822 4458 22874
rect 4470 22822 4522 22874
rect 7478 22822 7530 22874
rect 7542 22822 7594 22874
rect 7606 22822 7658 22874
rect 7670 22822 7722 22874
rect 7734 22822 7786 22874
rect 3056 22763 3108 22772
rect 3056 22729 3065 22763
rect 3065 22729 3099 22763
rect 3099 22729 3108 22763
rect 3056 22720 3108 22729
rect 3700 22652 3752 22704
rect 3976 22652 4028 22704
rect 5080 22652 5132 22704
rect 1216 22516 1268 22568
rect 3608 22627 3660 22636
rect 3608 22593 3617 22627
rect 3617 22593 3651 22627
rect 3651 22593 3660 22627
rect 3608 22584 3660 22593
rect 4160 22584 4212 22636
rect 3424 22516 3476 22568
rect 1676 22448 1728 22500
rect 10140 22491 10192 22500
rect 10140 22457 10149 22491
rect 10149 22457 10183 22491
rect 10183 22457 10192 22491
rect 10140 22448 10192 22457
rect 3700 22423 3752 22432
rect 3700 22389 3709 22423
rect 3709 22389 3743 22423
rect 3743 22389 3752 22423
rect 3700 22380 3752 22389
rect 940 22244 992 22296
rect 2582 22278 2634 22330
rect 2646 22278 2698 22330
rect 2710 22278 2762 22330
rect 2774 22278 2826 22330
rect 2838 22278 2890 22330
rect 5846 22278 5898 22330
rect 5910 22278 5962 22330
rect 5974 22278 6026 22330
rect 6038 22278 6090 22330
rect 6102 22278 6154 22330
rect 9110 22278 9162 22330
rect 9174 22278 9226 22330
rect 9238 22278 9290 22330
rect 9302 22278 9354 22330
rect 9366 22278 9418 22330
rect 2504 22176 2556 22228
rect 940 22108 992 22160
rect 1768 22108 1820 22160
rect 2320 22108 2372 22160
rect 2688 22108 2740 22160
rect 10140 22151 10192 22160
rect 10140 22117 10149 22151
rect 10149 22117 10183 22151
rect 10183 22117 10192 22151
rect 10140 22108 10192 22117
rect 1492 22040 1544 22092
rect 2228 22040 2280 22092
rect 2596 22040 2648 22092
rect 3148 22040 3200 22092
rect 4620 22040 4672 22092
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 2044 21972 2096 22024
rect 2964 21972 3016 22024
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 4214 21734 4266 21786
rect 4278 21734 4330 21786
rect 4342 21734 4394 21786
rect 4406 21734 4458 21786
rect 4470 21734 4522 21786
rect 7478 21734 7530 21786
rect 7542 21734 7594 21786
rect 7606 21734 7658 21786
rect 7670 21734 7722 21786
rect 7734 21734 7786 21786
rect 4068 21632 4120 21684
rect 940 21564 992 21616
rect 4804 21564 4856 21616
rect 2320 21496 2372 21548
rect 2964 21496 3016 21548
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 1768 21428 1820 21480
rect 2688 21428 2740 21480
rect 3424 21428 3476 21480
rect 2320 21360 2372 21412
rect 2596 21360 2648 21412
rect 2964 21403 3016 21412
rect 2964 21369 2973 21403
rect 2973 21369 3007 21403
rect 3007 21369 3016 21403
rect 2964 21360 3016 21369
rect 10140 21335 10192 21344
rect 10140 21301 10149 21335
rect 10149 21301 10183 21335
rect 10183 21301 10192 21335
rect 10140 21292 10192 21301
rect 2582 21190 2634 21242
rect 2646 21190 2698 21242
rect 2710 21190 2762 21242
rect 2774 21190 2826 21242
rect 2838 21190 2890 21242
rect 5846 21190 5898 21242
rect 5910 21190 5962 21242
rect 5974 21190 6026 21242
rect 6038 21190 6090 21242
rect 6102 21190 6154 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 9238 21190 9290 21242
rect 9302 21190 9354 21242
rect 9366 21190 9418 21242
rect 3608 21088 3660 21140
rect 2412 20952 2464 21004
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 1584 20884 1636 20936
rect 2964 20884 3016 20936
rect 4214 20646 4266 20698
rect 4278 20646 4330 20698
rect 4342 20646 4394 20698
rect 4406 20646 4458 20698
rect 4470 20646 4522 20698
rect 7478 20646 7530 20698
rect 7542 20646 7594 20698
rect 7606 20646 7658 20698
rect 7670 20646 7722 20698
rect 7734 20646 7786 20698
rect 7840 20544 7892 20596
rect 2228 20408 2280 20460
rect 3608 20408 3660 20460
rect 3976 20408 4028 20460
rect 9772 20408 9824 20460
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 1768 20340 1820 20392
rect 10048 20315 10100 20324
rect 10048 20281 10057 20315
rect 10057 20281 10091 20315
rect 10091 20281 10100 20315
rect 10048 20272 10100 20281
rect 2582 20102 2634 20154
rect 2646 20102 2698 20154
rect 2710 20102 2762 20154
rect 2774 20102 2826 20154
rect 2838 20102 2890 20154
rect 5846 20102 5898 20154
rect 5910 20102 5962 20154
rect 5974 20102 6026 20154
rect 6038 20102 6090 20154
rect 6102 20102 6154 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 9238 20102 9290 20154
rect 9302 20102 9354 20154
rect 9366 20102 9418 20154
rect 2504 20000 2556 20052
rect 3884 20000 3936 20052
rect 1860 19932 1912 19984
rect 2412 19932 2464 19984
rect 1768 19839 1820 19848
rect 1768 19805 1777 19839
rect 1777 19805 1811 19839
rect 1811 19805 1820 19839
rect 1768 19796 1820 19805
rect 2964 19864 3016 19916
rect 2872 19796 2924 19848
rect 3976 19839 4028 19848
rect 3976 19805 3985 19839
rect 3985 19805 4019 19839
rect 4019 19805 4028 19839
rect 3976 19796 4028 19805
rect 9864 19839 9916 19848
rect 9864 19805 9873 19839
rect 9873 19805 9907 19839
rect 9907 19805 9916 19839
rect 9864 19796 9916 19805
rect 1860 19660 1912 19712
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 4214 19558 4266 19610
rect 4278 19558 4330 19610
rect 4342 19558 4394 19610
rect 4406 19558 4458 19610
rect 4470 19558 4522 19610
rect 7478 19558 7530 19610
rect 7542 19558 7594 19610
rect 7606 19558 7658 19610
rect 7670 19558 7722 19610
rect 7734 19558 7786 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 2412 19456 2464 19508
rect 9864 19499 9916 19508
rect 9864 19465 9873 19499
rect 9873 19465 9907 19499
rect 9907 19465 9916 19499
rect 9864 19456 9916 19465
rect 1860 19431 1912 19440
rect 1860 19397 1869 19431
rect 1869 19397 1903 19431
rect 1903 19397 1912 19431
rect 1860 19388 1912 19397
rect 2412 19320 2464 19372
rect 2780 19320 2832 19372
rect 3148 19320 3200 19372
rect 5448 19320 5500 19372
rect 1400 19116 1452 19168
rect 1676 19116 1728 19168
rect 2582 19014 2634 19066
rect 2646 19014 2698 19066
rect 2710 19014 2762 19066
rect 2774 19014 2826 19066
rect 2838 19014 2890 19066
rect 5846 19014 5898 19066
rect 5910 19014 5962 19066
rect 5974 19014 6026 19066
rect 6038 19014 6090 19066
rect 6102 19014 6154 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 9238 19014 9290 19066
rect 9302 19014 9354 19066
rect 9366 19014 9418 19066
rect 1584 18912 1636 18964
rect 2044 18955 2096 18964
rect 2044 18921 2053 18955
rect 2053 18921 2087 18955
rect 2087 18921 2096 18955
rect 2044 18912 2096 18921
rect 3424 18912 3476 18964
rect 1492 18708 1544 18760
rect 2228 18751 2280 18760
rect 2228 18717 2237 18751
rect 2237 18717 2271 18751
rect 2271 18717 2280 18751
rect 2228 18708 2280 18717
rect 2872 18751 2924 18760
rect 2872 18717 2881 18751
rect 2881 18717 2915 18751
rect 2915 18717 2924 18751
rect 2872 18708 2924 18717
rect 9220 18708 9272 18760
rect 10048 18615 10100 18624
rect 10048 18581 10057 18615
rect 10057 18581 10091 18615
rect 10091 18581 10100 18615
rect 10048 18572 10100 18581
rect 4214 18470 4266 18522
rect 4278 18470 4330 18522
rect 4342 18470 4394 18522
rect 4406 18470 4458 18522
rect 4470 18470 4522 18522
rect 7478 18470 7530 18522
rect 7542 18470 7594 18522
rect 7606 18470 7658 18522
rect 7670 18470 7722 18522
rect 7734 18470 7786 18522
rect 1400 18411 1452 18420
rect 1400 18377 1409 18411
rect 1409 18377 1443 18411
rect 1443 18377 1452 18411
rect 1400 18368 1452 18377
rect 9220 18411 9272 18420
rect 9220 18377 9229 18411
rect 9229 18377 9263 18411
rect 9263 18377 9272 18411
rect 9220 18368 9272 18377
rect 1032 18300 1084 18352
rect 2412 18300 2464 18352
rect 5448 18300 5500 18352
rect 1400 18232 1452 18284
rect 9864 18275 9916 18284
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 1860 18028 1912 18080
rect 2964 18028 3016 18080
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 2582 17926 2634 17978
rect 2646 17926 2698 17978
rect 2710 17926 2762 17978
rect 2774 17926 2826 17978
rect 2838 17926 2890 17978
rect 5846 17926 5898 17978
rect 5910 17926 5962 17978
rect 5974 17926 6026 17978
rect 6038 17926 6090 17978
rect 6102 17926 6154 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 9238 17926 9290 17978
rect 9302 17926 9354 17978
rect 9366 17926 9418 17978
rect 1768 17824 1820 17876
rect 3792 17756 3844 17808
rect 4804 17688 4856 17740
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 2228 17663 2280 17672
rect 2228 17629 2237 17663
rect 2237 17629 2271 17663
rect 2271 17629 2280 17663
rect 2228 17620 2280 17629
rect 2780 17663 2832 17672
rect 2780 17629 2789 17663
rect 2789 17629 2823 17663
rect 2823 17629 2832 17663
rect 2780 17620 2832 17629
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 9496 17620 9548 17672
rect 3056 17552 3108 17604
rect 10048 17527 10100 17536
rect 10048 17493 10057 17527
rect 10057 17493 10091 17527
rect 10091 17493 10100 17527
rect 10048 17484 10100 17493
rect 4214 17382 4266 17434
rect 4278 17382 4330 17434
rect 4342 17382 4394 17434
rect 4406 17382 4458 17434
rect 4470 17382 4522 17434
rect 7478 17382 7530 17434
rect 7542 17382 7594 17434
rect 7606 17382 7658 17434
rect 7670 17382 7722 17434
rect 7734 17382 7786 17434
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 9864 17280 9916 17332
rect 2964 17212 3016 17264
rect 1492 17144 1544 17196
rect 4620 17144 4672 17196
rect 5448 17144 5500 17196
rect 2228 17008 2280 17060
rect 2780 17008 2832 17060
rect 1400 16983 1452 16992
rect 1400 16949 1409 16983
rect 1409 16949 1443 16983
rect 1443 16949 1452 16983
rect 1400 16940 1452 16949
rect 2582 16838 2634 16890
rect 2646 16838 2698 16890
rect 2710 16838 2762 16890
rect 2774 16838 2826 16890
rect 2838 16838 2890 16890
rect 5846 16838 5898 16890
rect 5910 16838 5962 16890
rect 5974 16838 6026 16890
rect 6038 16838 6090 16890
rect 6102 16838 6154 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 9238 16838 9290 16890
rect 9302 16838 9354 16890
rect 9366 16838 9418 16890
rect 5356 16736 5408 16788
rect 1584 16668 1636 16720
rect 1860 16668 1912 16720
rect 2872 16600 2924 16652
rect 5172 16600 5224 16652
rect 2780 16532 2832 16584
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 9956 16532 10008 16584
rect 2044 16464 2096 16516
rect 2504 16439 2556 16448
rect 2504 16405 2513 16439
rect 2513 16405 2547 16439
rect 2547 16405 2556 16439
rect 2504 16396 2556 16405
rect 3792 16439 3844 16448
rect 3792 16405 3801 16439
rect 3801 16405 3835 16439
rect 3835 16405 3844 16439
rect 3792 16396 3844 16405
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 4214 16294 4266 16346
rect 4278 16294 4330 16346
rect 4342 16294 4394 16346
rect 4406 16294 4458 16346
rect 4470 16294 4522 16346
rect 7478 16294 7530 16346
rect 7542 16294 7594 16346
rect 7606 16294 7658 16346
rect 7670 16294 7722 16346
rect 7734 16294 7786 16346
rect 2872 16192 2924 16244
rect 9496 16192 9548 16244
rect 1400 16056 1452 16108
rect 3792 16124 3844 16176
rect 4068 16056 4120 16108
rect 6184 16056 6236 16108
rect 9680 16056 9732 16108
rect 3792 15988 3844 16040
rect 2504 15920 2556 15972
rect 1952 15852 2004 15904
rect 10048 15895 10100 15904
rect 10048 15861 10057 15895
rect 10057 15861 10091 15895
rect 10091 15861 10100 15895
rect 10048 15852 10100 15861
rect 2582 15750 2634 15802
rect 2646 15750 2698 15802
rect 2710 15750 2762 15802
rect 2774 15750 2826 15802
rect 2838 15750 2890 15802
rect 5846 15750 5898 15802
rect 5910 15750 5962 15802
rect 5974 15750 6026 15802
rect 6038 15750 6090 15802
rect 6102 15750 6154 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 9238 15750 9290 15802
rect 9302 15750 9354 15802
rect 9366 15750 9418 15802
rect 1860 15691 1912 15700
rect 1860 15657 1869 15691
rect 1869 15657 1903 15691
rect 1903 15657 1912 15691
rect 1860 15648 1912 15657
rect 2228 15691 2280 15700
rect 2228 15657 2237 15691
rect 2237 15657 2271 15691
rect 2271 15657 2280 15691
rect 2228 15648 2280 15657
rect 3792 15691 3844 15700
rect 3792 15657 3801 15691
rect 3801 15657 3835 15691
rect 3835 15657 3844 15691
rect 3792 15648 3844 15657
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 1952 15555 2004 15564
rect 1952 15521 1961 15555
rect 1961 15521 1995 15555
rect 1995 15521 2004 15555
rect 1952 15512 2004 15521
rect 2228 15512 2280 15564
rect 6184 15512 6236 15564
rect 1768 15444 1820 15496
rect 2872 15487 2924 15496
rect 2872 15453 2881 15487
rect 2881 15453 2915 15487
rect 2915 15453 2924 15487
rect 2872 15444 2924 15453
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 4896 15444 4948 15496
rect 2320 15308 2372 15360
rect 4214 15206 4266 15258
rect 4278 15206 4330 15258
rect 4342 15206 4394 15258
rect 4406 15206 4458 15258
rect 4470 15206 4522 15258
rect 7478 15206 7530 15258
rect 7542 15206 7594 15258
rect 7606 15206 7658 15258
rect 7670 15206 7722 15258
rect 7734 15206 7786 15258
rect 2136 15147 2188 15156
rect 2136 15113 2145 15147
rect 2145 15113 2179 15147
rect 2179 15113 2188 15147
rect 2136 15104 2188 15113
rect 3148 15036 3200 15088
rect 2412 14968 2464 15020
rect 3424 14968 3476 15020
rect 9956 14968 10008 15020
rect 10048 14875 10100 14884
rect 10048 14841 10057 14875
rect 10057 14841 10091 14875
rect 10091 14841 10100 14875
rect 10048 14832 10100 14841
rect 2228 14764 2280 14816
rect 4804 14764 4856 14816
rect 2582 14662 2634 14714
rect 2646 14662 2698 14714
rect 2710 14662 2762 14714
rect 2774 14662 2826 14714
rect 2838 14662 2890 14714
rect 5846 14662 5898 14714
rect 5910 14662 5962 14714
rect 5974 14662 6026 14714
rect 6038 14662 6090 14714
rect 6102 14662 6154 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 9238 14662 9290 14714
rect 9302 14662 9354 14714
rect 9366 14662 9418 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 1952 14560 2004 14612
rect 2964 14603 3016 14612
rect 2320 14424 2372 14476
rect 2964 14569 2973 14603
rect 2973 14569 3007 14603
rect 3007 14569 3016 14603
rect 2964 14560 3016 14569
rect 2872 14492 2924 14544
rect 4896 14424 4948 14476
rect 3792 14356 3844 14408
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 2136 14288 2188 14340
rect 3056 14288 3108 14340
rect 2688 14220 2740 14272
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 4214 14118 4266 14170
rect 4278 14118 4330 14170
rect 4342 14118 4394 14170
rect 4406 14118 4458 14170
rect 4470 14118 4522 14170
rect 7478 14118 7530 14170
rect 7542 14118 7594 14170
rect 7606 14118 7658 14170
rect 7670 14118 7722 14170
rect 7734 14118 7786 14170
rect 1492 14016 1544 14068
rect 1676 14016 1728 14068
rect 2412 14059 2464 14068
rect 2412 14025 2421 14059
rect 2421 14025 2455 14059
rect 2455 14025 2464 14059
rect 2412 14016 2464 14025
rect 9588 14016 9640 14068
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 3240 13923 3292 13932
rect 3240 13889 3249 13923
rect 3249 13889 3283 13923
rect 3283 13889 3292 13923
rect 3240 13880 3292 13889
rect 3516 13880 3568 13932
rect 3884 13923 3936 13932
rect 3884 13889 3893 13923
rect 3893 13889 3927 13923
rect 3927 13889 3936 13923
rect 3884 13880 3936 13889
rect 1584 13744 1636 13796
rect 3608 13744 3660 13796
rect 2582 13574 2634 13626
rect 2646 13574 2698 13626
rect 2710 13574 2762 13626
rect 2774 13574 2826 13626
rect 2838 13574 2890 13626
rect 5846 13574 5898 13626
rect 5910 13574 5962 13626
rect 5974 13574 6026 13626
rect 6038 13574 6090 13626
rect 6102 13574 6154 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 9238 13574 9290 13626
rect 9302 13574 9354 13626
rect 9366 13574 9418 13626
rect 2412 13472 2464 13524
rect 3792 13447 3844 13456
rect 3792 13413 3801 13447
rect 3801 13413 3835 13447
rect 3835 13413 3844 13447
rect 3792 13404 3844 13413
rect 2320 13336 2372 13388
rect 2872 13336 2924 13388
rect 1308 13268 1360 13320
rect 2504 13268 2556 13320
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 9864 13472 9916 13524
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 1400 13175 1452 13184
rect 1400 13141 1409 13175
rect 1409 13141 1443 13175
rect 1443 13141 1452 13175
rect 1400 13132 1452 13141
rect 9864 13200 9916 13252
rect 2964 13132 3016 13184
rect 9680 13132 9732 13184
rect 4214 13030 4266 13082
rect 4278 13030 4330 13082
rect 4342 13030 4394 13082
rect 4406 13030 4458 13082
rect 4470 13030 4522 13082
rect 7478 13030 7530 13082
rect 7542 13030 7594 13082
rect 7606 13030 7658 13082
rect 7670 13030 7722 13082
rect 7734 13030 7786 13082
rect 3056 12928 3108 12980
rect 9772 12928 9824 12980
rect 1216 12792 1268 12844
rect 2596 12835 2648 12844
rect 2596 12801 2605 12835
rect 2605 12801 2639 12835
rect 2639 12801 2648 12835
rect 2596 12792 2648 12801
rect 9864 12835 9916 12844
rect 1952 12724 2004 12776
rect 9864 12801 9873 12835
rect 9873 12801 9907 12835
rect 9907 12801 9916 12835
rect 9864 12792 9916 12801
rect 10140 12724 10192 12776
rect 2412 12699 2464 12708
rect 2412 12665 2421 12699
rect 2421 12665 2455 12699
rect 2455 12665 2464 12699
rect 2412 12656 2464 12665
rect 2596 12656 2648 12708
rect 2872 12656 2924 12708
rect 3056 12656 3108 12708
rect 2228 12588 2280 12640
rect 10048 12631 10100 12640
rect 10048 12597 10057 12631
rect 10057 12597 10091 12631
rect 10091 12597 10100 12631
rect 10048 12588 10100 12597
rect 2582 12486 2634 12538
rect 2646 12486 2698 12538
rect 2710 12486 2762 12538
rect 2774 12486 2826 12538
rect 2838 12486 2890 12538
rect 5846 12486 5898 12538
rect 5910 12486 5962 12538
rect 5974 12486 6026 12538
rect 6038 12486 6090 12538
rect 6102 12486 6154 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 9238 12486 9290 12538
rect 9302 12486 9354 12538
rect 9366 12486 9418 12538
rect 1400 12427 1452 12436
rect 1400 12393 1409 12427
rect 1409 12393 1443 12427
rect 1443 12393 1452 12427
rect 1400 12384 1452 12393
rect 1768 12384 1820 12436
rect 2228 12384 2280 12436
rect 2964 12316 3016 12368
rect 9956 12384 10008 12436
rect 1492 12180 1544 12232
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 9864 12223 9916 12232
rect 9864 12189 9873 12223
rect 9873 12189 9907 12223
rect 9907 12189 9916 12223
rect 9864 12180 9916 12189
rect 3608 12112 3660 12164
rect 1124 12044 1176 12096
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 4214 11942 4266 11994
rect 4278 11942 4330 11994
rect 4342 11942 4394 11994
rect 4406 11942 4458 11994
rect 4470 11942 4522 11994
rect 7478 11942 7530 11994
rect 7542 11942 7594 11994
rect 7606 11942 7658 11994
rect 7670 11942 7722 11994
rect 7734 11942 7786 11994
rect 3148 11840 3200 11892
rect 9864 11840 9916 11892
rect 1032 11704 1084 11756
rect 1308 11636 1360 11688
rect 2320 11568 2372 11620
rect 3332 11704 3384 11756
rect 1768 11500 1820 11552
rect 2228 11500 2280 11552
rect 2582 11398 2634 11450
rect 2646 11398 2698 11450
rect 2710 11398 2762 11450
rect 2774 11398 2826 11450
rect 2838 11398 2890 11450
rect 5846 11398 5898 11450
rect 5910 11398 5962 11450
rect 5974 11398 6026 11450
rect 6038 11398 6090 11450
rect 6102 11398 6154 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 9238 11398 9290 11450
rect 9302 11398 9354 11450
rect 9366 11398 9418 11450
rect 2044 11296 2096 11348
rect 2228 11296 2280 11348
rect 4804 11296 4856 11348
rect 10048 11271 10100 11280
rect 1676 11203 1728 11212
rect 1676 11169 1685 11203
rect 1685 11169 1719 11203
rect 1719 11169 1728 11203
rect 1676 11160 1728 11169
rect 2044 11160 2096 11212
rect 10048 11237 10057 11271
rect 10057 11237 10091 11271
rect 10091 11237 10100 11271
rect 10048 11228 10100 11237
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 4712 11092 4764 11144
rect 4068 11024 4120 11076
rect 4214 10854 4266 10906
rect 4278 10854 4330 10906
rect 4342 10854 4394 10906
rect 4406 10854 4458 10906
rect 4470 10854 4522 10906
rect 7478 10854 7530 10906
rect 7542 10854 7594 10906
rect 7606 10854 7658 10906
rect 7670 10854 7722 10906
rect 7734 10854 7786 10906
rect 3148 10616 3200 10668
rect 3976 10616 4028 10668
rect 1308 10548 1360 10600
rect 4620 10548 4672 10600
rect 5264 10480 5316 10532
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 2582 10310 2634 10362
rect 2646 10310 2698 10362
rect 2710 10310 2762 10362
rect 2774 10310 2826 10362
rect 2838 10310 2890 10362
rect 5846 10310 5898 10362
rect 5910 10310 5962 10362
rect 5974 10310 6026 10362
rect 6038 10310 6090 10362
rect 6102 10310 6154 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 9238 10310 9290 10362
rect 9302 10310 9354 10362
rect 9366 10310 9418 10362
rect 3424 10208 3476 10260
rect 2136 10072 2188 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 3056 10004 3108 10056
rect 3240 10004 3292 10056
rect 3424 9936 3476 9988
rect 4214 9766 4266 9818
rect 4278 9766 4330 9818
rect 4342 9766 4394 9818
rect 4406 9766 4458 9818
rect 4470 9766 4522 9818
rect 7478 9766 7530 9818
rect 7542 9766 7594 9818
rect 7606 9766 7658 9818
rect 7670 9766 7722 9818
rect 7734 9766 7786 9818
rect 1860 9528 1912 9580
rect 3056 9528 3108 9580
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 3700 9528 3752 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 2872 9435 2924 9444
rect 2872 9401 2881 9435
rect 2881 9401 2915 9435
rect 2915 9401 2924 9435
rect 2872 9392 2924 9401
rect 10048 9435 10100 9444
rect 10048 9401 10057 9435
rect 10057 9401 10091 9435
rect 10091 9401 10100 9435
rect 10048 9392 10100 9401
rect 9864 9324 9916 9376
rect 2582 9222 2634 9274
rect 2646 9222 2698 9274
rect 2710 9222 2762 9274
rect 2774 9222 2826 9274
rect 2838 9222 2890 9274
rect 5846 9222 5898 9274
rect 5910 9222 5962 9274
rect 5974 9222 6026 9274
rect 6038 9222 6090 9274
rect 6102 9222 6154 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 9238 9222 9290 9274
rect 9302 9222 9354 9274
rect 9366 9222 9418 9274
rect 2964 9120 3016 9172
rect 2412 8984 2464 9036
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 3056 8916 3108 8968
rect 3148 8916 3200 8968
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 9864 8959 9916 8968
rect 9864 8925 9873 8959
rect 9873 8925 9907 8959
rect 9907 8925 9916 8959
rect 9864 8916 9916 8925
rect 9864 8780 9916 8832
rect 10048 8823 10100 8832
rect 10048 8789 10057 8823
rect 10057 8789 10091 8823
rect 10091 8789 10100 8823
rect 10048 8780 10100 8789
rect 4214 8678 4266 8730
rect 4278 8678 4330 8730
rect 4342 8678 4394 8730
rect 4406 8678 4458 8730
rect 4470 8678 4522 8730
rect 7478 8678 7530 8730
rect 7542 8678 7594 8730
rect 7606 8678 7658 8730
rect 7670 8678 7722 8730
rect 7734 8678 7786 8730
rect 3056 8619 3108 8628
rect 3056 8585 3065 8619
rect 3065 8585 3099 8619
rect 3099 8585 3108 8619
rect 3056 8576 3108 8585
rect 3700 8576 3752 8628
rect 1584 8508 1636 8560
rect 1768 8440 1820 8492
rect 3240 8440 3292 8492
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 2412 8372 2464 8424
rect 10048 8347 10100 8356
rect 10048 8313 10057 8347
rect 10057 8313 10091 8347
rect 10091 8313 10100 8347
rect 10048 8304 10100 8313
rect 2582 8134 2634 8186
rect 2646 8134 2698 8186
rect 2710 8134 2762 8186
rect 2774 8134 2826 8186
rect 2838 8134 2890 8186
rect 5846 8134 5898 8186
rect 5910 8134 5962 8186
rect 5974 8134 6026 8186
rect 6038 8134 6090 8186
rect 6102 8134 6154 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 9238 8134 9290 8186
rect 9302 8134 9354 8186
rect 9366 8134 9418 8186
rect 1952 7896 2004 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 3056 7828 3108 7880
rect 9864 7692 9916 7744
rect 4214 7590 4266 7642
rect 4278 7590 4330 7642
rect 4342 7590 4394 7642
rect 4406 7590 4458 7642
rect 4470 7590 4522 7642
rect 7478 7590 7530 7642
rect 7542 7590 7594 7642
rect 7606 7590 7658 7642
rect 7670 7590 7722 7642
rect 7734 7590 7786 7642
rect 3516 7488 3568 7540
rect 2504 7420 2556 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 10048 7191 10100 7200
rect 10048 7157 10057 7191
rect 10057 7157 10091 7191
rect 10091 7157 10100 7191
rect 10048 7148 10100 7157
rect 2582 7046 2634 7098
rect 2646 7046 2698 7098
rect 2710 7046 2762 7098
rect 2774 7046 2826 7098
rect 2838 7046 2890 7098
rect 5846 7046 5898 7098
rect 5910 7046 5962 7098
rect 5974 7046 6026 7098
rect 6038 7046 6090 7098
rect 6102 7046 6154 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 9238 7046 9290 7098
rect 9302 7046 9354 7098
rect 9366 7046 9418 7098
rect 3332 6808 3384 6860
rect 1676 6740 1728 6792
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 2228 6715 2280 6724
rect 2228 6681 2237 6715
rect 2237 6681 2271 6715
rect 2271 6681 2280 6715
rect 2228 6672 2280 6681
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 9864 6604 9916 6656
rect 10048 6647 10100 6656
rect 10048 6613 10057 6647
rect 10057 6613 10091 6647
rect 10091 6613 10100 6647
rect 10048 6604 10100 6613
rect 4214 6502 4266 6554
rect 4278 6502 4330 6554
rect 4342 6502 4394 6554
rect 4406 6502 4458 6554
rect 4470 6502 4522 6554
rect 7478 6502 7530 6554
rect 7542 6502 7594 6554
rect 7606 6502 7658 6554
rect 7670 6502 7722 6554
rect 7734 6502 7786 6554
rect 3976 6400 4028 6452
rect 2044 6375 2096 6384
rect 2044 6341 2053 6375
rect 2053 6341 2087 6375
rect 2087 6341 2096 6375
rect 2044 6332 2096 6341
rect 1860 6307 1912 6316
rect 1860 6273 1869 6307
rect 1869 6273 1903 6307
rect 1903 6273 1912 6307
rect 1860 6264 1912 6273
rect 2964 6264 3016 6316
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 3608 6128 3660 6180
rect 2582 5958 2634 6010
rect 2646 5958 2698 6010
rect 2710 5958 2762 6010
rect 2774 5958 2826 6010
rect 2838 5958 2890 6010
rect 5846 5958 5898 6010
rect 5910 5958 5962 6010
rect 5974 5958 6026 6010
rect 6038 5958 6090 6010
rect 6102 5958 6154 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 9238 5958 9290 6010
rect 9302 5958 9354 6010
rect 9366 5958 9418 6010
rect 2320 5856 2372 5908
rect 1492 5720 1544 5772
rect 3424 5720 3476 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 3240 5652 3292 5704
rect 3884 5652 3936 5704
rect 9864 5695 9916 5704
rect 9864 5661 9873 5695
rect 9873 5661 9907 5695
rect 9907 5661 9916 5695
rect 9864 5652 9916 5661
rect 3608 5584 3660 5636
rect 6828 5516 6880 5568
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 4214 5414 4266 5466
rect 4278 5414 4330 5466
rect 4342 5414 4394 5466
rect 4406 5414 4458 5466
rect 4470 5414 4522 5466
rect 7478 5414 7530 5466
rect 7542 5414 7594 5466
rect 7606 5414 7658 5466
rect 7670 5414 7722 5466
rect 7734 5414 7786 5466
rect 1308 5176 1360 5228
rect 3516 5312 3568 5364
rect 3700 5355 3752 5364
rect 3700 5321 3709 5355
rect 3709 5321 3743 5355
rect 3743 5321 3752 5355
rect 3700 5312 3752 5321
rect 3148 5244 3200 5296
rect 3884 5244 3936 5296
rect 3516 5219 3568 5228
rect 3516 5185 3525 5219
rect 3525 5185 3559 5219
rect 3559 5185 3568 5219
rect 3516 5176 3568 5185
rect 6828 5176 6880 5228
rect 2228 5108 2280 5160
rect 2412 5108 2464 5160
rect 5172 5040 5224 5092
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 2582 4870 2634 4922
rect 2646 4870 2698 4922
rect 2710 4870 2762 4922
rect 2774 4870 2826 4922
rect 2838 4870 2890 4922
rect 5846 4870 5898 4922
rect 5910 4870 5962 4922
rect 5974 4870 6026 4922
rect 6038 4870 6090 4922
rect 6102 4870 6154 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 9238 4870 9290 4922
rect 9302 4870 9354 4922
rect 9366 4870 9418 4922
rect 3976 4811 4028 4820
rect 3976 4777 3985 4811
rect 3985 4777 4019 4811
rect 4019 4777 4028 4811
rect 3976 4768 4028 4777
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 1768 4564 1820 4573
rect 3240 4700 3292 4752
rect 1952 4564 2004 4616
rect 3240 4564 3292 4616
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 9864 4607 9916 4616
rect 9864 4573 9873 4607
rect 9873 4573 9907 4607
rect 9907 4573 9916 4607
rect 9864 4564 9916 4573
rect 4620 4496 4672 4548
rect 3332 4428 3384 4480
rect 3792 4428 3844 4480
rect 9772 4428 9824 4480
rect 10048 4471 10100 4480
rect 10048 4437 10057 4471
rect 10057 4437 10091 4471
rect 10091 4437 10100 4471
rect 10048 4428 10100 4437
rect 4214 4326 4266 4378
rect 4278 4326 4330 4378
rect 4342 4326 4394 4378
rect 4406 4326 4458 4378
rect 4470 4326 4522 4378
rect 7478 4326 7530 4378
rect 7542 4326 7594 4378
rect 7606 4326 7658 4378
rect 7670 4326 7722 4378
rect 7734 4326 7786 4378
rect 9864 4224 9916 4276
rect 3148 4088 3200 4140
rect 3976 4088 4028 4140
rect 4068 4088 4120 4140
rect 4620 4088 4672 4140
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 1400 4063 1452 4072
rect 1400 4029 1409 4063
rect 1409 4029 1443 4063
rect 1443 4029 1452 4063
rect 1400 4020 1452 4029
rect 1768 4020 1820 4072
rect 2412 4020 2464 4072
rect 4712 4020 4764 4072
rect 4160 3952 4212 4004
rect 5632 3952 5684 4004
rect 3792 3884 3844 3936
rect 9036 3884 9088 3936
rect 2582 3782 2634 3834
rect 2646 3782 2698 3834
rect 2710 3782 2762 3834
rect 2774 3782 2826 3834
rect 2838 3782 2890 3834
rect 5846 3782 5898 3834
rect 5910 3782 5962 3834
rect 5974 3782 6026 3834
rect 6038 3782 6090 3834
rect 6102 3782 6154 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 9238 3782 9290 3834
rect 9302 3782 9354 3834
rect 9366 3782 9418 3834
rect 3516 3680 3568 3732
rect 10140 3680 10192 3732
rect 4160 3544 4212 3596
rect 4620 3544 4672 3596
rect 1952 3476 2004 3528
rect 2504 3476 2556 3528
rect 3608 3476 3660 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 9772 3476 9824 3528
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 10048 3383 10100 3392
rect 10048 3349 10057 3383
rect 10057 3349 10091 3383
rect 10091 3349 10100 3383
rect 10048 3340 10100 3349
rect 4214 3238 4266 3290
rect 4278 3238 4330 3290
rect 4342 3238 4394 3290
rect 4406 3238 4458 3290
rect 4470 3238 4522 3290
rect 7478 3238 7530 3290
rect 7542 3238 7594 3290
rect 7606 3238 7658 3290
rect 7670 3238 7722 3290
rect 7734 3238 7786 3290
rect 2136 3136 2188 3188
rect 3056 3136 3108 3188
rect 3608 3136 3660 3188
rect 2688 3068 2740 3120
rect 9680 3068 9732 3120
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 2964 3043 3016 3052
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 4436 3000 4488 3009
rect 2504 2932 2556 2984
rect 4160 2932 4212 2984
rect 9036 3000 9088 3052
rect 1676 2864 1728 2916
rect 3424 2796 3476 2848
rect 9496 2796 9548 2848
rect 10048 2839 10100 2848
rect 10048 2805 10057 2839
rect 10057 2805 10091 2839
rect 10091 2805 10100 2839
rect 10048 2796 10100 2805
rect 2582 2694 2634 2746
rect 2646 2694 2698 2746
rect 2710 2694 2762 2746
rect 2774 2694 2826 2746
rect 2838 2694 2890 2746
rect 5846 2694 5898 2746
rect 5910 2694 5962 2746
rect 5974 2694 6026 2746
rect 6038 2694 6090 2746
rect 6102 2694 6154 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 9238 2694 9290 2746
rect 9302 2694 9354 2746
rect 9366 2694 9418 2746
rect 2504 2592 2556 2644
rect 4620 2592 4672 2644
rect 2412 2524 2464 2576
rect 2780 2456 2832 2508
rect 4436 2456 4488 2508
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 4068 2388 4120 2440
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 5632 2388 5684 2440
rect 9680 2388 9732 2440
rect 3332 2320 3384 2372
rect 2228 2252 2280 2304
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 9588 2252 9640 2304
rect 4214 2150 4266 2202
rect 4278 2150 4330 2202
rect 4342 2150 4394 2202
rect 4406 2150 4458 2202
rect 4470 2150 4522 2202
rect 7478 2150 7530 2202
rect 7542 2150 7594 2202
rect 7606 2150 7658 2202
rect 7670 2150 7722 2202
rect 7734 2150 7786 2202
rect 2780 1028 2832 1080
rect 5264 1028 5316 1080
<< metal2 >>
rect 2962 79656 3018 79665
rect 2962 79591 3018 79600
rect 1398 79248 1454 79257
rect 1398 79183 1454 79192
rect 1412 77518 1440 79183
rect 2582 77820 2890 77840
rect 2582 77818 2588 77820
rect 2644 77818 2668 77820
rect 2724 77818 2748 77820
rect 2804 77818 2828 77820
rect 2884 77818 2890 77820
rect 2644 77766 2646 77818
rect 2826 77766 2828 77818
rect 2582 77764 2588 77766
rect 2644 77764 2668 77766
rect 2724 77764 2748 77766
rect 2804 77764 2828 77766
rect 2884 77764 2890 77766
rect 2582 77744 2890 77764
rect 2976 77654 3004 79591
rect 5998 79200 6054 80000
rect 9954 79520 10010 79529
rect 9954 79455 10010 79464
rect 3698 78840 3754 78849
rect 3698 78775 3754 78784
rect 3422 78024 3478 78033
rect 3422 77959 3478 77968
rect 2964 77648 3016 77654
rect 2964 77590 3016 77596
rect 1400 77512 1452 77518
rect 1400 77454 1452 77460
rect 2964 77512 3016 77518
rect 2964 77454 3016 77460
rect 2044 77376 2096 77382
rect 2044 77318 2096 77324
rect 2872 77376 2924 77382
rect 2872 77318 2924 77324
rect 1492 77036 1544 77042
rect 1492 76978 1544 76984
rect 1400 76424 1452 76430
rect 1400 76366 1452 76372
rect 1412 75041 1440 76366
rect 1504 75206 1532 76978
rect 1952 76832 2004 76838
rect 1952 76774 2004 76780
rect 1676 76288 1728 76294
rect 1676 76230 1728 76236
rect 1584 75948 1636 75954
rect 1584 75890 1636 75896
rect 1492 75200 1544 75206
rect 1492 75142 1544 75148
rect 1398 75032 1454 75041
rect 1398 74967 1454 74976
rect 1504 74866 1532 75142
rect 1492 74860 1544 74866
rect 1492 74802 1544 74808
rect 940 74384 992 74390
rect 940 74326 992 74332
rect 756 69760 808 69766
rect 756 69702 808 69708
rect 664 68332 716 68338
rect 664 68274 716 68280
rect 388 65408 440 65414
rect 388 65350 440 65356
rect 296 63980 348 63986
rect 296 63922 348 63928
rect 20 61056 72 61062
rect 20 60998 72 61004
rect 32 50130 60 60998
rect 112 60308 164 60314
rect 112 60250 164 60256
rect 124 51134 152 60250
rect 204 58540 256 58546
rect 204 58482 256 58488
rect 112 51128 164 51134
rect 112 51070 164 51076
rect 110 50416 166 50425
rect 110 50351 112 50360
rect 164 50351 166 50360
rect 112 50322 164 50328
rect 32 50102 152 50130
rect 20 49428 72 49434
rect 20 49370 72 49376
rect 32 45370 60 49370
rect 124 46714 152 50102
rect 112 46708 164 46714
rect 112 46650 164 46656
rect 110 46574 166 46583
rect 110 46509 166 46518
rect 32 45342 152 45370
rect 124 45286 152 45342
rect 20 45280 72 45286
rect 20 45222 72 45228
rect 112 45280 164 45286
rect 112 45222 164 45228
rect 32 40594 60 45222
rect 112 45076 164 45082
rect 112 45018 164 45024
rect 20 40588 72 40594
rect 20 40530 72 40536
rect 20 40452 72 40458
rect 20 40394 72 40400
rect 32 37670 60 40394
rect 20 37664 72 37670
rect 20 37606 72 37612
rect 124 29306 152 45018
rect 216 34134 244 58482
rect 308 45490 336 63922
rect 400 58886 428 65350
rect 572 63164 624 63170
rect 572 63106 624 63112
rect 584 60246 612 63106
rect 572 60240 624 60246
rect 572 60182 624 60188
rect 480 60104 532 60110
rect 480 60046 532 60052
rect 388 58880 440 58886
rect 388 58822 440 58828
rect 388 57860 440 57866
rect 388 57802 440 57808
rect 400 50522 428 57802
rect 492 53417 520 60046
rect 572 59152 624 59158
rect 572 59094 624 59100
rect 584 55554 612 59094
rect 572 55548 624 55554
rect 572 55490 624 55496
rect 676 55078 704 68274
rect 768 60178 796 69702
rect 848 67108 900 67114
rect 848 67050 900 67056
rect 860 60858 888 67050
rect 952 63170 980 74326
rect 1504 74118 1532 74802
rect 1596 74633 1624 75890
rect 1582 74624 1638 74633
rect 1582 74559 1638 74568
rect 1124 74112 1176 74118
rect 1124 74054 1176 74060
rect 1492 74112 1544 74118
rect 1492 74054 1544 74060
rect 1136 72758 1164 74054
rect 1400 73772 1452 73778
rect 1400 73714 1452 73720
rect 1308 73568 1360 73574
rect 1308 73510 1360 73516
rect 1216 73024 1268 73030
rect 1216 72966 1268 72972
rect 1124 72752 1176 72758
rect 1122 72720 1124 72729
rect 1176 72720 1178 72729
rect 1122 72655 1178 72664
rect 1032 71936 1084 71942
rect 1032 71878 1084 71884
rect 1044 66076 1072 71878
rect 1136 71670 1164 72655
rect 1124 71664 1176 71670
rect 1124 71606 1176 71612
rect 1136 70582 1164 71606
rect 1124 70576 1176 70582
rect 1124 70518 1176 70524
rect 1136 69494 1164 70518
rect 1124 69488 1176 69494
rect 1124 69430 1176 69436
rect 1124 69216 1176 69222
rect 1124 69158 1176 69164
rect 1136 66298 1164 69158
rect 1228 66722 1256 72966
rect 1320 72706 1348 73510
rect 1412 72865 1440 73714
rect 1492 73568 1544 73574
rect 1492 73510 1544 73516
rect 1398 72856 1454 72865
rect 1398 72791 1454 72800
rect 1320 72678 1440 72706
rect 1412 71074 1440 72678
rect 1320 71046 1440 71074
rect 1320 69834 1348 71046
rect 1504 70938 1532 73510
rect 1584 73160 1636 73166
rect 1584 73102 1636 73108
rect 1596 72457 1624 73102
rect 1582 72448 1638 72457
rect 1582 72383 1638 72392
rect 1584 72072 1636 72078
rect 1584 72014 1636 72020
rect 1596 71097 1624 72014
rect 1688 71670 1716 76230
rect 1768 76084 1820 76090
rect 1768 76026 1820 76032
rect 1676 71664 1728 71670
rect 1676 71606 1728 71612
rect 1676 71460 1728 71466
rect 1676 71402 1728 71408
rect 1582 71088 1638 71097
rect 1582 71023 1638 71032
rect 1412 70910 1532 70938
rect 1584 70984 1636 70990
rect 1584 70926 1636 70932
rect 1308 69828 1360 69834
rect 1308 69770 1360 69776
rect 1412 68490 1440 70910
rect 1492 70848 1544 70854
rect 1492 70790 1544 70796
rect 1504 70310 1532 70790
rect 1596 70689 1624 70926
rect 1582 70680 1638 70689
rect 1582 70615 1638 70624
rect 1492 70304 1544 70310
rect 1492 70246 1544 70252
rect 1582 70272 1638 70281
rect 1582 70207 1638 70216
rect 1596 69902 1624 70207
rect 1584 69896 1636 69902
rect 1584 69838 1636 69844
rect 1584 69760 1636 69766
rect 1584 69702 1636 69708
rect 1492 69420 1544 69426
rect 1492 69362 1544 69368
rect 1504 68746 1532 69362
rect 1596 69306 1624 69702
rect 1688 69494 1716 71402
rect 1780 70650 1808 76026
rect 1860 75268 1912 75274
rect 1860 75210 1912 75216
rect 1872 74866 1900 75210
rect 1860 74860 1912 74866
rect 1860 74802 1912 74808
rect 1872 74186 1900 74802
rect 1860 74180 1912 74186
rect 1860 74122 1912 74128
rect 1872 72690 1900 74122
rect 1860 72684 1912 72690
rect 1860 72626 1912 72632
rect 1872 72486 1900 72626
rect 1860 72480 1912 72486
rect 1860 72422 1912 72428
rect 1860 72208 1912 72214
rect 1860 72150 1912 72156
rect 1768 70644 1820 70650
rect 1768 70586 1820 70592
rect 1872 70394 1900 72150
rect 1780 70366 1900 70394
rect 1676 69488 1728 69494
rect 1676 69430 1728 69436
rect 1596 69278 1716 69306
rect 1584 68808 1636 68814
rect 1584 68750 1636 68756
rect 1492 68740 1544 68746
rect 1492 68682 1544 68688
rect 1412 68462 1532 68490
rect 1308 68264 1360 68270
rect 1308 68206 1360 68212
rect 1320 67697 1348 68206
rect 1400 67720 1452 67726
rect 1306 67688 1362 67697
rect 1400 67662 1452 67668
rect 1306 67623 1362 67632
rect 1412 67289 1440 67662
rect 1398 67280 1454 67289
rect 1398 67215 1454 67224
rect 1400 67176 1452 67182
rect 1400 67118 1452 67124
rect 1412 66881 1440 67118
rect 1398 66872 1454 66881
rect 1398 66807 1454 66816
rect 1228 66694 1440 66722
rect 1504 66706 1532 68462
rect 1596 68105 1624 68750
rect 1582 68096 1638 68105
rect 1582 68031 1638 68040
rect 1688 67946 1716 69278
rect 1596 67918 1716 67946
rect 1308 66564 1360 66570
rect 1308 66506 1360 66512
rect 1124 66292 1176 66298
rect 1124 66234 1176 66240
rect 1044 66048 1164 66076
rect 1032 65952 1084 65958
rect 1032 65894 1084 65900
rect 940 63164 992 63170
rect 940 63106 992 63112
rect 1044 63050 1072 65894
rect 952 63022 1072 63050
rect 848 60852 900 60858
rect 848 60794 900 60800
rect 952 60738 980 63022
rect 1032 62892 1084 62898
rect 1032 62834 1084 62840
rect 860 60710 980 60738
rect 756 60172 808 60178
rect 756 60114 808 60120
rect 756 59424 808 59430
rect 756 59366 808 59372
rect 768 58614 796 59366
rect 756 58608 808 58614
rect 756 58550 808 58556
rect 756 57928 808 57934
rect 756 57870 808 57876
rect 664 55072 716 55078
rect 664 55014 716 55020
rect 572 54120 624 54126
rect 572 54062 624 54068
rect 478 53408 534 53417
rect 478 53343 534 53352
rect 480 52488 532 52494
rect 480 52430 532 52436
rect 388 50516 440 50522
rect 388 50458 440 50464
rect 388 50380 440 50386
rect 388 50322 440 50328
rect 296 45484 348 45490
rect 296 45426 348 45432
rect 296 45280 348 45286
rect 296 45222 348 45228
rect 308 44441 336 45222
rect 294 44432 350 44441
rect 294 44367 350 44376
rect 296 44328 348 44334
rect 296 44270 348 44276
rect 204 34128 256 34134
rect 204 34070 256 34076
rect 112 29300 164 29306
rect 112 29242 164 29248
rect 308 25770 336 44270
rect 400 34610 428 50322
rect 492 35698 520 52430
rect 584 51270 612 54062
rect 664 53100 716 53106
rect 664 53042 716 53048
rect 572 51264 624 51270
rect 572 51206 624 51212
rect 572 51128 624 51134
rect 572 51070 624 51076
rect 584 45626 612 51070
rect 572 45620 624 45626
rect 572 45562 624 45568
rect 572 45416 624 45422
rect 572 45358 624 45364
rect 584 42838 612 45358
rect 572 42832 624 42838
rect 572 42774 624 42780
rect 572 42084 624 42090
rect 572 42026 624 42032
rect 584 40458 612 42026
rect 572 40452 624 40458
rect 572 40394 624 40400
rect 572 38548 624 38554
rect 572 38490 624 38496
rect 584 37398 612 38490
rect 572 37392 624 37398
rect 572 37334 624 37340
rect 480 35692 532 35698
rect 480 35634 532 35640
rect 388 34604 440 34610
rect 388 34546 440 34552
rect 676 31890 704 53042
rect 768 36242 796 57870
rect 860 57050 888 60710
rect 938 60616 994 60625
rect 938 60551 994 60560
rect 848 57044 900 57050
rect 848 56986 900 56992
rect 848 55752 900 55758
rect 848 55694 900 55700
rect 756 36236 808 36242
rect 756 36178 808 36184
rect 754 32872 810 32881
rect 754 32807 810 32816
rect 664 31884 716 31890
rect 664 31826 716 31832
rect 664 31340 716 31346
rect 664 31282 716 31288
rect 676 28150 704 31282
rect 768 29850 796 32807
rect 860 32026 888 55694
rect 952 50250 980 60551
rect 1044 50538 1072 62834
rect 1136 62218 1164 66048
rect 1320 66026 1348 66506
rect 1308 66020 1360 66026
rect 1308 65962 1360 65968
rect 1320 65006 1348 65962
rect 1308 65000 1360 65006
rect 1308 64942 1360 64948
rect 1320 64054 1348 64942
rect 1412 64938 1440 66694
rect 1492 66700 1544 66706
rect 1492 66642 1544 66648
rect 1596 66298 1624 67918
rect 1676 67720 1728 67726
rect 1674 67688 1676 67697
rect 1728 67688 1730 67697
rect 1674 67623 1730 67632
rect 1676 67040 1728 67046
rect 1676 66982 1728 66988
rect 1492 66292 1544 66298
rect 1492 66234 1544 66240
rect 1584 66292 1636 66298
rect 1584 66234 1636 66240
rect 1504 65226 1532 66234
rect 1582 66192 1638 66201
rect 1582 66127 1584 66136
rect 1636 66127 1638 66136
rect 1584 66098 1636 66104
rect 1582 66056 1638 66065
rect 1582 65991 1638 66000
rect 1596 65550 1624 65991
rect 1584 65544 1636 65550
rect 1584 65486 1636 65492
rect 1504 65198 1624 65226
rect 1492 65136 1544 65142
rect 1492 65078 1544 65084
rect 1504 64977 1532 65078
rect 1490 64968 1546 64977
rect 1400 64932 1452 64938
rect 1490 64903 1546 64912
rect 1400 64874 1452 64880
rect 1308 64048 1360 64054
rect 1308 63990 1360 63996
rect 1596 63968 1624 65198
rect 1412 63940 1624 63968
rect 1412 63322 1440 63940
rect 1688 63900 1716 66982
rect 1780 65618 1808 70366
rect 1860 70304 1912 70310
rect 1860 70246 1912 70252
rect 1872 67046 1900 70246
rect 1860 67040 1912 67046
rect 1860 66982 1912 66988
rect 1768 65612 1820 65618
rect 1768 65554 1820 65560
rect 1860 65408 1912 65414
rect 1860 65350 1912 65356
rect 1872 65006 1900 65350
rect 1860 65000 1912 65006
rect 1860 64942 1912 64948
rect 1768 64592 1820 64598
rect 1768 64534 1820 64540
rect 1228 63294 1440 63322
rect 1504 63872 1716 63900
rect 1124 62212 1176 62218
rect 1124 62154 1176 62160
rect 1124 61124 1176 61130
rect 1124 61066 1176 61072
rect 1136 59770 1164 61066
rect 1228 60858 1256 63294
rect 1400 63232 1452 63238
rect 1400 63174 1452 63180
rect 1412 62121 1440 63174
rect 1398 62112 1454 62121
rect 1398 62047 1454 62056
rect 1504 61962 1532 63872
rect 1584 63776 1636 63782
rect 1584 63718 1636 63724
rect 1596 63073 1624 63718
rect 1676 63504 1728 63510
rect 1674 63472 1676 63481
rect 1728 63472 1730 63481
rect 1674 63407 1730 63416
rect 1676 63368 1728 63374
rect 1676 63310 1728 63316
rect 1582 63064 1638 63073
rect 1582 62999 1638 63008
rect 1584 62688 1636 62694
rect 1584 62630 1636 62636
rect 1412 61934 1532 61962
rect 1216 60852 1268 60858
rect 1216 60794 1268 60800
rect 1216 60512 1268 60518
rect 1216 60454 1268 60460
rect 1124 59764 1176 59770
rect 1124 59706 1176 59712
rect 1124 59628 1176 59634
rect 1124 59570 1176 59576
rect 1136 58993 1164 59570
rect 1122 58984 1178 58993
rect 1122 58919 1178 58928
rect 1122 58848 1178 58857
rect 1122 58783 1178 58792
rect 1136 56409 1164 58783
rect 1228 56594 1256 60454
rect 1308 60240 1360 60246
rect 1308 60182 1360 60188
rect 1320 56658 1348 60182
rect 1412 58954 1440 61934
rect 1492 61804 1544 61810
rect 1492 61746 1544 61752
rect 1504 61130 1532 61746
rect 1596 61441 1624 62630
rect 1688 62257 1716 63310
rect 1674 62248 1730 62257
rect 1674 62183 1730 62192
rect 1780 62098 1808 64534
rect 1872 64394 1900 64942
rect 1860 64388 1912 64394
rect 1860 64330 1912 64336
rect 1872 62150 1900 64330
rect 1688 62070 1808 62098
rect 1860 62144 1912 62150
rect 1860 62086 1912 62092
rect 1582 61432 1638 61441
rect 1582 61367 1638 61376
rect 1688 61130 1716 62070
rect 1768 61804 1820 61810
rect 1768 61746 1820 61752
rect 1780 61305 1808 61746
rect 1860 61600 1912 61606
rect 1860 61542 1912 61548
rect 1766 61296 1822 61305
rect 1766 61231 1822 61240
rect 1780 61198 1808 61231
rect 1768 61192 1820 61198
rect 1768 61134 1820 61140
rect 1492 61124 1544 61130
rect 1492 61066 1544 61072
rect 1676 61124 1728 61130
rect 1676 61066 1728 61072
rect 1676 60852 1728 60858
rect 1676 60794 1728 60800
rect 1492 60784 1544 60790
rect 1492 60726 1544 60732
rect 1400 58948 1452 58954
rect 1400 58890 1452 58896
rect 1400 58336 1452 58342
rect 1400 58278 1452 58284
rect 1412 57497 1440 58278
rect 1398 57488 1454 57497
rect 1398 57423 1454 57432
rect 1320 56630 1440 56658
rect 1228 56566 1348 56594
rect 1122 56400 1178 56409
rect 1122 56335 1178 56344
rect 1216 56296 1268 56302
rect 1216 56238 1268 56244
rect 1124 55072 1176 55078
rect 1124 55014 1176 55020
rect 1136 51066 1164 55014
rect 1228 51074 1256 56238
rect 1320 55350 1348 56566
rect 1308 55344 1360 55350
rect 1308 55286 1360 55292
rect 1306 55176 1362 55185
rect 1306 55111 1308 55120
rect 1360 55111 1362 55120
rect 1308 55082 1360 55088
rect 1412 54330 1440 56630
rect 1504 56370 1532 60726
rect 1584 60512 1636 60518
rect 1584 60454 1636 60460
rect 1596 59129 1624 60454
rect 1582 59120 1638 59129
rect 1582 59055 1638 59064
rect 1584 59016 1636 59022
rect 1584 58958 1636 58964
rect 1596 58682 1624 58958
rect 1584 58676 1636 58682
rect 1584 58618 1636 58624
rect 1584 57792 1636 57798
rect 1584 57734 1636 57740
rect 1596 57089 1624 57734
rect 1582 57080 1638 57089
rect 1582 57015 1638 57024
rect 1688 56846 1716 60794
rect 1768 60716 1820 60722
rect 1768 60658 1820 60664
rect 1780 60314 1808 60658
rect 1768 60308 1820 60314
rect 1768 60250 1820 60256
rect 1768 60036 1820 60042
rect 1768 59978 1820 59984
rect 1780 57594 1808 59978
rect 1768 57588 1820 57594
rect 1768 57530 1820 57536
rect 1768 57452 1820 57458
rect 1768 57394 1820 57400
rect 1780 56846 1808 57394
rect 1676 56840 1728 56846
rect 1676 56782 1728 56788
rect 1768 56840 1820 56846
rect 1768 56782 1820 56788
rect 1584 56772 1636 56778
rect 1584 56714 1636 56720
rect 1492 56364 1544 56370
rect 1492 56306 1544 56312
rect 1596 55706 1624 56714
rect 1674 56672 1730 56681
rect 1674 56607 1730 56616
rect 1688 56506 1716 56607
rect 1676 56500 1728 56506
rect 1676 56442 1728 56448
rect 1768 56432 1820 56438
rect 1768 56374 1820 56380
rect 1676 56364 1728 56370
rect 1676 56306 1728 56312
rect 1504 55678 1624 55706
rect 1504 55162 1532 55678
rect 1584 55616 1636 55622
rect 1584 55558 1636 55564
rect 1596 55457 1624 55558
rect 1582 55448 1638 55457
rect 1582 55383 1638 55392
rect 1504 55134 1624 55162
rect 1492 55072 1544 55078
rect 1492 55014 1544 55020
rect 1400 54324 1452 54330
rect 1400 54266 1452 54272
rect 1504 54097 1532 55014
rect 1596 54602 1624 55134
rect 1688 54806 1716 56306
rect 1780 55457 1808 56374
rect 1766 55448 1822 55457
rect 1766 55383 1822 55392
rect 1768 55276 1820 55282
rect 1768 55218 1820 55224
rect 1676 54800 1728 54806
rect 1676 54742 1728 54748
rect 1584 54596 1636 54602
rect 1584 54538 1636 54544
rect 1596 54194 1624 54538
rect 1780 54369 1808 55218
rect 1766 54360 1822 54369
rect 1676 54324 1728 54330
rect 1766 54295 1822 54304
rect 1676 54266 1728 54272
rect 1584 54188 1636 54194
rect 1584 54130 1636 54136
rect 1490 54088 1546 54097
rect 1308 54052 1360 54058
rect 1490 54023 1546 54032
rect 1308 53994 1360 54000
rect 1320 51649 1348 53994
rect 1400 53440 1452 53446
rect 1400 53382 1452 53388
rect 1412 52737 1440 53382
rect 1584 52896 1636 52902
rect 1584 52838 1636 52844
rect 1398 52728 1454 52737
rect 1398 52663 1454 52672
rect 1492 52352 1544 52358
rect 1596 52329 1624 52838
rect 1492 52294 1544 52300
rect 1582 52320 1638 52329
rect 1400 52012 1452 52018
rect 1400 51954 1452 51960
rect 1306 51640 1362 51649
rect 1306 51575 1362 51584
rect 1308 51536 1360 51542
rect 1308 51478 1360 51484
rect 1320 51241 1348 51478
rect 1306 51232 1362 51241
rect 1306 51167 1362 51176
rect 1124 51060 1176 51066
rect 1228 51046 1348 51074
rect 1124 51002 1176 51008
rect 1214 50960 1270 50969
rect 1214 50895 1270 50904
rect 1124 50788 1176 50794
rect 1124 50730 1176 50736
rect 1136 50697 1164 50730
rect 1122 50688 1178 50697
rect 1122 50623 1178 50632
rect 1044 50510 1164 50538
rect 1032 50448 1084 50454
rect 1032 50390 1084 50396
rect 940 50244 992 50250
rect 940 50186 992 50192
rect 1044 50130 1072 50390
rect 952 50102 1072 50130
rect 952 38962 980 50102
rect 1136 49994 1164 50510
rect 1044 49966 1164 49994
rect 1044 45626 1072 49966
rect 1122 49872 1178 49881
rect 1122 49807 1124 49816
rect 1176 49807 1178 49816
rect 1124 49778 1176 49784
rect 1124 49632 1176 49638
rect 1124 49574 1176 49580
rect 1136 48550 1164 49574
rect 1124 48544 1176 48550
rect 1124 48486 1176 48492
rect 1122 48376 1178 48385
rect 1122 48311 1178 48320
rect 1032 45620 1084 45626
rect 1032 45562 1084 45568
rect 1032 45484 1084 45490
rect 1032 45426 1084 45432
rect 1044 41546 1072 45426
rect 1032 41540 1084 41546
rect 1032 41482 1084 41488
rect 1030 41440 1086 41449
rect 1030 41375 1086 41384
rect 940 38956 992 38962
rect 940 38898 992 38904
rect 938 38584 994 38593
rect 938 38519 994 38528
rect 952 38418 980 38519
rect 940 38412 992 38418
rect 940 38354 992 38360
rect 940 38208 992 38214
rect 940 38150 992 38156
rect 952 36961 980 38150
rect 938 36952 994 36961
rect 938 36887 994 36896
rect 940 32360 992 32366
rect 940 32302 992 32308
rect 848 32020 900 32026
rect 848 31962 900 31968
rect 848 31272 900 31278
rect 848 31214 900 31220
rect 860 30054 888 31214
rect 848 30048 900 30054
rect 848 29990 900 29996
rect 756 29844 808 29850
rect 756 29786 808 29792
rect 664 28144 716 28150
rect 664 28086 716 28092
rect 296 25764 348 25770
rect 296 25706 348 25712
rect 952 22302 980 32302
rect 1044 27470 1072 41375
rect 1136 41206 1164 48311
rect 1124 41200 1176 41206
rect 1124 41142 1176 41148
rect 1124 39432 1176 39438
rect 1124 39374 1176 39380
rect 1136 39273 1164 39374
rect 1122 39264 1178 39273
rect 1122 39199 1178 39208
rect 1124 39092 1176 39098
rect 1124 39034 1176 39040
rect 1136 38729 1164 39034
rect 1122 38720 1178 38729
rect 1122 38655 1178 38664
rect 1228 38570 1256 50895
rect 1320 45082 1348 51046
rect 1412 50969 1440 51954
rect 1398 50960 1454 50969
rect 1398 50895 1454 50904
rect 1504 50794 1532 52294
rect 1582 52255 1638 52264
rect 1582 52184 1638 52193
rect 1582 52119 1584 52128
rect 1636 52119 1638 52128
rect 1584 52090 1636 52096
rect 1688 52034 1716 54266
rect 1768 53984 1820 53990
rect 1768 53926 1820 53932
rect 1596 52006 1716 52034
rect 1596 51388 1624 52006
rect 1676 51808 1728 51814
rect 1676 51750 1728 51756
rect 1688 51542 1716 51750
rect 1676 51536 1728 51542
rect 1676 51478 1728 51484
rect 1596 51360 1716 51388
rect 1780 51377 1808 53926
rect 1584 51264 1636 51270
rect 1584 51206 1636 51212
rect 1492 50788 1544 50794
rect 1492 50730 1544 50736
rect 1400 50720 1452 50726
rect 1596 50674 1624 51206
rect 1688 51105 1716 51360
rect 1766 51368 1822 51377
rect 1766 51303 1822 51312
rect 1766 51232 1822 51241
rect 1766 51167 1822 51176
rect 1674 51096 1730 51105
rect 1674 51031 1730 51040
rect 1780 50930 1808 51167
rect 1768 50924 1820 50930
rect 1768 50866 1820 50872
rect 1400 50662 1452 50668
rect 1412 49366 1440 50662
rect 1504 50646 1624 50674
rect 1504 50289 1532 50646
rect 1584 50516 1636 50522
rect 1584 50458 1636 50464
rect 1596 50318 1624 50458
rect 1674 50416 1730 50425
rect 1674 50351 1730 50360
rect 1584 50312 1636 50318
rect 1490 50280 1546 50289
rect 1584 50254 1636 50260
rect 1490 50215 1546 50224
rect 1492 50176 1544 50182
rect 1492 50118 1544 50124
rect 1400 49360 1452 49366
rect 1400 49302 1452 49308
rect 1400 49088 1452 49094
rect 1400 49030 1452 49036
rect 1412 48521 1440 49030
rect 1398 48512 1454 48521
rect 1398 48447 1454 48456
rect 1400 48136 1452 48142
rect 1400 48078 1452 48084
rect 1412 47433 1440 48078
rect 1504 47546 1532 50118
rect 1596 49842 1624 50254
rect 1688 49910 1716 50351
rect 1780 50318 1808 50866
rect 1768 50312 1820 50318
rect 1768 50254 1820 50260
rect 1676 49904 1728 49910
rect 1676 49846 1728 49852
rect 1780 49842 1808 50254
rect 1584 49836 1636 49842
rect 1584 49778 1636 49784
rect 1768 49836 1820 49842
rect 1768 49778 1820 49784
rect 1768 49700 1820 49706
rect 1768 49642 1820 49648
rect 1676 49360 1728 49366
rect 1676 49302 1728 49308
rect 1584 48544 1636 48550
rect 1584 48486 1636 48492
rect 1596 48113 1624 48486
rect 1582 48104 1638 48113
rect 1582 48039 1638 48048
rect 1584 48000 1636 48006
rect 1584 47942 1636 47948
rect 1596 47705 1624 47942
rect 1582 47696 1638 47705
rect 1582 47631 1638 47640
rect 1504 47518 1624 47546
rect 1492 47456 1544 47462
rect 1398 47424 1454 47433
rect 1492 47398 1544 47404
rect 1398 47359 1454 47368
rect 1504 47122 1532 47398
rect 1492 47116 1544 47122
rect 1492 47058 1544 47064
rect 1492 46980 1544 46986
rect 1492 46922 1544 46928
rect 1400 46708 1452 46714
rect 1400 46650 1452 46656
rect 1412 46617 1440 46650
rect 1398 46608 1454 46617
rect 1398 46543 1454 46552
rect 1400 46368 1452 46374
rect 1400 46310 1452 46316
rect 1412 46034 1440 46310
rect 1400 46028 1452 46034
rect 1400 45970 1452 45976
rect 1398 45656 1454 45665
rect 1398 45591 1454 45600
rect 1308 45076 1360 45082
rect 1308 45018 1360 45024
rect 1412 44962 1440 45591
rect 1504 45490 1532 46922
rect 1596 45914 1624 47518
rect 1688 46986 1716 49302
rect 1780 48346 1808 49642
rect 1768 48340 1820 48346
rect 1768 48282 1820 48288
rect 1766 48240 1822 48249
rect 1766 48175 1822 48184
rect 1780 47122 1808 48175
rect 1768 47116 1820 47122
rect 1768 47058 1820 47064
rect 1676 46980 1728 46986
rect 1676 46922 1728 46928
rect 1674 46880 1730 46889
rect 1674 46815 1730 46824
rect 1688 46034 1716 46815
rect 1768 46708 1820 46714
rect 1768 46650 1820 46656
rect 1676 46028 1728 46034
rect 1676 45970 1728 45976
rect 1596 45886 1716 45914
rect 1492 45484 1544 45490
rect 1492 45426 1544 45432
rect 1490 45384 1546 45393
rect 1490 45319 1546 45328
rect 1320 44934 1440 44962
rect 1320 43246 1348 44934
rect 1400 44872 1452 44878
rect 1400 44814 1452 44820
rect 1412 44305 1440 44814
rect 1398 44296 1454 44305
rect 1398 44231 1454 44240
rect 1504 44180 1532 45319
rect 1582 45112 1638 45121
rect 1582 45047 1584 45056
rect 1636 45047 1638 45056
rect 1584 45018 1636 45024
rect 1582 44704 1638 44713
rect 1582 44639 1638 44648
rect 1596 44538 1624 44639
rect 1584 44532 1636 44538
rect 1584 44474 1636 44480
rect 1412 44152 1532 44180
rect 1582 44160 1638 44169
rect 1308 43240 1360 43246
rect 1308 43182 1360 43188
rect 1306 42800 1362 42809
rect 1306 42735 1362 42744
rect 1320 42294 1348 42735
rect 1308 42288 1360 42294
rect 1308 42230 1360 42236
rect 1412 42242 1440 44152
rect 1582 44095 1638 44104
rect 1492 43716 1544 43722
rect 1492 43658 1544 43664
rect 1504 43314 1532 43658
rect 1596 43450 1624 44095
rect 1584 43444 1636 43450
rect 1584 43386 1636 43392
rect 1688 43330 1716 45886
rect 1492 43308 1544 43314
rect 1492 43250 1544 43256
rect 1596 43302 1716 43330
rect 1492 43172 1544 43178
rect 1492 43114 1544 43120
rect 1504 43081 1532 43114
rect 1490 43072 1546 43081
rect 1490 43007 1546 43016
rect 1492 42696 1544 42702
rect 1492 42638 1544 42644
rect 1504 42362 1532 42638
rect 1492 42356 1544 42362
rect 1492 42298 1544 42304
rect 1412 42214 1532 42242
rect 1400 42152 1452 42158
rect 1400 42094 1452 42100
rect 1308 41608 1360 41614
rect 1306 41576 1308 41585
rect 1360 41576 1362 41585
rect 1306 41511 1362 41520
rect 1306 41440 1362 41449
rect 1306 41375 1362 41384
rect 1320 39284 1348 41375
rect 1412 41274 1440 42094
rect 1400 41268 1452 41274
rect 1400 41210 1452 41216
rect 1400 41132 1452 41138
rect 1400 41074 1452 41080
rect 1412 39409 1440 41074
rect 1398 39400 1454 39409
rect 1398 39335 1454 39344
rect 1320 39256 1440 39284
rect 1306 38856 1362 38865
rect 1306 38791 1362 38800
rect 1320 38593 1348 38791
rect 1136 38542 1256 38570
rect 1306 38584 1362 38593
rect 1136 38350 1164 38542
rect 1412 38554 1440 39256
rect 1504 38554 1532 42214
rect 1596 38593 1624 43302
rect 1676 43240 1728 43246
rect 1676 43182 1728 43188
rect 1688 41449 1716 43182
rect 1780 42401 1808 46650
rect 1872 46186 1900 61542
rect 1964 61033 1992 76774
rect 2056 75970 2084 77318
rect 2320 77036 2372 77042
rect 2320 76978 2372 76984
rect 2504 77036 2556 77042
rect 2504 76978 2556 76984
rect 2056 75942 2176 75970
rect 2044 75880 2096 75886
rect 2044 75822 2096 75828
rect 2056 75206 2084 75822
rect 2044 75200 2096 75206
rect 2044 75142 2096 75148
rect 2044 74724 2096 74730
rect 2044 74666 2096 74672
rect 2056 71466 2084 74666
rect 2044 71460 2096 71466
rect 2044 71402 2096 71408
rect 2044 70508 2096 70514
rect 2044 70450 2096 70456
rect 2056 69873 2084 70450
rect 2042 69864 2098 69873
rect 2042 69799 2098 69808
rect 2044 69760 2096 69766
rect 2044 69702 2096 69708
rect 1950 61024 2006 61033
rect 1950 60959 2006 60968
rect 1952 60852 2004 60858
rect 1952 60794 2004 60800
rect 1964 59226 1992 60794
rect 2056 59974 2084 69702
rect 2148 61606 2176 75942
rect 2332 75818 2360 76978
rect 2412 76832 2464 76838
rect 2412 76774 2464 76780
rect 2320 75812 2372 75818
rect 2320 75754 2372 75760
rect 2332 75342 2360 75754
rect 2320 75336 2372 75342
rect 2320 75278 2372 75284
rect 2320 74656 2372 74662
rect 2320 74598 2372 74604
rect 2228 73772 2280 73778
rect 2228 73714 2280 73720
rect 2240 73273 2268 73714
rect 2226 73264 2282 73273
rect 2332 73234 2360 74598
rect 2226 73199 2282 73208
rect 2320 73228 2372 73234
rect 2320 73170 2372 73176
rect 2228 72072 2280 72078
rect 2228 72014 2280 72020
rect 2240 71641 2268 72014
rect 2320 71936 2372 71942
rect 2320 71878 2372 71884
rect 2226 71632 2282 71641
rect 2226 71567 2282 71576
rect 2228 69896 2280 69902
rect 2228 69838 2280 69844
rect 2240 69057 2268 69838
rect 2226 69048 2282 69057
rect 2226 68983 2282 68992
rect 2228 68672 2280 68678
rect 2228 68614 2280 68620
rect 2240 67425 2268 68614
rect 2226 67416 2282 67425
rect 2226 67351 2282 67360
rect 2228 67312 2280 67318
rect 2228 67254 2280 67260
rect 2240 64598 2268 67254
rect 2228 64592 2280 64598
rect 2228 64534 2280 64540
rect 2228 64456 2280 64462
rect 2332 64444 2360 71878
rect 2424 71738 2452 76774
rect 2516 75857 2544 76978
rect 2884 76820 2912 77318
rect 2976 77081 3004 77454
rect 3148 77376 3200 77382
rect 3148 77318 3200 77324
rect 2962 77072 3018 77081
rect 2962 77007 3018 77016
rect 3056 76968 3108 76974
rect 3056 76910 3108 76916
rect 3068 76838 3096 76910
rect 3056 76832 3108 76838
rect 2884 76792 3004 76820
rect 2582 76732 2890 76752
rect 2582 76730 2588 76732
rect 2644 76730 2668 76732
rect 2724 76730 2748 76732
rect 2804 76730 2828 76732
rect 2884 76730 2890 76732
rect 2644 76678 2646 76730
rect 2826 76678 2828 76730
rect 2582 76676 2588 76678
rect 2644 76676 2668 76678
rect 2724 76676 2748 76678
rect 2804 76676 2828 76678
rect 2884 76676 2890 76678
rect 2582 76656 2890 76676
rect 2780 76424 2832 76430
rect 2780 76366 2832 76372
rect 2596 76288 2648 76294
rect 2596 76230 2648 76236
rect 2608 75954 2636 76230
rect 2792 75954 2820 76366
rect 2596 75948 2648 75954
rect 2596 75890 2648 75896
rect 2780 75948 2832 75954
rect 2780 75890 2832 75896
rect 2502 75848 2558 75857
rect 2792 75818 2820 75890
rect 2502 75783 2558 75792
rect 2780 75812 2832 75818
rect 2780 75754 2832 75760
rect 2582 75644 2890 75664
rect 2582 75642 2588 75644
rect 2644 75642 2668 75644
rect 2724 75642 2748 75644
rect 2804 75642 2828 75644
rect 2884 75642 2890 75644
rect 2644 75590 2646 75642
rect 2826 75590 2828 75642
rect 2582 75588 2588 75590
rect 2644 75588 2668 75590
rect 2724 75588 2748 75590
rect 2804 75588 2828 75590
rect 2884 75588 2890 75590
rect 2582 75568 2890 75588
rect 2504 75472 2556 75478
rect 2504 75414 2556 75420
rect 2516 75041 2544 75414
rect 2976 75274 3004 76792
rect 3056 76774 3108 76780
rect 3056 76560 3108 76566
rect 3056 76502 3108 76508
rect 2964 75268 3016 75274
rect 2964 75210 3016 75216
rect 2502 75032 2558 75041
rect 2502 74967 2558 74976
rect 2964 74860 3016 74866
rect 2964 74802 3016 74808
rect 2582 74556 2890 74576
rect 2582 74554 2588 74556
rect 2644 74554 2668 74556
rect 2724 74554 2748 74556
rect 2804 74554 2828 74556
rect 2884 74554 2890 74556
rect 2644 74502 2646 74554
rect 2826 74502 2828 74554
rect 2582 74500 2588 74502
rect 2644 74500 2668 74502
rect 2724 74500 2748 74502
rect 2804 74500 2828 74502
rect 2884 74500 2890 74502
rect 2582 74480 2890 74500
rect 2976 74089 3004 74802
rect 2962 74080 3018 74089
rect 2962 74015 3018 74024
rect 2872 73772 2924 73778
rect 2872 73714 2924 73720
rect 2884 73681 2912 73714
rect 2870 73672 2926 73681
rect 2870 73607 2926 73616
rect 2582 73468 2890 73488
rect 2582 73466 2588 73468
rect 2644 73466 2668 73468
rect 2724 73466 2748 73468
rect 2804 73466 2828 73468
rect 2884 73466 2890 73468
rect 2644 73414 2646 73466
rect 2826 73414 2828 73466
rect 2582 73412 2588 73414
rect 2644 73412 2668 73414
rect 2724 73412 2748 73414
rect 2804 73412 2828 73414
rect 2884 73412 2890 73414
rect 2582 73392 2890 73412
rect 2780 73092 2832 73098
rect 2780 73034 2832 73040
rect 2686 72720 2742 72729
rect 2792 72690 2820 73034
rect 2686 72655 2688 72664
rect 2740 72655 2742 72664
rect 2780 72684 2832 72690
rect 2688 72626 2740 72632
rect 2780 72626 2832 72632
rect 2964 72684 3016 72690
rect 2964 72626 3016 72632
rect 2976 72486 3004 72626
rect 2964 72480 3016 72486
rect 2964 72422 3016 72428
rect 2582 72380 2890 72400
rect 2582 72378 2588 72380
rect 2644 72378 2668 72380
rect 2724 72378 2748 72380
rect 2804 72378 2828 72380
rect 2884 72378 2890 72380
rect 2644 72326 2646 72378
rect 2826 72326 2828 72378
rect 2582 72324 2588 72326
rect 2644 72324 2668 72326
rect 2724 72324 2748 72326
rect 2804 72324 2828 72326
rect 2884 72324 2890 72326
rect 2582 72304 2890 72324
rect 2872 72072 2924 72078
rect 2870 72040 2872 72049
rect 2924 72040 2926 72049
rect 2870 71975 2926 71984
rect 2596 71936 2648 71942
rect 2596 71878 2648 71884
rect 2412 71732 2464 71738
rect 2412 71674 2464 71680
rect 2608 71602 2636 71878
rect 2976 71602 3004 72422
rect 2412 71596 2464 71602
rect 2412 71538 2464 71544
rect 2596 71596 2648 71602
rect 2596 71538 2648 71544
rect 2964 71596 3016 71602
rect 2964 71538 3016 71544
rect 2424 70582 2452 71538
rect 2582 71292 2890 71312
rect 2582 71290 2588 71292
rect 2644 71290 2668 71292
rect 2724 71290 2748 71292
rect 2804 71290 2828 71292
rect 2884 71290 2890 71292
rect 2644 71238 2646 71290
rect 2826 71238 2828 71290
rect 2582 71236 2588 71238
rect 2644 71236 2668 71238
rect 2724 71236 2748 71238
rect 2804 71236 2828 71238
rect 2884 71236 2890 71238
rect 2582 71216 2890 71236
rect 2976 70582 3004 71538
rect 2412 70576 2464 70582
rect 2412 70518 2464 70524
rect 2964 70576 3016 70582
rect 2964 70518 3016 70524
rect 2412 70304 2464 70310
rect 2412 70246 2464 70252
rect 2424 67318 2452 70246
rect 2582 70204 2890 70224
rect 2582 70202 2588 70204
rect 2644 70202 2668 70204
rect 2724 70202 2748 70204
rect 2804 70202 2828 70204
rect 2884 70202 2890 70204
rect 2644 70150 2646 70202
rect 2826 70150 2828 70202
rect 2582 70148 2588 70150
rect 2644 70148 2668 70150
rect 2724 70148 2748 70150
rect 2804 70148 2828 70150
rect 2884 70148 2890 70150
rect 2582 70128 2890 70148
rect 2872 69896 2924 69902
rect 2872 69838 2924 69844
rect 2688 69760 2740 69766
rect 2688 69702 2740 69708
rect 2700 69329 2728 69702
rect 2884 69465 2912 69838
rect 2976 69578 3004 70518
rect 3068 69766 3096 76502
rect 3160 75954 3188 77318
rect 3436 77042 3464 77959
rect 3516 77716 3568 77722
rect 3516 77658 3568 77664
rect 3332 77036 3384 77042
rect 3332 76978 3384 76984
rect 3424 77036 3476 77042
rect 3424 76978 3476 76984
rect 3240 76832 3292 76838
rect 3240 76774 3292 76780
rect 3252 76362 3280 76774
rect 3344 76537 3372 76978
rect 3330 76528 3386 76537
rect 3330 76463 3386 76472
rect 3240 76356 3292 76362
rect 3240 76298 3292 76304
rect 3528 76242 3556 77658
rect 3712 77110 3740 78775
rect 9586 78704 9642 78713
rect 9586 78639 9642 78648
rect 4066 78432 4122 78441
rect 4066 78367 4122 78376
rect 3974 77616 4030 77625
rect 3974 77551 4030 77560
rect 3988 77518 4016 77551
rect 4080 77518 4108 78367
rect 9494 78024 9550 78033
rect 9494 77959 9550 77968
rect 5846 77820 6154 77840
rect 5846 77818 5852 77820
rect 5908 77818 5932 77820
rect 5988 77818 6012 77820
rect 6068 77818 6092 77820
rect 6148 77818 6154 77820
rect 5908 77766 5910 77818
rect 6090 77766 6092 77818
rect 5846 77764 5852 77766
rect 5908 77764 5932 77766
rect 5988 77764 6012 77766
rect 6068 77764 6092 77766
rect 6148 77764 6154 77766
rect 5846 77744 6154 77764
rect 9110 77820 9418 77840
rect 9110 77818 9116 77820
rect 9172 77818 9196 77820
rect 9252 77818 9276 77820
rect 9332 77818 9356 77820
rect 9412 77818 9418 77820
rect 9172 77766 9174 77818
rect 9354 77766 9356 77818
rect 9110 77764 9116 77766
rect 9172 77764 9196 77766
rect 9252 77764 9276 77766
rect 9332 77764 9356 77766
rect 9412 77764 9418 77766
rect 9110 77744 9418 77764
rect 3976 77512 4028 77518
rect 3976 77454 4028 77460
rect 4068 77512 4120 77518
rect 4068 77454 4120 77460
rect 9404 77512 9456 77518
rect 9404 77454 9456 77460
rect 7840 77444 7892 77450
rect 7840 77386 7892 77392
rect 3884 77376 3936 77382
rect 3884 77318 3936 77324
rect 3700 77104 3752 77110
rect 3700 77046 3752 77052
rect 3608 76968 3660 76974
rect 3608 76910 3660 76916
rect 3252 76214 3556 76242
rect 3148 75948 3200 75954
rect 3148 75890 3200 75896
rect 3148 73568 3200 73574
rect 3148 73510 3200 73516
rect 3056 69760 3108 69766
rect 3056 69702 3108 69708
rect 2976 69550 3096 69578
rect 3068 69494 3096 69550
rect 3056 69488 3108 69494
rect 2870 69456 2926 69465
rect 3056 69430 3108 69436
rect 2870 69391 2926 69400
rect 2964 69420 3016 69426
rect 2964 69362 3016 69368
rect 2686 69320 2742 69329
rect 2686 69255 2742 69264
rect 2582 69116 2890 69136
rect 2582 69114 2588 69116
rect 2644 69114 2668 69116
rect 2724 69114 2748 69116
rect 2804 69114 2828 69116
rect 2884 69114 2890 69116
rect 2644 69062 2646 69114
rect 2826 69062 2828 69114
rect 2582 69060 2588 69062
rect 2644 69060 2668 69062
rect 2724 69060 2748 69062
rect 2804 69060 2828 69062
rect 2884 69060 2890 69062
rect 2582 69040 2890 69060
rect 2872 68808 2924 68814
rect 2872 68750 2924 68756
rect 2504 68740 2556 68746
rect 2504 68682 2556 68688
rect 2412 67312 2464 67318
rect 2412 67254 2464 67260
rect 2412 67176 2464 67182
rect 2412 67118 2464 67124
rect 2280 64416 2360 64444
rect 2228 64398 2280 64404
rect 2226 64152 2282 64161
rect 2226 64087 2282 64096
rect 2240 61742 2268 64087
rect 2320 62688 2372 62694
rect 2318 62656 2320 62665
rect 2372 62656 2374 62665
rect 2318 62591 2374 62600
rect 2424 62370 2452 67118
rect 2516 66722 2544 68682
rect 2884 68490 2912 68750
rect 2976 68649 3004 69362
rect 3068 68814 3096 69430
rect 3056 68808 3108 68814
rect 3056 68750 3108 68756
rect 3160 68746 3188 73510
rect 3148 68740 3200 68746
rect 3148 68682 3200 68688
rect 2962 68640 3018 68649
rect 2962 68575 3018 68584
rect 2884 68462 3004 68490
rect 2582 68028 2890 68048
rect 2582 68026 2588 68028
rect 2644 68026 2668 68028
rect 2724 68026 2748 68028
rect 2804 68026 2828 68028
rect 2884 68026 2890 68028
rect 2644 67974 2646 68026
rect 2826 67974 2828 68026
rect 2582 67972 2588 67974
rect 2644 67972 2668 67974
rect 2724 67972 2748 67974
rect 2804 67972 2828 67974
rect 2884 67972 2890 67974
rect 2582 67952 2890 67972
rect 2582 66940 2890 66960
rect 2582 66938 2588 66940
rect 2644 66938 2668 66940
rect 2724 66938 2748 66940
rect 2804 66938 2828 66940
rect 2884 66938 2890 66940
rect 2644 66886 2646 66938
rect 2826 66886 2828 66938
rect 2582 66884 2588 66886
rect 2644 66884 2668 66886
rect 2724 66884 2748 66886
rect 2804 66884 2828 66886
rect 2884 66884 2890 66886
rect 2582 66864 2890 66884
rect 2516 66694 2636 66722
rect 2976 66706 3004 68462
rect 3056 67244 3108 67250
rect 3056 67186 3108 67192
rect 2504 66632 2556 66638
rect 2504 66574 2556 66580
rect 2332 62342 2452 62370
rect 2228 61736 2280 61742
rect 2228 61678 2280 61684
rect 2136 61600 2188 61606
rect 2136 61542 2188 61548
rect 2228 61328 2280 61334
rect 2228 61270 2280 61276
rect 2240 60246 2268 61270
rect 2332 60761 2360 62342
rect 2412 62280 2464 62286
rect 2412 62222 2464 62228
rect 2424 61810 2452 62222
rect 2412 61804 2464 61810
rect 2412 61746 2464 61752
rect 2412 61600 2464 61606
rect 2412 61542 2464 61548
rect 2318 60752 2374 60761
rect 2318 60687 2374 60696
rect 2320 60512 2372 60518
rect 2320 60454 2372 60460
rect 2228 60240 2280 60246
rect 2228 60182 2280 60188
rect 2332 60081 2360 60454
rect 2318 60072 2374 60081
rect 2318 60007 2374 60016
rect 2044 59968 2096 59974
rect 2044 59910 2096 59916
rect 2318 59936 2374 59945
rect 2424 59922 2452 61542
rect 2516 61282 2544 66574
rect 2608 66502 2636 66694
rect 2964 66700 3016 66706
rect 2964 66642 3016 66648
rect 2596 66496 2648 66502
rect 2596 66438 2648 66444
rect 2964 66496 3016 66502
rect 3068 66473 3096 67186
rect 3148 66700 3200 66706
rect 3148 66642 3200 66648
rect 2964 66438 3016 66444
rect 3054 66464 3110 66473
rect 2582 65852 2890 65872
rect 2582 65850 2588 65852
rect 2644 65850 2668 65852
rect 2724 65850 2748 65852
rect 2804 65850 2828 65852
rect 2884 65850 2890 65852
rect 2644 65798 2646 65850
rect 2826 65798 2828 65850
rect 2582 65796 2588 65798
rect 2644 65796 2668 65798
rect 2724 65796 2748 65798
rect 2804 65796 2828 65798
rect 2884 65796 2890 65798
rect 2582 65776 2890 65796
rect 2976 65657 3004 66438
rect 3054 66399 3110 66408
rect 3160 66230 3188 66642
rect 3148 66224 3200 66230
rect 3148 66166 3200 66172
rect 3056 65952 3108 65958
rect 3056 65894 3108 65900
rect 2962 65648 3018 65657
rect 2962 65583 3018 65592
rect 2964 65544 3016 65550
rect 2964 65486 3016 65492
rect 2780 65476 2832 65482
rect 2780 65418 2832 65424
rect 2792 65006 2820 65418
rect 2976 65074 3004 65486
rect 2964 65068 3016 65074
rect 2964 65010 3016 65016
rect 2780 65000 2832 65006
rect 2780 64942 2832 64948
rect 2582 64764 2890 64784
rect 2582 64762 2588 64764
rect 2644 64762 2668 64764
rect 2724 64762 2748 64764
rect 2804 64762 2828 64764
rect 2884 64762 2890 64764
rect 2644 64710 2646 64762
rect 2826 64710 2828 64762
rect 2582 64708 2588 64710
rect 2644 64708 2668 64710
rect 2724 64708 2748 64710
rect 2804 64708 2828 64710
rect 2884 64708 2890 64710
rect 2582 64688 2890 64708
rect 2976 64462 3004 65010
rect 3068 64569 3096 65894
rect 3160 65074 3188 66166
rect 3252 65142 3280 76214
rect 3516 75744 3568 75750
rect 3516 75686 3568 75692
rect 3332 73228 3384 73234
rect 3332 73170 3384 73176
rect 3240 65136 3292 65142
rect 3240 65078 3292 65084
rect 3148 65068 3200 65074
rect 3148 65010 3200 65016
rect 3148 64932 3200 64938
rect 3148 64874 3200 64880
rect 3054 64560 3110 64569
rect 3054 64495 3110 64504
rect 2964 64456 3016 64462
rect 2964 64398 3016 64404
rect 2976 63918 3004 64398
rect 3056 64320 3108 64326
rect 3054 64288 3056 64297
rect 3108 64288 3110 64297
rect 3054 64223 3110 64232
rect 2964 63912 3016 63918
rect 2964 63854 3016 63860
rect 3054 63880 3110 63889
rect 2582 63676 2890 63696
rect 2582 63674 2588 63676
rect 2644 63674 2668 63676
rect 2724 63674 2748 63676
rect 2804 63674 2828 63676
rect 2884 63674 2890 63676
rect 2644 63622 2646 63674
rect 2826 63622 2828 63674
rect 2582 63620 2588 63622
rect 2644 63620 2668 63622
rect 2724 63620 2748 63622
rect 2804 63620 2828 63622
rect 2884 63620 2890 63622
rect 2582 63600 2890 63620
rect 2872 63368 2924 63374
rect 2872 63310 2924 63316
rect 2884 62937 2912 63310
rect 2870 62928 2926 62937
rect 2870 62863 2926 62872
rect 2582 62588 2890 62608
rect 2582 62586 2588 62588
rect 2644 62586 2668 62588
rect 2724 62586 2748 62588
rect 2804 62586 2828 62588
rect 2884 62586 2890 62588
rect 2644 62534 2646 62586
rect 2826 62534 2828 62586
rect 2582 62532 2588 62534
rect 2644 62532 2668 62534
rect 2724 62532 2748 62534
rect 2804 62532 2828 62534
rect 2884 62532 2890 62534
rect 2582 62512 2890 62532
rect 2976 62286 3004 63854
rect 3054 63815 3110 63824
rect 3068 63510 3096 63815
rect 3056 63504 3108 63510
rect 3056 63446 3108 63452
rect 3056 62892 3108 62898
rect 3056 62834 3108 62840
rect 2964 62280 3016 62286
rect 2964 62222 3016 62228
rect 2596 62212 2648 62218
rect 2596 62154 2648 62160
rect 2608 61674 2636 62154
rect 2964 62144 3016 62150
rect 2964 62086 3016 62092
rect 2686 61840 2742 61849
rect 2686 61775 2688 61784
rect 2740 61775 2742 61784
rect 2688 61746 2740 61752
rect 2596 61668 2648 61674
rect 2596 61610 2648 61616
rect 2582 61500 2890 61520
rect 2582 61498 2588 61500
rect 2644 61498 2668 61500
rect 2724 61498 2748 61500
rect 2804 61498 2828 61500
rect 2884 61498 2890 61500
rect 2644 61446 2646 61498
rect 2826 61446 2828 61498
rect 2582 61444 2588 61446
rect 2644 61444 2668 61446
rect 2724 61444 2748 61446
rect 2804 61444 2828 61446
rect 2884 61444 2890 61446
rect 2582 61424 2890 61444
rect 2516 61254 2728 61282
rect 2502 61024 2558 61033
rect 2502 60959 2558 60968
rect 2516 60042 2544 60959
rect 2700 60858 2728 61254
rect 2780 61056 2832 61062
rect 2780 60998 2832 61004
rect 2792 60897 2820 60998
rect 2778 60888 2834 60897
rect 2688 60852 2740 60858
rect 2778 60823 2834 60832
rect 2688 60794 2740 60800
rect 2976 60761 3004 62086
rect 2962 60752 3018 60761
rect 2962 60687 3018 60696
rect 2962 60616 3018 60625
rect 2962 60551 2964 60560
rect 3016 60551 3018 60560
rect 2964 60522 3016 60528
rect 3068 60466 3096 62834
rect 2976 60438 3096 60466
rect 2582 60412 2890 60432
rect 2582 60410 2588 60412
rect 2644 60410 2668 60412
rect 2724 60410 2748 60412
rect 2804 60410 2828 60412
rect 2884 60410 2890 60412
rect 2644 60358 2646 60410
rect 2826 60358 2828 60410
rect 2582 60356 2588 60358
rect 2644 60356 2668 60358
rect 2724 60356 2748 60358
rect 2804 60356 2828 60358
rect 2884 60356 2890 60358
rect 2582 60336 2890 60356
rect 2688 60240 2740 60246
rect 2688 60182 2740 60188
rect 2596 60172 2648 60178
rect 2596 60114 2648 60120
rect 2504 60036 2556 60042
rect 2504 59978 2556 59984
rect 2424 59894 2544 59922
rect 2318 59871 2374 59880
rect 2044 59764 2096 59770
rect 2332 59752 2360 59871
rect 2044 59706 2096 59712
rect 2148 59724 2360 59752
rect 2056 59226 2084 59706
rect 2148 59634 2176 59724
rect 2136 59628 2188 59634
rect 2136 59570 2188 59576
rect 2134 59528 2190 59537
rect 2134 59463 2190 59472
rect 2320 59492 2372 59498
rect 2148 59430 2176 59463
rect 2320 59434 2372 59440
rect 2412 59492 2464 59498
rect 2412 59434 2464 59440
rect 2136 59424 2188 59430
rect 2136 59366 2188 59372
rect 2228 59424 2280 59430
rect 2228 59366 2280 59372
rect 1952 59220 2004 59226
rect 1952 59162 2004 59168
rect 2044 59220 2096 59226
rect 2044 59162 2096 59168
rect 2148 58886 2176 59366
rect 2044 58880 2096 58886
rect 2044 58822 2096 58828
rect 2136 58880 2188 58886
rect 2240 58857 2268 59366
rect 2332 59226 2360 59434
rect 2320 59220 2372 59226
rect 2320 59162 2372 59168
rect 2136 58822 2188 58828
rect 2226 58848 2282 58857
rect 1952 58540 2004 58546
rect 1952 58482 2004 58488
rect 1964 57497 1992 58482
rect 1950 57488 2006 57497
rect 1950 57423 2006 57432
rect 1952 56976 2004 56982
rect 1952 56918 2004 56924
rect 1964 46714 1992 56918
rect 2056 54126 2084 58822
rect 2148 57458 2176 58822
rect 2226 58783 2282 58792
rect 2332 58614 2360 59162
rect 2228 58608 2280 58614
rect 2228 58550 2280 58556
rect 2320 58608 2372 58614
rect 2320 58550 2372 58556
rect 2136 57452 2188 57458
rect 2136 57394 2188 57400
rect 2136 57248 2188 57254
rect 2136 57190 2188 57196
rect 2044 54120 2096 54126
rect 2044 54062 2096 54068
rect 2044 53984 2096 53990
rect 2044 53926 2096 53932
rect 2056 53689 2084 53926
rect 2042 53680 2098 53689
rect 2042 53615 2098 53624
rect 2044 53236 2096 53242
rect 2044 53178 2096 53184
rect 1952 46708 2004 46714
rect 1952 46650 2004 46656
rect 1872 46158 1992 46186
rect 1860 45416 1912 45422
rect 1860 45358 1912 45364
rect 1872 45082 1900 45358
rect 1860 45076 1912 45082
rect 1860 45018 1912 45024
rect 1860 44736 1912 44742
rect 1860 44678 1912 44684
rect 1766 42392 1822 42401
rect 1766 42327 1822 42336
rect 1768 42288 1820 42294
rect 1768 42230 1820 42236
rect 1780 41732 1808 42230
rect 1872 41857 1900 44678
rect 1964 42945 1992 46158
rect 1950 42936 2006 42945
rect 1950 42871 2006 42880
rect 1950 42800 2006 42809
rect 1950 42735 2006 42744
rect 1858 41848 1914 41857
rect 1858 41783 1914 41792
rect 1780 41704 1900 41732
rect 1768 41472 1820 41478
rect 1674 41440 1730 41449
rect 1768 41414 1820 41420
rect 1674 41375 1730 41384
rect 1676 41200 1728 41206
rect 1676 41142 1728 41148
rect 1688 38978 1716 41142
rect 1780 39098 1808 41414
rect 1768 39092 1820 39098
rect 1768 39034 1820 39040
rect 1688 38950 1808 38978
rect 1676 38888 1728 38894
rect 1676 38830 1728 38836
rect 1582 38584 1638 38593
rect 1306 38519 1362 38528
rect 1400 38548 1452 38554
rect 1400 38490 1452 38496
rect 1492 38548 1544 38554
rect 1688 38554 1716 38830
rect 1780 38554 1808 38950
rect 1582 38519 1638 38528
rect 1676 38548 1728 38554
rect 1492 38490 1544 38496
rect 1676 38490 1728 38496
rect 1768 38548 1820 38554
rect 1768 38490 1820 38496
rect 1582 38448 1638 38457
rect 1308 38412 1360 38418
rect 1360 38372 1532 38400
rect 1582 38383 1638 38392
rect 1676 38412 1728 38418
rect 1308 38354 1360 38360
rect 1124 38344 1176 38350
rect 1504 38321 1532 38372
rect 1124 38286 1176 38292
rect 1306 38312 1362 38321
rect 1306 38247 1362 38256
rect 1490 38312 1546 38321
rect 1490 38247 1546 38256
rect 1124 38004 1176 38010
rect 1124 37946 1176 37952
rect 1136 36922 1164 37946
rect 1216 37936 1268 37942
rect 1216 37878 1268 37884
rect 1124 36916 1176 36922
rect 1124 36858 1176 36864
rect 1124 36712 1176 36718
rect 1124 36654 1176 36660
rect 1136 31822 1164 36654
rect 1124 31816 1176 31822
rect 1124 31758 1176 31764
rect 1124 31680 1176 31686
rect 1124 31622 1176 31628
rect 1136 31385 1164 31622
rect 1122 31376 1178 31385
rect 1122 31311 1178 31320
rect 1124 30320 1176 30326
rect 1122 30288 1124 30297
rect 1176 30288 1178 30297
rect 1122 30223 1178 30232
rect 1228 28200 1256 37878
rect 1136 28172 1256 28200
rect 1032 27464 1084 27470
rect 1032 27406 1084 27412
rect 1136 24614 1164 28172
rect 1214 27976 1270 27985
rect 1214 27911 1270 27920
rect 1228 27538 1256 27911
rect 1216 27532 1268 27538
rect 1216 27474 1268 27480
rect 1124 24608 1176 24614
rect 1124 24550 1176 24556
rect 1216 23656 1268 23662
rect 1216 23598 1268 23604
rect 1228 22817 1256 23598
rect 1214 22808 1270 22817
rect 1214 22743 1270 22752
rect 1216 22568 1268 22574
rect 1216 22510 1268 22516
rect 940 22296 992 22302
rect 940 22238 992 22244
rect 940 22160 992 22166
rect 940 22102 992 22108
rect 952 21622 980 22102
rect 1228 22001 1256 22510
rect 1214 21992 1270 22001
rect 1214 21927 1270 21936
rect 940 21616 992 21622
rect 940 21558 992 21564
rect 1032 18352 1084 18358
rect 1032 18294 1084 18300
rect 1044 11762 1072 18294
rect 1320 17252 1348 38247
rect 1400 37800 1452 37806
rect 1400 37742 1452 37748
rect 1412 35018 1440 37742
rect 1492 37460 1544 37466
rect 1492 37402 1544 37408
rect 1504 37262 1532 37402
rect 1492 37256 1544 37262
rect 1492 37198 1544 37204
rect 1596 37210 1624 38383
rect 1676 38354 1728 38360
rect 1688 38010 1716 38354
rect 1768 38344 1820 38350
rect 1768 38286 1820 38292
rect 1676 38004 1728 38010
rect 1676 37946 1728 37952
rect 1676 37732 1728 37738
rect 1676 37674 1728 37680
rect 1688 37330 1716 37674
rect 1676 37324 1728 37330
rect 1676 37266 1728 37272
rect 1596 37182 1716 37210
rect 1584 37120 1636 37126
rect 1584 37062 1636 37068
rect 1492 36168 1544 36174
rect 1596 36145 1624 37062
rect 1492 36110 1544 36116
rect 1582 36136 1638 36145
rect 1504 35290 1532 36110
rect 1582 36071 1638 36080
rect 1584 35488 1636 35494
rect 1584 35430 1636 35436
rect 1492 35284 1544 35290
rect 1492 35226 1544 35232
rect 1596 35193 1624 35430
rect 1582 35184 1638 35193
rect 1582 35119 1638 35128
rect 1492 35080 1544 35086
rect 1492 35022 1544 35028
rect 1400 35012 1452 35018
rect 1400 34954 1452 34960
rect 1400 34400 1452 34406
rect 1400 34342 1452 34348
rect 1412 33561 1440 34342
rect 1398 33552 1454 33561
rect 1398 33487 1454 33496
rect 1504 33402 1532 35022
rect 1582 34776 1638 34785
rect 1582 34711 1584 34720
rect 1636 34711 1638 34720
rect 1584 34682 1636 34688
rect 1412 33374 1532 33402
rect 1412 31929 1440 33374
rect 1490 33280 1546 33289
rect 1490 33215 1546 33224
rect 1504 32978 1532 33215
rect 1492 32972 1544 32978
rect 1492 32914 1544 32920
rect 1688 32910 1716 37182
rect 1676 32904 1728 32910
rect 1490 32872 1546 32881
rect 1676 32846 1728 32852
rect 1490 32807 1546 32816
rect 1398 31920 1454 31929
rect 1398 31855 1454 31864
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 28218 1440 31758
rect 1504 31634 1532 32807
rect 1584 32564 1636 32570
rect 1584 32506 1636 32512
rect 1596 31754 1624 32506
rect 1674 32192 1730 32201
rect 1674 32127 1730 32136
rect 1584 31748 1636 31754
rect 1584 31690 1636 31696
rect 1504 31606 1624 31634
rect 1490 31512 1546 31521
rect 1490 31447 1546 31456
rect 1400 28212 1452 28218
rect 1400 28154 1452 28160
rect 1400 28008 1452 28014
rect 1400 27950 1452 27956
rect 1412 27577 1440 27950
rect 1398 27568 1454 27577
rect 1398 27503 1454 27512
rect 1400 25832 1452 25838
rect 1400 25774 1452 25780
rect 1412 25401 1440 25774
rect 1398 25392 1454 25401
rect 1398 25327 1454 25336
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1412 24993 1440 25230
rect 1398 24984 1454 24993
rect 1398 24919 1454 24928
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 23225 1440 24142
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 22409 1440 23054
rect 1398 22400 1454 22409
rect 1398 22335 1454 22344
rect 1504 22098 1532 31447
rect 1492 22092 1544 22098
rect 1492 22034 1544 22040
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1412 21593 1440 21966
rect 1398 21584 1454 21593
rect 1398 21519 1454 21528
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 21185 1440 21422
rect 1398 21176 1454 21185
rect 1398 21111 1454 21120
rect 1596 21026 1624 31606
rect 1688 30410 1716 32127
rect 1780 30734 1808 38286
rect 1872 38282 1900 41704
rect 1964 41546 1992 42735
rect 1952 41540 2004 41546
rect 1952 41482 2004 41488
rect 1952 41132 2004 41138
rect 1952 41074 2004 41080
rect 1964 40118 1992 41074
rect 1952 40112 2004 40118
rect 1952 40054 2004 40060
rect 1952 39092 2004 39098
rect 1952 39034 2004 39040
rect 1964 38554 1992 39034
rect 2056 38554 2084 53178
rect 2148 52902 2176 57190
rect 2240 53242 2268 58550
rect 2332 57390 2360 58550
rect 2424 57633 2452 59434
rect 2410 57624 2466 57633
rect 2410 57559 2466 57568
rect 2320 57384 2372 57390
rect 2372 57344 2452 57372
rect 2320 57326 2372 57332
rect 2320 56840 2372 56846
rect 2320 56782 2372 56788
rect 2332 56250 2360 56782
rect 2424 56778 2452 57344
rect 2412 56772 2464 56778
rect 2412 56714 2464 56720
rect 2332 56222 2452 56250
rect 2320 56160 2372 56166
rect 2320 56102 2372 56108
rect 2332 55729 2360 56102
rect 2318 55720 2374 55729
rect 2318 55655 2374 55664
rect 2320 55616 2372 55622
rect 2320 55558 2372 55564
rect 2332 55321 2360 55558
rect 2318 55312 2374 55321
rect 2318 55247 2374 55256
rect 2424 54890 2452 56222
rect 2332 54862 2452 54890
rect 2332 54670 2360 54862
rect 2412 54800 2464 54806
rect 2412 54742 2464 54748
rect 2320 54664 2372 54670
rect 2320 54606 2372 54612
rect 2332 54126 2360 54606
rect 2320 54120 2372 54126
rect 2320 54062 2372 54068
rect 2332 53650 2360 54062
rect 2320 53644 2372 53650
rect 2320 53586 2372 53592
rect 2320 53440 2372 53446
rect 2320 53382 2372 53388
rect 2228 53236 2280 53242
rect 2228 53178 2280 53184
rect 2332 53145 2360 53382
rect 2318 53136 2374 53145
rect 2228 53100 2280 53106
rect 2318 53071 2374 53080
rect 2228 53042 2280 53048
rect 2136 52896 2188 52902
rect 2136 52838 2188 52844
rect 2134 52728 2190 52737
rect 2134 52663 2190 52672
rect 2148 51241 2176 52663
rect 2134 51232 2190 51241
rect 2134 51167 2190 51176
rect 2136 51060 2188 51066
rect 2136 51002 2188 51008
rect 2148 50930 2176 51002
rect 2136 50924 2188 50930
rect 2136 50866 2188 50872
rect 2134 50824 2190 50833
rect 2134 50759 2190 50768
rect 2148 43858 2176 50759
rect 2240 43926 2268 53042
rect 2320 52488 2372 52494
rect 2320 52430 2372 52436
rect 2332 51610 2360 52430
rect 2320 51604 2372 51610
rect 2320 51546 2372 51552
rect 2424 51456 2452 54742
rect 2516 53106 2544 59894
rect 2608 59770 2636 60114
rect 2596 59764 2648 59770
rect 2596 59706 2648 59712
rect 2596 59628 2648 59634
rect 2596 59570 2648 59576
rect 2608 59537 2636 59570
rect 2700 59566 2728 60182
rect 2780 59968 2832 59974
rect 2780 59910 2832 59916
rect 2792 59673 2820 59910
rect 2778 59664 2834 59673
rect 2778 59599 2834 59608
rect 2688 59560 2740 59566
rect 2594 59528 2650 59537
rect 2688 59502 2740 59508
rect 2594 59463 2650 59472
rect 2582 59324 2890 59344
rect 2582 59322 2588 59324
rect 2644 59322 2668 59324
rect 2724 59322 2748 59324
rect 2804 59322 2828 59324
rect 2884 59322 2890 59324
rect 2644 59270 2646 59322
rect 2826 59270 2828 59322
rect 2582 59268 2588 59270
rect 2644 59268 2668 59270
rect 2724 59268 2748 59270
rect 2804 59268 2828 59270
rect 2884 59268 2890 59270
rect 2582 59248 2890 59268
rect 2596 58948 2648 58954
rect 2596 58890 2648 58896
rect 2608 58614 2636 58890
rect 2596 58608 2648 58614
rect 2596 58550 2648 58556
rect 2686 58576 2742 58585
rect 2686 58511 2688 58520
rect 2740 58511 2742 58520
rect 2688 58482 2740 58488
rect 2582 58236 2890 58256
rect 2582 58234 2588 58236
rect 2644 58234 2668 58236
rect 2724 58234 2748 58236
rect 2804 58234 2828 58236
rect 2884 58234 2890 58236
rect 2644 58182 2646 58234
rect 2826 58182 2828 58234
rect 2582 58180 2588 58182
rect 2644 58180 2668 58182
rect 2724 58180 2748 58182
rect 2804 58180 2828 58182
rect 2884 58180 2890 58182
rect 2582 58160 2890 58180
rect 2780 58064 2832 58070
rect 2700 58012 2780 58018
rect 2700 58006 2832 58012
rect 2700 57990 2820 58006
rect 2594 57896 2650 57905
rect 2594 57831 2650 57840
rect 2608 57798 2636 57831
rect 2596 57792 2648 57798
rect 2596 57734 2648 57740
rect 2700 57361 2728 57990
rect 2686 57352 2742 57361
rect 2686 57287 2742 57296
rect 2582 57148 2890 57168
rect 2582 57146 2588 57148
rect 2644 57146 2668 57148
rect 2724 57146 2748 57148
rect 2804 57146 2828 57148
rect 2884 57146 2890 57148
rect 2644 57094 2646 57146
rect 2826 57094 2828 57146
rect 2582 57092 2588 57094
rect 2644 57092 2668 57094
rect 2724 57092 2748 57094
rect 2804 57092 2828 57094
rect 2884 57092 2890 57094
rect 2582 57072 2890 57092
rect 2686 56264 2742 56273
rect 2686 56199 2688 56208
rect 2740 56199 2742 56208
rect 2688 56170 2740 56176
rect 2582 56060 2890 56080
rect 2582 56058 2588 56060
rect 2644 56058 2668 56060
rect 2724 56058 2748 56060
rect 2804 56058 2828 56060
rect 2884 56058 2890 56060
rect 2644 56006 2646 56058
rect 2826 56006 2828 56058
rect 2582 56004 2588 56006
rect 2644 56004 2668 56006
rect 2724 56004 2748 56006
rect 2804 56004 2828 56006
rect 2884 56004 2890 56006
rect 2582 55984 2890 56004
rect 2872 55752 2924 55758
rect 2870 55720 2872 55729
rect 2924 55720 2926 55729
rect 2870 55655 2926 55664
rect 2976 55298 3004 60438
rect 3054 60344 3110 60353
rect 3054 60279 3110 60288
rect 3068 57390 3096 60279
rect 3056 57384 3108 57390
rect 3056 57326 3108 57332
rect 3056 56840 3108 56846
rect 3056 56782 3108 56788
rect 3068 55418 3096 56782
rect 3056 55412 3108 55418
rect 3056 55354 3108 55360
rect 2884 55270 3004 55298
rect 3054 55312 3110 55321
rect 2884 55060 2912 55270
rect 3160 55298 3188 64874
rect 3240 64864 3292 64870
rect 3240 64806 3292 64812
rect 3252 63986 3280 64806
rect 3240 63980 3292 63986
rect 3240 63922 3292 63928
rect 3252 63481 3280 63922
rect 3238 63472 3294 63481
rect 3238 63407 3294 63416
rect 3240 63300 3292 63306
rect 3240 63242 3292 63248
rect 3252 60897 3280 63242
rect 3238 60888 3294 60897
rect 3238 60823 3294 60832
rect 3238 60752 3294 60761
rect 3238 60687 3240 60696
rect 3292 60687 3294 60696
rect 3240 60658 3292 60664
rect 3240 59424 3292 59430
rect 3240 59366 3292 59372
rect 3252 58070 3280 59366
rect 3240 58064 3292 58070
rect 3240 58006 3292 58012
rect 3240 57384 3292 57390
rect 3240 57326 3292 57332
rect 3252 55826 3280 57326
rect 3240 55820 3292 55826
rect 3240 55762 3292 55768
rect 3240 55616 3292 55622
rect 3240 55558 3292 55564
rect 3252 55418 3280 55558
rect 3240 55412 3292 55418
rect 3240 55354 3292 55360
rect 3160 55270 3280 55298
rect 3054 55247 3110 55256
rect 2884 55032 3004 55060
rect 2582 54972 2890 54992
rect 2582 54970 2588 54972
rect 2644 54970 2668 54972
rect 2724 54970 2748 54972
rect 2804 54970 2828 54972
rect 2884 54970 2890 54972
rect 2644 54918 2646 54970
rect 2826 54918 2828 54970
rect 2582 54916 2588 54918
rect 2644 54916 2668 54918
rect 2724 54916 2748 54918
rect 2804 54916 2828 54918
rect 2884 54916 2890 54918
rect 2582 54896 2890 54916
rect 2780 54528 2832 54534
rect 2778 54496 2780 54505
rect 2832 54496 2834 54505
rect 2778 54431 2834 54440
rect 2582 53884 2890 53904
rect 2582 53882 2588 53884
rect 2644 53882 2668 53884
rect 2724 53882 2748 53884
rect 2804 53882 2828 53884
rect 2884 53882 2890 53884
rect 2644 53830 2646 53882
rect 2826 53830 2828 53882
rect 2582 53828 2588 53830
rect 2644 53828 2668 53830
rect 2724 53828 2748 53830
rect 2804 53828 2828 53830
rect 2884 53828 2890 53830
rect 2582 53808 2890 53828
rect 2596 53644 2648 53650
rect 2596 53586 2648 53592
rect 2504 53100 2556 53106
rect 2504 53042 2556 53048
rect 2608 53009 2636 53586
rect 2594 53000 2650 53009
rect 2594 52935 2650 52944
rect 2504 52896 2556 52902
rect 2504 52838 2556 52844
rect 2332 51428 2452 51456
rect 2332 51066 2360 51428
rect 2320 51060 2372 51066
rect 2320 51002 2372 51008
rect 2516 50946 2544 52838
rect 2582 52796 2890 52816
rect 2582 52794 2588 52796
rect 2644 52794 2668 52796
rect 2724 52794 2748 52796
rect 2804 52794 2828 52796
rect 2884 52794 2890 52796
rect 2644 52742 2646 52794
rect 2826 52742 2828 52794
rect 2582 52740 2588 52742
rect 2644 52740 2668 52742
rect 2724 52740 2748 52742
rect 2804 52740 2828 52742
rect 2884 52740 2890 52742
rect 2582 52720 2890 52740
rect 2872 52148 2924 52154
rect 2872 52090 2924 52096
rect 2884 51921 2912 52090
rect 2870 51912 2926 51921
rect 2870 51847 2926 51856
rect 2582 51708 2890 51728
rect 2582 51706 2588 51708
rect 2644 51706 2668 51708
rect 2724 51706 2748 51708
rect 2804 51706 2828 51708
rect 2884 51706 2890 51708
rect 2644 51654 2646 51706
rect 2826 51654 2828 51706
rect 2582 51652 2588 51654
rect 2644 51652 2668 51654
rect 2724 51652 2748 51654
rect 2804 51652 2828 51654
rect 2884 51652 2890 51654
rect 2582 51632 2890 51652
rect 2976 51610 3004 55032
rect 2964 51604 3016 51610
rect 2964 51546 3016 51552
rect 2596 51400 2648 51406
rect 2596 51342 2648 51348
rect 2332 50918 2544 50946
rect 2332 49178 2360 50918
rect 2608 50862 2636 51342
rect 2780 51332 2832 51338
rect 2780 51274 2832 51280
rect 2792 50862 2820 51274
rect 2596 50856 2648 50862
rect 2516 50816 2596 50844
rect 2516 50504 2544 50816
rect 2596 50798 2648 50804
rect 2780 50856 2832 50862
rect 2780 50798 2832 50804
rect 2964 50720 3016 50726
rect 2964 50662 3016 50668
rect 2582 50620 2890 50640
rect 2582 50618 2588 50620
rect 2644 50618 2668 50620
rect 2724 50618 2748 50620
rect 2804 50618 2828 50620
rect 2884 50618 2890 50620
rect 2644 50566 2646 50618
rect 2826 50566 2828 50618
rect 2582 50564 2588 50566
rect 2644 50564 2668 50566
rect 2724 50564 2748 50566
rect 2804 50564 2828 50566
rect 2884 50564 2890 50566
rect 2582 50544 2890 50564
rect 2516 50476 2636 50504
rect 2504 49836 2556 49842
rect 2504 49778 2556 49784
rect 2516 49722 2544 49778
rect 2608 49774 2636 50476
rect 2872 50448 2924 50454
rect 2872 50390 2924 50396
rect 2780 50176 2832 50182
rect 2780 50118 2832 50124
rect 2424 49694 2544 49722
rect 2596 49768 2648 49774
rect 2792 49745 2820 50118
rect 2884 49994 2912 50390
rect 2976 50153 3004 50662
rect 2962 50144 3018 50153
rect 2962 50079 3018 50088
rect 2884 49966 3004 49994
rect 2596 49710 2648 49716
rect 2778 49736 2834 49745
rect 2424 49434 2452 49694
rect 2778 49671 2834 49680
rect 2504 49632 2556 49638
rect 2504 49574 2556 49580
rect 2412 49428 2464 49434
rect 2412 49370 2464 49376
rect 2516 49337 2544 49574
rect 2582 49532 2890 49552
rect 2582 49530 2588 49532
rect 2644 49530 2668 49532
rect 2724 49530 2748 49532
rect 2804 49530 2828 49532
rect 2884 49530 2890 49532
rect 2644 49478 2646 49530
rect 2826 49478 2828 49530
rect 2582 49476 2588 49478
rect 2644 49476 2668 49478
rect 2724 49476 2748 49478
rect 2804 49476 2828 49478
rect 2884 49476 2890 49478
rect 2582 49456 2890 49476
rect 2688 49360 2740 49366
rect 2502 49328 2558 49337
rect 2688 49302 2740 49308
rect 2778 49328 2834 49337
rect 2502 49263 2558 49272
rect 2594 49192 2650 49201
rect 2332 49150 2452 49178
rect 2320 49088 2372 49094
rect 2320 49030 2372 49036
rect 2332 48929 2360 49030
rect 2318 48920 2374 48929
rect 2318 48855 2374 48864
rect 2424 48804 2452 49150
rect 2594 49127 2650 49136
rect 2502 49056 2558 49065
rect 2502 48991 2558 49000
rect 2332 48776 2452 48804
rect 2228 43920 2280 43926
rect 2228 43862 2280 43868
rect 2136 43852 2188 43858
rect 2136 43794 2188 43800
rect 2332 43772 2360 48776
rect 2516 48736 2544 48991
rect 2424 48708 2544 48736
rect 2424 48249 2452 48708
rect 2608 48668 2636 49127
rect 2700 48822 2728 49302
rect 2778 49263 2834 49272
rect 2872 49292 2924 49298
rect 2688 48816 2740 48822
rect 2688 48758 2740 48764
rect 2792 48754 2820 49263
rect 2872 49234 2924 49240
rect 2884 49201 2912 49234
rect 2870 49192 2926 49201
rect 2870 49127 2926 49136
rect 2976 48822 3004 49966
rect 2964 48816 3016 48822
rect 2964 48758 3016 48764
rect 2780 48748 2832 48754
rect 2780 48690 2832 48696
rect 2516 48640 2636 48668
rect 2964 48680 3016 48686
rect 2962 48648 2964 48657
rect 3016 48648 3018 48657
rect 2410 48240 2466 48249
rect 2410 48175 2466 48184
rect 2412 48136 2464 48142
rect 2412 48078 2464 48084
rect 2424 47977 2452 48078
rect 2410 47968 2466 47977
rect 2410 47903 2466 47912
rect 2412 47592 2464 47598
rect 2412 47534 2464 47540
rect 2424 47258 2452 47534
rect 2412 47252 2464 47258
rect 2412 47194 2464 47200
rect 2412 47116 2464 47122
rect 2412 47058 2464 47064
rect 2424 46578 2452 47058
rect 2412 46572 2464 46578
rect 2412 46514 2464 46520
rect 2424 44878 2452 46514
rect 2412 44872 2464 44878
rect 2412 44814 2464 44820
rect 2516 44248 2544 48640
rect 2962 48583 3018 48592
rect 2582 48444 2890 48464
rect 2582 48442 2588 48444
rect 2644 48442 2668 48444
rect 2724 48442 2748 48444
rect 2804 48442 2828 48444
rect 2884 48442 2890 48444
rect 2644 48390 2646 48442
rect 2826 48390 2828 48442
rect 2582 48388 2588 48390
rect 2644 48388 2668 48390
rect 2724 48388 2748 48390
rect 2804 48388 2828 48390
rect 2884 48388 2890 48390
rect 2582 48368 2890 48388
rect 2688 48326 2740 48332
rect 2688 48268 2740 48274
rect 2780 48272 2832 48278
rect 2596 48136 2648 48142
rect 2596 48078 2648 48084
rect 2608 47734 2636 48078
rect 2700 47841 2728 48268
rect 2778 48240 2780 48249
rect 2832 48240 2834 48249
rect 2778 48175 2834 48184
rect 2964 48068 3016 48074
rect 2964 48010 3016 48016
rect 2686 47832 2742 47841
rect 2686 47767 2742 47776
rect 2596 47728 2648 47734
rect 2596 47670 2648 47676
rect 2582 47356 2890 47376
rect 2582 47354 2588 47356
rect 2644 47354 2668 47356
rect 2724 47354 2748 47356
rect 2804 47354 2828 47356
rect 2884 47354 2890 47356
rect 2644 47302 2646 47354
rect 2826 47302 2828 47354
rect 2582 47300 2588 47302
rect 2644 47300 2668 47302
rect 2724 47300 2748 47302
rect 2804 47300 2828 47302
rect 2884 47300 2890 47302
rect 2582 47280 2890 47300
rect 2582 46268 2890 46288
rect 2582 46266 2588 46268
rect 2644 46266 2668 46268
rect 2724 46266 2748 46268
rect 2804 46266 2828 46268
rect 2884 46266 2890 46268
rect 2644 46214 2646 46266
rect 2826 46214 2828 46266
rect 2582 46212 2588 46214
rect 2644 46212 2668 46214
rect 2724 46212 2748 46214
rect 2804 46212 2828 46214
rect 2884 46212 2890 46214
rect 2582 46192 2890 46212
rect 2686 46064 2742 46073
rect 2686 45999 2742 46008
rect 2700 45966 2728 45999
rect 2688 45960 2740 45966
rect 2688 45902 2740 45908
rect 2870 45928 2926 45937
rect 2870 45863 2926 45872
rect 2884 45830 2912 45863
rect 2872 45824 2924 45830
rect 2872 45766 2924 45772
rect 2870 45656 2926 45665
rect 2870 45591 2926 45600
rect 2884 45558 2912 45591
rect 2872 45552 2924 45558
rect 2872 45494 2924 45500
rect 2582 45180 2890 45200
rect 2582 45178 2588 45180
rect 2644 45178 2668 45180
rect 2724 45178 2748 45180
rect 2804 45178 2828 45180
rect 2884 45178 2890 45180
rect 2644 45126 2646 45178
rect 2826 45126 2828 45178
rect 2582 45124 2588 45126
rect 2644 45124 2668 45126
rect 2724 45124 2748 45126
rect 2804 45124 2828 45126
rect 2884 45124 2890 45126
rect 2582 45104 2890 45124
rect 2596 44872 2648 44878
rect 2596 44814 2648 44820
rect 2240 43744 2360 43772
rect 2424 44220 2544 44248
rect 2240 43738 2268 43744
rect 2148 43710 2268 43738
rect 2148 38554 2176 43710
rect 2424 43704 2452 44220
rect 2608 44180 2636 44814
rect 2976 44384 3004 48010
rect 3068 46102 3096 55247
rect 3148 55140 3200 55146
rect 3148 55082 3200 55088
rect 3160 51524 3188 55082
rect 3252 51649 3280 55270
rect 3238 51640 3294 51649
rect 3238 51575 3294 51584
rect 3160 51496 3280 51524
rect 3148 51400 3200 51406
rect 3148 51342 3200 51348
rect 3160 51066 3188 51342
rect 3148 51060 3200 51066
rect 3148 51002 3200 51008
rect 3146 50960 3202 50969
rect 3146 50895 3202 50904
rect 3160 49065 3188 50895
rect 3146 49056 3202 49065
rect 3146 48991 3202 49000
rect 3148 48748 3200 48754
rect 3148 48690 3200 48696
rect 3160 47705 3188 48690
rect 3146 47696 3202 47705
rect 3146 47631 3202 47640
rect 3148 47592 3200 47598
rect 3148 47534 3200 47540
rect 3056 46096 3108 46102
rect 3056 46038 3108 46044
rect 3056 45892 3108 45898
rect 3056 45834 3108 45840
rect 3068 44538 3096 45834
rect 3056 44532 3108 44538
rect 3056 44474 3108 44480
rect 2976 44356 3096 44384
rect 2964 44260 3016 44266
rect 2964 44202 3016 44208
rect 2516 44152 2636 44180
rect 2516 43874 2544 44152
rect 2582 44092 2890 44112
rect 2582 44090 2588 44092
rect 2644 44090 2668 44092
rect 2724 44090 2748 44092
rect 2804 44090 2828 44092
rect 2884 44090 2890 44092
rect 2644 44038 2646 44090
rect 2826 44038 2828 44090
rect 2582 44036 2588 44038
rect 2644 44036 2668 44038
rect 2724 44036 2748 44038
rect 2804 44036 2828 44038
rect 2884 44036 2890 44038
rect 2582 44016 2890 44036
rect 2686 43888 2742 43897
rect 2516 43846 2636 43874
rect 2504 43784 2556 43790
rect 2504 43726 2556 43732
rect 2332 43676 2452 43704
rect 2228 43648 2280 43654
rect 2228 43590 2280 43596
rect 2240 42158 2268 43590
rect 2228 42152 2280 42158
rect 2228 42094 2280 42100
rect 2228 42016 2280 42022
rect 2228 41958 2280 41964
rect 2240 41138 2268 41958
rect 2228 41132 2280 41138
rect 2228 41074 2280 41080
rect 2228 40656 2280 40662
rect 2228 40598 2280 40604
rect 2240 40186 2268 40598
rect 2228 40180 2280 40186
rect 2228 40122 2280 40128
rect 2240 39574 2268 40122
rect 2228 39568 2280 39574
rect 2228 39510 2280 39516
rect 2226 38992 2282 39001
rect 2226 38927 2282 38936
rect 2240 38554 2268 38927
rect 1952 38548 2004 38554
rect 1952 38490 2004 38496
rect 2044 38548 2096 38554
rect 2044 38490 2096 38496
rect 2136 38548 2188 38554
rect 2136 38490 2188 38496
rect 2228 38548 2280 38554
rect 2228 38490 2280 38496
rect 1952 38412 2004 38418
rect 2332 38400 2360 43676
rect 2516 43314 2544 43726
rect 2504 43308 2556 43314
rect 2504 43250 2556 43256
rect 2412 43240 2464 43246
rect 2412 43182 2464 43188
rect 2424 42242 2452 43182
rect 2608 43092 2636 43846
rect 2686 43823 2742 43832
rect 2872 43852 2924 43858
rect 2700 43314 2728 43823
rect 2872 43794 2924 43800
rect 2780 43716 2832 43722
rect 2780 43658 2832 43664
rect 2688 43308 2740 43314
rect 2688 43250 2740 43256
rect 2792 43246 2820 43658
rect 2884 43330 2912 43794
rect 2976 43654 3004 44202
rect 2964 43648 3016 43654
rect 2964 43590 3016 43596
rect 3068 43489 3096 44356
rect 3160 43858 3188 47534
rect 3252 46186 3280 51496
rect 3344 48793 3372 73170
rect 3528 72826 3556 75686
rect 3620 74186 3648 76910
rect 3792 76288 3844 76294
rect 3792 76230 3844 76236
rect 3700 75948 3752 75954
rect 3700 75890 3752 75896
rect 3712 75449 3740 75890
rect 3698 75440 3754 75449
rect 3698 75375 3754 75384
rect 3608 74180 3660 74186
rect 3608 74122 3660 74128
rect 3804 73098 3832 76230
rect 3896 74934 3924 77318
rect 4214 77276 4522 77296
rect 4214 77274 4220 77276
rect 4276 77274 4300 77276
rect 4356 77274 4380 77276
rect 4436 77274 4460 77276
rect 4516 77274 4522 77276
rect 4276 77222 4278 77274
rect 4458 77222 4460 77274
rect 4214 77220 4220 77222
rect 4276 77220 4300 77222
rect 4356 77220 4380 77222
rect 4436 77220 4460 77222
rect 4516 77220 4522 77222
rect 4214 77200 4522 77220
rect 7478 77276 7786 77296
rect 7478 77274 7484 77276
rect 7540 77274 7564 77276
rect 7620 77274 7644 77276
rect 7700 77274 7724 77276
rect 7780 77274 7786 77276
rect 7540 77222 7542 77274
rect 7722 77222 7724 77274
rect 7478 77220 7484 77222
rect 7540 77220 7564 77222
rect 7620 77220 7644 77222
rect 7700 77220 7724 77222
rect 7780 77220 7786 77222
rect 7478 77200 7786 77220
rect 5846 76732 6154 76752
rect 5846 76730 5852 76732
rect 5908 76730 5932 76732
rect 5988 76730 6012 76732
rect 6068 76730 6092 76732
rect 6148 76730 6154 76732
rect 5908 76678 5910 76730
rect 6090 76678 6092 76730
rect 5846 76676 5852 76678
rect 5908 76676 5932 76678
rect 5988 76676 6012 76678
rect 6068 76676 6092 76678
rect 6148 76676 6154 76678
rect 5846 76656 6154 76676
rect 3976 76424 4028 76430
rect 3976 76366 4028 76372
rect 3988 76265 4016 76366
rect 3974 76256 4030 76265
rect 3974 76191 4030 76200
rect 4214 76188 4522 76208
rect 4214 76186 4220 76188
rect 4276 76186 4300 76188
rect 4356 76186 4380 76188
rect 4436 76186 4460 76188
rect 4516 76186 4522 76188
rect 4276 76134 4278 76186
rect 4458 76134 4460 76186
rect 4214 76132 4220 76134
rect 4276 76132 4300 76134
rect 4356 76132 4380 76134
rect 4436 76132 4460 76134
rect 4516 76132 4522 76134
rect 4214 76112 4522 76132
rect 7478 76188 7786 76208
rect 7478 76186 7484 76188
rect 7540 76186 7564 76188
rect 7620 76186 7644 76188
rect 7700 76186 7724 76188
rect 7780 76186 7786 76188
rect 7540 76134 7542 76186
rect 7722 76134 7724 76186
rect 7478 76132 7484 76134
rect 7540 76132 7564 76134
rect 7620 76132 7644 76134
rect 7700 76132 7724 76134
rect 7780 76132 7786 76134
rect 7478 76112 7786 76132
rect 5264 76016 5316 76022
rect 5264 75958 5316 75964
rect 4214 75100 4522 75120
rect 4214 75098 4220 75100
rect 4276 75098 4300 75100
rect 4356 75098 4380 75100
rect 4436 75098 4460 75100
rect 4516 75098 4522 75100
rect 4276 75046 4278 75098
rect 4458 75046 4460 75098
rect 4214 75044 4220 75046
rect 4276 75044 4300 75046
rect 4356 75044 4380 75046
rect 4436 75044 4460 75046
rect 4516 75044 4522 75046
rect 4214 75024 4522 75044
rect 3884 74928 3936 74934
rect 3884 74870 3936 74876
rect 4214 74012 4522 74032
rect 4214 74010 4220 74012
rect 4276 74010 4300 74012
rect 4356 74010 4380 74012
rect 4436 74010 4460 74012
rect 4516 74010 4522 74012
rect 4276 73958 4278 74010
rect 4458 73958 4460 74010
rect 4214 73956 4220 73958
rect 4276 73956 4300 73958
rect 4356 73956 4380 73958
rect 4436 73956 4460 73958
rect 4516 73956 4522 73958
rect 4214 73936 4522 73956
rect 3792 73092 3844 73098
rect 3792 73034 3844 73040
rect 4214 72924 4522 72944
rect 4214 72922 4220 72924
rect 4276 72922 4300 72924
rect 4356 72922 4380 72924
rect 4436 72922 4460 72924
rect 4516 72922 4522 72924
rect 4276 72870 4278 72922
rect 4458 72870 4460 72922
rect 4214 72868 4220 72870
rect 4276 72868 4300 72870
rect 4356 72868 4380 72870
rect 4436 72868 4460 72870
rect 4516 72868 4522 72870
rect 4214 72848 4522 72868
rect 3516 72820 3568 72826
rect 3516 72762 3568 72768
rect 3884 72480 3936 72486
rect 3884 72422 3936 72428
rect 4620 72480 4672 72486
rect 4620 72422 4672 72428
rect 3700 71596 3752 71602
rect 3700 71538 3752 71544
rect 3516 70644 3568 70650
rect 3516 70586 3568 70592
rect 3528 67658 3556 70586
rect 3516 67652 3568 67658
rect 3516 67594 3568 67600
rect 3712 65634 3740 71538
rect 3792 69760 3844 69766
rect 3792 69702 3844 69708
rect 3436 65606 3740 65634
rect 3436 61033 3464 65606
rect 3608 65544 3660 65550
rect 3608 65486 3660 65492
rect 3516 65068 3568 65074
rect 3516 65010 3568 65016
rect 3528 64870 3556 65010
rect 3516 64864 3568 64870
rect 3516 64806 3568 64812
rect 3516 64592 3568 64598
rect 3516 64534 3568 64540
rect 3528 62150 3556 64534
rect 3516 62144 3568 62150
rect 3516 62086 3568 62092
rect 3516 61804 3568 61810
rect 3516 61746 3568 61752
rect 3422 61024 3478 61033
rect 3422 60959 3478 60968
rect 3424 60716 3476 60722
rect 3424 60658 3476 60664
rect 3436 49638 3464 60658
rect 3528 58614 3556 61746
rect 3516 58608 3568 58614
rect 3516 58550 3568 58556
rect 3514 58440 3570 58449
rect 3514 58375 3516 58384
rect 3568 58375 3570 58384
rect 3516 58346 3568 58352
rect 3516 58132 3568 58138
rect 3516 58074 3568 58080
rect 3528 55865 3556 58074
rect 3620 56506 3648 65486
rect 3700 65408 3752 65414
rect 3700 65350 3752 65356
rect 3712 65142 3740 65350
rect 3700 65136 3752 65142
rect 3700 65078 3752 65084
rect 3700 63980 3752 63986
rect 3700 63922 3752 63928
rect 3712 61849 3740 63922
rect 3698 61840 3754 61849
rect 3698 61775 3754 61784
rect 3698 61704 3754 61713
rect 3698 61639 3700 61648
rect 3752 61639 3754 61648
rect 3700 61610 3752 61616
rect 3804 61554 3832 69702
rect 3712 61526 3832 61554
rect 3712 59430 3740 61526
rect 3790 61432 3846 61441
rect 3790 61367 3846 61376
rect 3700 59424 3752 59430
rect 3700 59366 3752 59372
rect 3700 58540 3752 58546
rect 3700 58482 3752 58488
rect 3608 56500 3660 56506
rect 3608 56442 3660 56448
rect 3608 56364 3660 56370
rect 3608 56306 3660 56312
rect 3514 55856 3570 55865
rect 3514 55791 3570 55800
rect 3516 55752 3568 55758
rect 3516 55694 3568 55700
rect 3528 55214 3556 55694
rect 3620 55418 3648 56306
rect 3608 55412 3660 55418
rect 3608 55354 3660 55360
rect 3608 55276 3660 55282
rect 3608 55218 3660 55224
rect 3516 55208 3568 55214
rect 3516 55150 3568 55156
rect 3528 55049 3556 55150
rect 3514 55040 3570 55049
rect 3514 54975 3570 54984
rect 3516 54868 3568 54874
rect 3516 54810 3568 54816
rect 3424 49632 3476 49638
rect 3528 49609 3556 54810
rect 3620 51474 3648 55218
rect 3608 51468 3660 51474
rect 3608 51410 3660 51416
rect 3606 51368 3662 51377
rect 3606 51303 3662 51312
rect 3424 49574 3476 49580
rect 3514 49600 3570 49609
rect 3514 49535 3570 49544
rect 3516 49428 3568 49434
rect 3516 49370 3568 49376
rect 3330 48784 3386 48793
rect 3330 48719 3386 48728
rect 3528 48634 3556 49370
rect 3436 48606 3556 48634
rect 3330 48104 3386 48113
rect 3330 48039 3386 48048
rect 3344 47444 3372 48039
rect 3436 47598 3464 48606
rect 3516 48544 3568 48550
rect 3516 48486 3568 48492
rect 3528 47841 3556 48486
rect 3514 47832 3570 47841
rect 3514 47767 3516 47776
rect 3568 47767 3570 47776
rect 3516 47738 3568 47744
rect 3620 47648 3648 51303
rect 3528 47620 3648 47648
rect 3424 47592 3476 47598
rect 3424 47534 3476 47540
rect 3344 47416 3464 47444
rect 3330 47288 3386 47297
rect 3330 47223 3386 47232
rect 3344 46510 3372 47223
rect 3332 46504 3384 46510
rect 3332 46446 3384 46452
rect 3252 46158 3372 46186
rect 3240 46096 3292 46102
rect 3240 46038 3292 46044
rect 3148 43852 3200 43858
rect 3148 43794 3200 43800
rect 3148 43648 3200 43654
rect 3148 43590 3200 43596
rect 3054 43480 3110 43489
rect 3054 43415 3110 43424
rect 2884 43302 3004 43330
rect 2780 43240 2832 43246
rect 2780 43182 2832 43188
rect 2516 43064 2636 43092
rect 2516 42888 2544 43064
rect 2582 43004 2890 43024
rect 2582 43002 2588 43004
rect 2644 43002 2668 43004
rect 2724 43002 2748 43004
rect 2804 43002 2828 43004
rect 2884 43002 2890 43004
rect 2644 42950 2646 43002
rect 2826 42950 2828 43002
rect 2582 42948 2588 42950
rect 2644 42948 2668 42950
rect 2724 42948 2748 42950
rect 2804 42948 2828 42950
rect 2884 42948 2890 42950
rect 2582 42928 2890 42948
rect 2516 42860 2728 42888
rect 2700 42294 2728 42860
rect 2778 42800 2834 42809
rect 2778 42735 2834 42744
rect 2688 42288 2740 42294
rect 2424 42214 2544 42242
rect 2688 42230 2740 42236
rect 2792 42226 2820 42735
rect 2976 42702 3004 43302
rect 3160 43217 3188 43590
rect 3146 43208 3202 43217
rect 3146 43143 3202 43152
rect 3056 43104 3108 43110
rect 3056 43046 3108 43052
rect 2964 42696 3016 42702
rect 2964 42638 3016 42644
rect 2964 42560 3016 42566
rect 2964 42502 3016 42508
rect 2516 41596 2544 42214
rect 2780 42220 2832 42226
rect 2780 42162 2832 42168
rect 2582 41916 2890 41936
rect 2582 41914 2588 41916
rect 2644 41914 2668 41916
rect 2724 41914 2748 41916
rect 2804 41914 2828 41916
rect 2884 41914 2890 41916
rect 2644 41862 2646 41914
rect 2826 41862 2828 41914
rect 2582 41860 2588 41862
rect 2644 41860 2668 41862
rect 2724 41860 2748 41862
rect 2804 41860 2828 41862
rect 2884 41860 2890 41862
rect 2582 41840 2890 41860
rect 2780 41744 2832 41750
rect 2976 41698 3004 42502
rect 2780 41686 2832 41692
rect 2516 41568 2636 41596
rect 2608 41274 2636 41568
rect 2688 41540 2740 41546
rect 2688 41482 2740 41488
rect 2412 41268 2464 41274
rect 2412 41210 2464 41216
rect 2596 41268 2648 41274
rect 2596 41210 2648 41216
rect 2424 38468 2452 41210
rect 2700 41138 2728 41482
rect 2792 41274 2820 41686
rect 2884 41670 3004 41698
rect 2780 41268 2832 41274
rect 2780 41210 2832 41216
rect 2688 41132 2740 41138
rect 2688 41074 2740 41080
rect 2884 41041 2912 41670
rect 3068 41562 3096 43046
rect 3148 42764 3200 42770
rect 3148 42706 3200 42712
rect 2976 41534 3096 41562
rect 2976 41177 3004 41534
rect 3160 41460 3188 42706
rect 3068 41432 3188 41460
rect 2962 41168 3018 41177
rect 2962 41103 3018 41112
rect 2870 41032 2926 41041
rect 2870 40967 2926 40976
rect 2582 40828 2890 40848
rect 2582 40826 2588 40828
rect 2644 40826 2668 40828
rect 2724 40826 2748 40828
rect 2804 40826 2828 40828
rect 2884 40826 2890 40828
rect 2644 40774 2646 40826
rect 2826 40774 2828 40826
rect 2582 40772 2588 40774
rect 2644 40772 2668 40774
rect 2724 40772 2748 40774
rect 2804 40772 2828 40774
rect 2884 40772 2890 40774
rect 2582 40752 2890 40772
rect 2594 40488 2650 40497
rect 2594 40423 2650 40432
rect 2608 39982 2636 40423
rect 2964 40112 3016 40118
rect 2964 40054 3016 40060
rect 2596 39976 2648 39982
rect 2596 39918 2648 39924
rect 2582 39740 2890 39760
rect 2582 39738 2588 39740
rect 2644 39738 2668 39740
rect 2724 39738 2748 39740
rect 2804 39738 2828 39740
rect 2884 39738 2890 39740
rect 2644 39686 2646 39738
rect 2826 39686 2828 39738
rect 2582 39684 2588 39686
rect 2644 39684 2668 39686
rect 2724 39684 2748 39686
rect 2804 39684 2828 39686
rect 2884 39684 2890 39686
rect 2582 39664 2890 39684
rect 2976 39438 3004 40054
rect 2780 39432 2832 39438
rect 2780 39374 2832 39380
rect 2964 39432 3016 39438
rect 2964 39374 3016 39380
rect 2504 39364 2556 39370
rect 2504 39306 2556 39312
rect 2516 38842 2544 39306
rect 2792 38865 2820 39374
rect 2976 38894 3004 39374
rect 3068 38944 3096 41432
rect 3252 40390 3280 46038
rect 3148 40384 3200 40390
rect 3148 40326 3200 40332
rect 3240 40384 3292 40390
rect 3240 40326 3292 40332
rect 3160 39642 3188 40326
rect 3344 40202 3372 46158
rect 3436 43790 3464 47416
rect 3424 43784 3476 43790
rect 3424 43726 3476 43732
rect 3424 43648 3476 43654
rect 3422 43616 3424 43625
rect 3476 43616 3478 43625
rect 3422 43551 3478 43560
rect 3424 43240 3476 43246
rect 3424 43182 3476 43188
rect 3436 42650 3464 43182
rect 3528 42770 3556 47620
rect 3712 47580 3740 58482
rect 3804 50017 3832 61367
rect 3790 50008 3846 50017
rect 3790 49943 3846 49952
rect 3792 49768 3844 49774
rect 3792 49710 3844 49716
rect 3804 48668 3832 49710
rect 3896 49434 3924 72422
rect 4632 71942 4660 72422
rect 4620 71936 4672 71942
rect 4620 71878 4672 71884
rect 4214 71836 4522 71856
rect 4214 71834 4220 71836
rect 4276 71834 4300 71836
rect 4356 71834 4380 71836
rect 4436 71834 4460 71836
rect 4516 71834 4522 71836
rect 4276 71782 4278 71834
rect 4458 71782 4460 71834
rect 4214 71780 4220 71782
rect 4276 71780 4300 71782
rect 4356 71780 4380 71782
rect 4436 71780 4460 71782
rect 4516 71780 4522 71782
rect 4214 71760 4522 71780
rect 4214 70748 4522 70768
rect 4214 70746 4220 70748
rect 4276 70746 4300 70748
rect 4356 70746 4380 70748
rect 4436 70746 4460 70748
rect 4516 70746 4522 70748
rect 4276 70694 4278 70746
rect 4458 70694 4460 70746
rect 4214 70692 4220 70694
rect 4276 70692 4300 70694
rect 4356 70692 4380 70694
rect 4436 70692 4460 70694
rect 4516 70692 4522 70694
rect 4214 70672 4522 70692
rect 4214 69660 4522 69680
rect 4214 69658 4220 69660
rect 4276 69658 4300 69660
rect 4356 69658 4380 69660
rect 4436 69658 4460 69660
rect 4516 69658 4522 69660
rect 4276 69606 4278 69658
rect 4458 69606 4460 69658
rect 4214 69604 4220 69606
rect 4276 69604 4300 69606
rect 4356 69604 4380 69606
rect 4436 69604 4460 69606
rect 4516 69604 4522 69606
rect 4214 69584 4522 69604
rect 4068 68944 4120 68950
rect 4068 68886 4120 68892
rect 3976 65408 4028 65414
rect 3976 65350 4028 65356
rect 3988 65113 4016 65350
rect 3974 65104 4030 65113
rect 3974 65039 4030 65048
rect 4080 64546 4108 68886
rect 4214 68572 4522 68592
rect 4214 68570 4220 68572
rect 4276 68570 4300 68572
rect 4356 68570 4380 68572
rect 4436 68570 4460 68572
rect 4516 68570 4522 68572
rect 4276 68518 4278 68570
rect 4458 68518 4460 68570
rect 4214 68516 4220 68518
rect 4276 68516 4300 68518
rect 4356 68516 4380 68518
rect 4436 68516 4460 68518
rect 4516 68516 4522 68518
rect 4214 68496 4522 68516
rect 4804 67652 4856 67658
rect 4804 67594 4856 67600
rect 4214 67484 4522 67504
rect 4214 67482 4220 67484
rect 4276 67482 4300 67484
rect 4356 67482 4380 67484
rect 4436 67482 4460 67484
rect 4516 67482 4522 67484
rect 4276 67430 4278 67482
rect 4458 67430 4460 67482
rect 4214 67428 4220 67430
rect 4276 67428 4300 67430
rect 4356 67428 4380 67430
rect 4436 67428 4460 67430
rect 4516 67428 4522 67430
rect 4214 67408 4522 67428
rect 4214 66396 4522 66416
rect 4214 66394 4220 66396
rect 4276 66394 4300 66396
rect 4356 66394 4380 66396
rect 4436 66394 4460 66396
rect 4516 66394 4522 66396
rect 4276 66342 4278 66394
rect 4458 66342 4460 66394
rect 4214 66340 4220 66342
rect 4276 66340 4300 66342
rect 4356 66340 4380 66342
rect 4436 66340 4460 66342
rect 4516 66340 4522 66342
rect 4214 66320 4522 66340
rect 4214 65308 4522 65328
rect 4214 65306 4220 65308
rect 4276 65306 4300 65308
rect 4356 65306 4380 65308
rect 4436 65306 4460 65308
rect 4516 65306 4522 65308
rect 4276 65254 4278 65306
rect 4458 65254 4460 65306
rect 4214 65252 4220 65254
rect 4276 65252 4300 65254
rect 4356 65252 4380 65254
rect 4436 65252 4460 65254
rect 4516 65252 4522 65254
rect 4214 65232 4522 65252
rect 3988 64518 4108 64546
rect 3988 61441 4016 64518
rect 4068 64456 4120 64462
rect 4068 64398 4120 64404
rect 3974 61432 4030 61441
rect 3974 61367 4030 61376
rect 3976 60648 4028 60654
rect 4080 60625 4108 64398
rect 4214 64220 4522 64240
rect 4214 64218 4220 64220
rect 4276 64218 4300 64220
rect 4356 64218 4380 64220
rect 4436 64218 4460 64220
rect 4516 64218 4522 64220
rect 4276 64166 4278 64218
rect 4458 64166 4460 64218
rect 4214 64164 4220 64166
rect 4276 64164 4300 64166
rect 4356 64164 4380 64166
rect 4436 64164 4460 64166
rect 4516 64164 4522 64166
rect 4214 64144 4522 64164
rect 4214 63132 4522 63152
rect 4214 63130 4220 63132
rect 4276 63130 4300 63132
rect 4356 63130 4380 63132
rect 4436 63130 4460 63132
rect 4516 63130 4522 63132
rect 4276 63078 4278 63130
rect 4458 63078 4460 63130
rect 4214 63076 4220 63078
rect 4276 63076 4300 63078
rect 4356 63076 4380 63078
rect 4436 63076 4460 63078
rect 4516 63076 4522 63078
rect 4214 63056 4522 63076
rect 4214 62044 4522 62064
rect 4214 62042 4220 62044
rect 4276 62042 4300 62044
rect 4356 62042 4380 62044
rect 4436 62042 4460 62044
rect 4516 62042 4522 62044
rect 4276 61990 4278 62042
rect 4458 61990 4460 62042
rect 4214 61988 4220 61990
rect 4276 61988 4300 61990
rect 4356 61988 4380 61990
rect 4436 61988 4460 61990
rect 4516 61988 4522 61990
rect 4214 61968 4522 61988
rect 4214 60956 4522 60976
rect 4214 60954 4220 60956
rect 4276 60954 4300 60956
rect 4356 60954 4380 60956
rect 4436 60954 4460 60956
rect 4516 60954 4522 60956
rect 4276 60902 4278 60954
rect 4458 60902 4460 60954
rect 4214 60900 4220 60902
rect 4276 60900 4300 60902
rect 4356 60900 4380 60902
rect 4436 60900 4460 60902
rect 4516 60900 4522 60902
rect 4214 60880 4522 60900
rect 3976 60590 4028 60596
rect 4066 60616 4122 60625
rect 3988 59430 4016 60590
rect 4066 60551 4122 60560
rect 4066 60480 4122 60489
rect 4066 60415 4122 60424
rect 3976 59424 4028 59430
rect 3976 59366 4028 59372
rect 3976 58880 4028 58886
rect 3976 58822 4028 58828
rect 3988 58721 4016 58822
rect 3974 58712 4030 58721
rect 3974 58647 4030 58656
rect 3976 58608 4028 58614
rect 3976 58550 4028 58556
rect 3988 49774 4016 58550
rect 4080 54874 4108 60415
rect 4214 59868 4522 59888
rect 4214 59866 4220 59868
rect 4276 59866 4300 59868
rect 4356 59866 4380 59868
rect 4436 59866 4460 59868
rect 4516 59866 4522 59868
rect 4276 59814 4278 59866
rect 4458 59814 4460 59866
rect 4214 59812 4220 59814
rect 4276 59812 4300 59814
rect 4356 59812 4380 59814
rect 4436 59812 4460 59814
rect 4516 59812 4522 59814
rect 4214 59792 4522 59812
rect 4620 59424 4672 59430
rect 4620 59366 4672 59372
rect 4214 58780 4522 58800
rect 4214 58778 4220 58780
rect 4276 58778 4300 58780
rect 4356 58778 4380 58780
rect 4436 58778 4460 58780
rect 4516 58778 4522 58780
rect 4276 58726 4278 58778
rect 4458 58726 4460 58778
rect 4214 58724 4220 58726
rect 4276 58724 4300 58726
rect 4356 58724 4380 58726
rect 4436 58724 4460 58726
rect 4516 58724 4522 58726
rect 4214 58704 4522 58724
rect 4160 58472 4212 58478
rect 4160 58414 4212 58420
rect 4172 58138 4200 58414
rect 4160 58132 4212 58138
rect 4160 58074 4212 58080
rect 4214 57692 4522 57712
rect 4214 57690 4220 57692
rect 4276 57690 4300 57692
rect 4356 57690 4380 57692
rect 4436 57690 4460 57692
rect 4516 57690 4522 57692
rect 4276 57638 4278 57690
rect 4458 57638 4460 57690
rect 4214 57636 4220 57638
rect 4276 57636 4300 57638
rect 4356 57636 4380 57638
rect 4436 57636 4460 57638
rect 4516 57636 4522 57638
rect 4214 57616 4522 57636
rect 4214 56604 4522 56624
rect 4214 56602 4220 56604
rect 4276 56602 4300 56604
rect 4356 56602 4380 56604
rect 4436 56602 4460 56604
rect 4516 56602 4522 56604
rect 4276 56550 4278 56602
rect 4458 56550 4460 56602
rect 4214 56548 4220 56550
rect 4276 56548 4300 56550
rect 4356 56548 4380 56550
rect 4436 56548 4460 56550
rect 4516 56548 4522 56550
rect 4214 56528 4522 56548
rect 4160 55752 4212 55758
rect 4158 55720 4160 55729
rect 4212 55720 4214 55729
rect 4158 55655 4214 55664
rect 4214 55516 4522 55536
rect 4214 55514 4220 55516
rect 4276 55514 4300 55516
rect 4356 55514 4380 55516
rect 4436 55514 4460 55516
rect 4516 55514 4522 55516
rect 4276 55462 4278 55514
rect 4458 55462 4460 55514
rect 4214 55460 4220 55462
rect 4276 55460 4300 55462
rect 4356 55460 4380 55462
rect 4436 55460 4460 55462
rect 4516 55460 4522 55462
rect 4214 55440 4522 55460
rect 4632 55298 4660 59366
rect 4712 59016 4764 59022
rect 4712 58958 4764 58964
rect 4172 55270 4660 55298
rect 4068 54868 4120 54874
rect 4068 54810 4120 54816
rect 4172 54754 4200 55270
rect 4344 55208 4396 55214
rect 4342 55176 4344 55185
rect 4396 55176 4398 55185
rect 4342 55111 4398 55120
rect 4080 54726 4200 54754
rect 4080 50969 4108 54726
rect 4214 54428 4522 54448
rect 4214 54426 4220 54428
rect 4276 54426 4300 54428
rect 4356 54426 4380 54428
rect 4436 54426 4460 54428
rect 4516 54426 4522 54428
rect 4276 54374 4278 54426
rect 4458 54374 4460 54426
rect 4214 54372 4220 54374
rect 4276 54372 4300 54374
rect 4356 54372 4380 54374
rect 4436 54372 4460 54374
rect 4516 54372 4522 54374
rect 4214 54352 4522 54372
rect 4620 53576 4672 53582
rect 4620 53518 4672 53524
rect 4214 53340 4522 53360
rect 4214 53338 4220 53340
rect 4276 53338 4300 53340
rect 4356 53338 4380 53340
rect 4436 53338 4460 53340
rect 4516 53338 4522 53340
rect 4276 53286 4278 53338
rect 4458 53286 4460 53338
rect 4214 53284 4220 53286
rect 4276 53284 4300 53286
rect 4356 53284 4380 53286
rect 4436 53284 4460 53286
rect 4516 53284 4522 53286
rect 4214 53264 4522 53284
rect 4158 52728 4214 52737
rect 4158 52663 4160 52672
rect 4212 52663 4214 52672
rect 4160 52634 4212 52640
rect 4214 52252 4522 52272
rect 4214 52250 4220 52252
rect 4276 52250 4300 52252
rect 4356 52250 4380 52252
rect 4436 52250 4460 52252
rect 4516 52250 4522 52252
rect 4276 52198 4278 52250
rect 4458 52198 4460 52250
rect 4214 52196 4220 52198
rect 4276 52196 4300 52198
rect 4356 52196 4380 52198
rect 4436 52196 4460 52198
rect 4516 52196 4522 52198
rect 4214 52176 4522 52196
rect 4632 51513 4660 53518
rect 4724 53174 4752 58958
rect 4712 53168 4764 53174
rect 4712 53110 4764 53116
rect 4816 52986 4844 67594
rect 5172 66768 5224 66774
rect 5172 66710 5224 66716
rect 4988 66020 5040 66026
rect 4988 65962 5040 65968
rect 4896 65136 4948 65142
rect 4896 65078 4948 65084
rect 4724 52958 4844 52986
rect 4618 51504 4674 51513
rect 4618 51439 4674 51448
rect 4214 51164 4522 51184
rect 4214 51162 4220 51164
rect 4276 51162 4300 51164
rect 4356 51162 4380 51164
rect 4436 51162 4460 51164
rect 4516 51162 4522 51164
rect 4276 51110 4278 51162
rect 4458 51110 4460 51162
rect 4724 51116 4752 52958
rect 4802 52864 4858 52873
rect 4802 52799 4858 52808
rect 4214 51108 4220 51110
rect 4276 51108 4300 51110
rect 4356 51108 4380 51110
rect 4436 51108 4460 51110
rect 4516 51108 4522 51110
rect 4214 51088 4522 51108
rect 4632 51088 4752 51116
rect 4066 50960 4122 50969
rect 4632 50946 4660 51088
rect 4066 50895 4122 50904
rect 4160 50924 4212 50930
rect 4632 50918 4752 50946
rect 4816 50930 4844 52799
rect 4160 50866 4212 50872
rect 4068 50856 4120 50862
rect 4068 50798 4120 50804
rect 3976 49768 4028 49774
rect 3976 49710 4028 49716
rect 3976 49632 4028 49638
rect 3976 49574 4028 49580
rect 3884 49428 3936 49434
rect 3884 49370 3936 49376
rect 3804 48640 3924 48668
rect 3790 48240 3846 48249
rect 3790 48175 3846 48184
rect 3620 47552 3740 47580
rect 3516 42764 3568 42770
rect 3516 42706 3568 42712
rect 3436 42622 3556 42650
rect 3424 42560 3476 42566
rect 3424 42502 3476 42508
rect 3436 41721 3464 42502
rect 3422 41712 3478 41721
rect 3422 41647 3478 41656
rect 3424 41608 3476 41614
rect 3528 41585 3556 42622
rect 3424 41550 3476 41556
rect 3514 41576 3570 41585
rect 3436 41041 3464 41550
rect 3514 41511 3570 41520
rect 3516 41472 3568 41478
rect 3620 41449 3648 47552
rect 3700 47456 3752 47462
rect 3700 47398 3752 47404
rect 3712 47161 3740 47398
rect 3698 47152 3754 47161
rect 3698 47087 3754 47096
rect 3698 46608 3754 46617
rect 3698 46543 3700 46552
rect 3752 46543 3754 46552
rect 3700 46514 3752 46520
rect 3804 46186 3832 48175
rect 3896 47734 3924 48640
rect 3884 47728 3936 47734
rect 3884 47670 3936 47676
rect 3884 47592 3936 47598
rect 3884 47534 3936 47540
rect 3896 47161 3924 47534
rect 3882 47152 3938 47161
rect 3882 47087 3938 47096
rect 3988 47036 4016 49574
rect 3896 47008 4016 47036
rect 3896 46560 3924 47008
rect 3976 46912 4028 46918
rect 3976 46854 4028 46860
rect 3988 46753 4016 46854
rect 3974 46744 4030 46753
rect 3974 46679 4030 46688
rect 3896 46532 4016 46560
rect 3882 46472 3938 46481
rect 3882 46407 3884 46416
rect 3936 46407 3938 46416
rect 3884 46378 3936 46384
rect 3712 46158 3832 46186
rect 3516 41414 3568 41420
rect 3606 41440 3662 41449
rect 3528 41274 3556 41414
rect 3606 41375 3662 41384
rect 3606 41304 3662 41313
rect 3516 41268 3568 41274
rect 3606 41239 3662 41248
rect 3516 41210 3568 41216
rect 3514 41168 3570 41177
rect 3514 41103 3570 41112
rect 3422 41032 3478 41041
rect 3422 40967 3478 40976
rect 3424 40928 3476 40934
rect 3424 40870 3476 40876
rect 3436 40497 3464 40870
rect 3422 40488 3478 40497
rect 3422 40423 3478 40432
rect 3424 40384 3476 40390
rect 3424 40326 3476 40332
rect 3252 40174 3372 40202
rect 3148 39636 3200 39642
rect 3148 39578 3200 39584
rect 3252 39030 3280 40174
rect 3330 39944 3386 39953
rect 3330 39879 3332 39888
rect 3384 39879 3386 39888
rect 3332 39850 3384 39856
rect 3332 39568 3384 39574
rect 3332 39510 3384 39516
rect 3240 39024 3292 39030
rect 3240 38966 3292 38972
rect 3068 38916 3188 38944
rect 2964 38888 3016 38894
rect 2594 38856 2650 38865
rect 2516 38814 2594 38842
rect 2594 38791 2650 38800
rect 2778 38856 2834 38865
rect 2964 38830 3016 38836
rect 2778 38791 2834 38800
rect 3056 38820 3108 38826
rect 3056 38762 3108 38768
rect 3068 38706 3096 38762
rect 3160 38729 3188 38916
rect 2976 38678 3096 38706
rect 3146 38720 3202 38729
rect 2582 38652 2890 38672
rect 2582 38650 2588 38652
rect 2644 38650 2668 38652
rect 2724 38650 2748 38652
rect 2804 38650 2828 38652
rect 2884 38650 2890 38652
rect 2644 38598 2646 38650
rect 2826 38598 2828 38650
rect 2582 38596 2588 38598
rect 2644 38596 2668 38598
rect 2724 38596 2748 38598
rect 2804 38596 2828 38598
rect 2884 38596 2890 38598
rect 2582 38576 2890 38596
rect 2976 38554 3004 38678
rect 3146 38655 3202 38664
rect 3146 38584 3202 38593
rect 2964 38548 3016 38554
rect 3146 38519 3148 38528
rect 2964 38490 3016 38496
rect 3200 38519 3202 38528
rect 3148 38490 3200 38496
rect 3056 38480 3108 38486
rect 2424 38440 2636 38468
rect 2332 38372 2452 38400
rect 1952 38354 2004 38360
rect 1860 38276 1912 38282
rect 1860 38218 1912 38224
rect 1858 37904 1914 37913
rect 1858 37839 1914 37848
rect 1872 37398 1900 37839
rect 1964 37806 1992 38354
rect 2136 38276 2188 38282
rect 2136 38218 2188 38224
rect 2320 38276 2372 38282
rect 2320 38218 2372 38224
rect 2044 38208 2096 38214
rect 2044 38150 2096 38156
rect 1952 37800 2004 37806
rect 1952 37742 2004 37748
rect 1952 37664 2004 37670
rect 1952 37606 2004 37612
rect 1860 37392 1912 37398
rect 1860 37334 1912 37340
rect 1860 36712 1912 36718
rect 1860 36654 1912 36660
rect 1872 31958 1900 36654
rect 1860 31952 1912 31958
rect 1860 31894 1912 31900
rect 1860 31748 1912 31754
rect 1860 31690 1912 31696
rect 1872 31482 1900 31690
rect 1860 31476 1912 31482
rect 1860 31418 1912 31424
rect 1768 30728 1820 30734
rect 1768 30670 1820 30676
rect 1860 30660 1912 30666
rect 1860 30602 1912 30608
rect 1688 30382 1808 30410
rect 1676 30252 1728 30258
rect 1676 30194 1728 30200
rect 1688 29209 1716 30194
rect 1674 29200 1730 29209
rect 1674 29135 1730 29144
rect 1676 28212 1728 28218
rect 1676 28154 1728 28160
rect 1688 23730 1716 28154
rect 1780 25906 1808 30382
rect 1872 30161 1900 30602
rect 1858 30152 1914 30161
rect 1858 30087 1914 30096
rect 1860 30048 1912 30054
rect 1860 29990 1912 29996
rect 1872 26897 1900 29990
rect 1964 28082 1992 37606
rect 2056 34610 2084 38150
rect 2044 34604 2096 34610
rect 2044 34546 2096 34552
rect 2044 34468 2096 34474
rect 2044 34410 2096 34416
rect 2056 30326 2084 34410
rect 2148 32910 2176 38218
rect 2228 38208 2280 38214
rect 2332 38185 2360 38218
rect 2228 38150 2280 38156
rect 2318 38176 2374 38185
rect 2240 37466 2268 38150
rect 2318 38111 2374 38120
rect 2320 37800 2372 37806
rect 2320 37742 2372 37748
rect 2228 37460 2280 37466
rect 2228 37402 2280 37408
rect 2332 37194 2360 37742
rect 2228 37188 2280 37194
rect 2228 37130 2280 37136
rect 2320 37188 2372 37194
rect 2320 37130 2372 37136
rect 2240 34474 2268 37130
rect 2320 36916 2372 36922
rect 2320 36858 2372 36864
rect 2332 36553 2360 36858
rect 2318 36544 2374 36553
rect 2318 36479 2374 36488
rect 2318 35592 2374 35601
rect 2318 35527 2320 35536
rect 2372 35527 2374 35536
rect 2320 35498 2372 35504
rect 2424 35086 2452 38372
rect 2504 38344 2556 38350
rect 2504 38286 2556 38292
rect 2516 37466 2544 38286
rect 2608 37874 2636 38440
rect 2778 38448 2834 38457
rect 3056 38422 3108 38428
rect 2778 38383 2834 38392
rect 2688 38208 2740 38214
rect 2688 38150 2740 38156
rect 2596 37868 2648 37874
rect 2596 37810 2648 37816
rect 2700 37806 2728 38150
rect 2792 38010 2820 38383
rect 2964 38276 3016 38282
rect 2964 38218 3016 38224
rect 2780 38004 2832 38010
rect 2780 37946 2832 37952
rect 2976 37942 3004 38218
rect 2964 37936 3016 37942
rect 2964 37878 3016 37884
rect 2688 37800 2740 37806
rect 2688 37742 2740 37748
rect 2582 37564 2890 37584
rect 2582 37562 2588 37564
rect 2644 37562 2668 37564
rect 2724 37562 2748 37564
rect 2804 37562 2828 37564
rect 2884 37562 2890 37564
rect 2644 37510 2646 37562
rect 2826 37510 2828 37562
rect 2582 37508 2588 37510
rect 2644 37508 2668 37510
rect 2724 37508 2748 37510
rect 2804 37508 2828 37510
rect 2884 37508 2890 37510
rect 2582 37488 2890 37508
rect 2504 37460 2556 37466
rect 2504 37402 2556 37408
rect 2516 36786 2544 37402
rect 2688 37188 2740 37194
rect 2688 37130 2740 37136
rect 2700 36922 2728 37130
rect 2976 37126 3004 37878
rect 2964 37120 3016 37126
rect 2964 37062 3016 37068
rect 2688 36916 2740 36922
rect 2688 36858 2740 36864
rect 2872 36848 2924 36854
rect 2872 36790 2924 36796
rect 2504 36780 2556 36786
rect 2504 36722 2556 36728
rect 2884 36666 2912 36790
rect 2884 36638 3004 36666
rect 2504 36576 2556 36582
rect 2504 36518 2556 36524
rect 2516 36174 2544 36518
rect 2582 36476 2890 36496
rect 2582 36474 2588 36476
rect 2644 36474 2668 36476
rect 2724 36474 2748 36476
rect 2804 36474 2828 36476
rect 2884 36474 2890 36476
rect 2644 36422 2646 36474
rect 2826 36422 2828 36474
rect 2582 36420 2588 36422
rect 2644 36420 2668 36422
rect 2724 36420 2748 36422
rect 2804 36420 2828 36422
rect 2884 36420 2890 36422
rect 2582 36400 2890 36420
rect 2976 36394 3004 36638
rect 3068 36582 3096 38422
rect 3344 38321 3372 39510
rect 3330 38312 3386 38321
rect 3330 38247 3386 38256
rect 3436 38026 3464 40326
rect 3252 37998 3464 38026
rect 3146 37904 3202 37913
rect 3146 37839 3202 37848
rect 3056 36576 3108 36582
rect 3056 36518 3108 36524
rect 2976 36366 3096 36394
rect 2504 36168 2556 36174
rect 2504 36110 2556 36116
rect 2962 36136 3018 36145
rect 2962 36071 3018 36080
rect 2582 35388 2890 35408
rect 2582 35386 2588 35388
rect 2644 35386 2668 35388
rect 2724 35386 2748 35388
rect 2804 35386 2828 35388
rect 2884 35386 2890 35388
rect 2644 35334 2646 35386
rect 2826 35334 2828 35386
rect 2582 35332 2588 35334
rect 2644 35332 2668 35334
rect 2724 35332 2748 35334
rect 2804 35332 2828 35334
rect 2884 35332 2890 35334
rect 2582 35312 2890 35332
rect 2412 35080 2464 35086
rect 2412 35022 2464 35028
rect 2504 35012 2556 35018
rect 2504 34954 2556 34960
rect 2228 34468 2280 34474
rect 2228 34410 2280 34416
rect 2412 33992 2464 33998
rect 2412 33934 2464 33940
rect 2228 33924 2280 33930
rect 2228 33866 2280 33872
rect 2320 33924 2372 33930
rect 2320 33866 2372 33872
rect 2240 33658 2268 33866
rect 2228 33652 2280 33658
rect 2228 33594 2280 33600
rect 2332 33590 2360 33866
rect 2320 33584 2372 33590
rect 2320 33526 2372 33532
rect 2228 33516 2280 33522
rect 2228 33458 2280 33464
rect 2136 32904 2188 32910
rect 2136 32846 2188 32852
rect 2134 32736 2190 32745
rect 2134 32671 2190 32680
rect 2148 31906 2176 32671
rect 2240 32434 2268 33458
rect 2320 32768 2372 32774
rect 2320 32710 2372 32716
rect 2332 32609 2360 32710
rect 2318 32600 2374 32609
rect 2318 32535 2374 32544
rect 2228 32428 2280 32434
rect 2280 32388 2360 32416
rect 2228 32370 2280 32376
rect 2148 31890 2268 31906
rect 2148 31884 2280 31890
rect 2148 31878 2228 31884
rect 2228 31826 2280 31832
rect 2136 31816 2188 31822
rect 2136 31758 2188 31764
rect 2044 30320 2096 30326
rect 2044 30262 2096 30268
rect 2042 30152 2098 30161
rect 2042 30087 2098 30096
rect 1952 28076 2004 28082
rect 1952 28018 2004 28024
rect 1952 27940 2004 27946
rect 1952 27882 2004 27888
rect 1964 27470 1992 27882
rect 1952 27464 2004 27470
rect 1952 27406 2004 27412
rect 1964 26994 1992 27406
rect 1952 26988 2004 26994
rect 1952 26930 2004 26936
rect 1858 26888 1914 26897
rect 1858 26823 1914 26832
rect 1952 26852 2004 26858
rect 1952 26794 2004 26800
rect 1860 26784 1912 26790
rect 1860 26726 1912 26732
rect 1872 26382 1900 26726
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 1860 26240 1912 26246
rect 1860 26182 1912 26188
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 1768 25764 1820 25770
rect 1768 25706 1820 25712
rect 1780 24070 1808 25706
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1766 23896 1822 23905
rect 1766 23831 1822 23840
rect 1676 23724 1728 23730
rect 1676 23666 1728 23672
rect 1676 22500 1728 22506
rect 1676 22442 1728 22448
rect 1504 20998 1624 21026
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 20641 1440 20878
rect 1398 20632 1454 20641
rect 1398 20567 1454 20576
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1412 20233 1440 20334
rect 1398 20224 1454 20233
rect 1398 20159 1454 20168
rect 1400 19168 1452 19174
rect 1400 19110 1452 19116
rect 1412 18426 1440 19110
rect 1504 18850 1532 20998
rect 1584 20936 1636 20942
rect 1688 20924 1716 22442
rect 1780 22166 1808 23831
rect 1768 22160 1820 22166
rect 1768 22102 1820 22108
rect 1768 21480 1820 21486
rect 1768 21422 1820 21428
rect 1636 20896 1716 20924
rect 1584 20878 1636 20884
rect 1596 18970 1624 20878
rect 1780 20482 1808 21422
rect 1688 20454 1808 20482
rect 1688 19174 1716 20454
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 1780 19854 1808 20334
rect 1872 19990 1900 26182
rect 1860 19984 1912 19990
rect 1860 19926 1912 19932
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1504 18822 1716 18850
rect 1492 18760 1544 18766
rect 1492 18702 1544 18708
rect 1400 18420 1452 18426
rect 1400 18362 1452 18368
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1136 17224 1348 17252
rect 1412 17241 1440 18226
rect 1504 17649 1532 18702
rect 1584 17672 1636 17678
rect 1490 17640 1546 17649
rect 1584 17614 1636 17620
rect 1490 17575 1546 17584
rect 1398 17232 1454 17241
rect 1136 12102 1164 17224
rect 1398 17167 1454 17176
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16114 1440 16934
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1504 15609 1532 17138
rect 1596 16833 1624 17614
rect 1582 16824 1638 16833
rect 1582 16759 1638 16768
rect 1584 16720 1636 16726
rect 1584 16662 1636 16668
rect 1490 15600 1546 15609
rect 1490 15535 1546 15544
rect 1492 14068 1544 14074
rect 1492 14010 1544 14016
rect 1308 13320 1360 13326
rect 1308 13262 1360 13268
rect 1216 12844 1268 12850
rect 1216 12786 1268 12792
rect 1124 12096 1176 12102
rect 1124 12038 1176 12044
rect 1032 11756 1084 11762
rect 1032 11698 1084 11704
rect 1228 11257 1256 12786
rect 1320 11801 1348 13262
rect 1400 13184 1452 13190
rect 1400 13126 1452 13132
rect 1412 12442 1440 13126
rect 1400 12436 1452 12442
rect 1400 12378 1452 12384
rect 1504 12238 1532 14010
rect 1596 13954 1624 16662
rect 1688 14793 1716 18822
rect 1780 17882 1808 19790
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1872 19446 1900 19654
rect 1964 19514 1992 26794
rect 2056 24274 2084 30087
rect 2148 26858 2176 31758
rect 2228 31748 2280 31754
rect 2228 31690 2280 31696
rect 2136 26852 2188 26858
rect 2136 26794 2188 26800
rect 2134 26752 2190 26761
rect 2134 26687 2190 26696
rect 2044 24268 2096 24274
rect 2044 24210 2096 24216
rect 2148 24154 2176 26687
rect 2056 24126 2176 24154
rect 2056 22137 2084 24126
rect 2136 24064 2188 24070
rect 2136 24006 2188 24012
rect 2042 22128 2098 22137
rect 2042 22063 2098 22072
rect 2044 22024 2096 22030
rect 2044 21966 2096 21972
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1860 19440 1912 19446
rect 1860 19382 1912 19388
rect 2056 18970 2084 21966
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1872 16726 1900 18022
rect 1860 16720 1912 16726
rect 1860 16662 1912 16668
rect 2044 16516 2096 16522
rect 2044 16458 2096 16464
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1674 14784 1730 14793
rect 1674 14719 1730 14728
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1688 14074 1716 14554
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1596 13926 1716 13954
rect 1584 13796 1636 13802
rect 1584 13738 1636 13744
rect 1596 12617 1624 13738
rect 1582 12608 1638 12617
rect 1582 12543 1638 12552
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1306 11792 1362 11801
rect 1306 11727 1362 11736
rect 1308 11688 1360 11694
rect 1308 11630 1360 11636
rect 1214 11248 1270 11257
rect 1214 11183 1270 11192
rect 1320 10849 1348 11630
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1306 10840 1362 10849
rect 1306 10775 1362 10784
rect 1308 10600 1360 10606
rect 1308 10542 1360 10548
rect 1320 10033 1348 10542
rect 1412 10441 1440 11086
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 1400 10056 1452 10062
rect 1306 10024 1362 10033
rect 1400 9998 1452 10004
rect 1306 9959 1362 9968
rect 1412 9625 1440 9998
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 9217 1440 9454
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 8673 1440 8910
rect 1398 8664 1454 8673
rect 1398 8599 1454 8608
rect 1596 8566 1624 12271
rect 1688 11218 1716 13926
rect 1780 12442 1808 15438
rect 1872 14618 1900 15642
rect 1964 15570 1992 15846
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1964 14464 1992 14554
rect 1872 14436 1992 14464
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8265 1440 8366
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1400 7880 1452 7886
rect 1398 7848 1400 7857
rect 1452 7848 1454 7857
rect 1398 7783 1454 7792
rect 1398 7440 1454 7449
rect 1398 7375 1400 7384
rect 1452 7375 1454 7384
rect 1400 7346 1452 7352
rect 1596 6882 1624 8502
rect 1780 8498 1808 11494
rect 1872 9586 1900 14436
rect 1950 14376 2006 14385
rect 1950 14311 2006 14320
rect 1964 12866 1992 14311
rect 2056 13161 2084 16458
rect 2148 15162 2176 24006
rect 2240 22098 2268 31690
rect 2332 31686 2360 32388
rect 2320 31680 2372 31686
rect 2320 31622 2372 31628
rect 2320 31476 2372 31482
rect 2320 31418 2372 31424
rect 2332 30297 2360 31418
rect 2424 31328 2452 33934
rect 2516 33590 2544 34954
rect 2780 34944 2832 34950
rect 2780 34886 2832 34892
rect 2792 34513 2820 34886
rect 2976 34610 3004 36071
rect 2964 34604 3016 34610
rect 2964 34546 3016 34552
rect 2778 34504 2834 34513
rect 3068 34490 3096 36366
rect 2778 34439 2834 34448
rect 2976 34462 3096 34490
rect 2582 34300 2890 34320
rect 2582 34298 2588 34300
rect 2644 34298 2668 34300
rect 2724 34298 2748 34300
rect 2804 34298 2828 34300
rect 2884 34298 2890 34300
rect 2644 34246 2646 34298
rect 2826 34246 2828 34298
rect 2582 34244 2588 34246
rect 2644 34244 2668 34246
rect 2724 34244 2748 34246
rect 2804 34244 2828 34246
rect 2884 34244 2890 34246
rect 2582 34224 2890 34244
rect 2872 33992 2924 33998
rect 2872 33934 2924 33940
rect 2504 33584 2556 33590
rect 2504 33526 2556 33532
rect 2504 33448 2556 33454
rect 2504 33390 2556 33396
rect 2516 32026 2544 33390
rect 2884 33386 2912 33934
rect 2976 33810 3004 34462
rect 3056 34400 3108 34406
rect 3056 34342 3108 34348
rect 3068 33969 3096 34342
rect 3054 33960 3110 33969
rect 3054 33895 3110 33904
rect 2976 33782 3096 33810
rect 3068 33522 3096 33782
rect 2964 33516 3016 33522
rect 2964 33458 3016 33464
rect 3056 33516 3108 33522
rect 3056 33458 3108 33464
rect 2872 33380 2924 33386
rect 2872 33322 2924 33328
rect 2582 33212 2890 33232
rect 2582 33210 2588 33212
rect 2644 33210 2668 33212
rect 2724 33210 2748 33212
rect 2804 33210 2828 33212
rect 2884 33210 2890 33212
rect 2644 33158 2646 33210
rect 2826 33158 2828 33210
rect 2582 33156 2588 33158
rect 2644 33156 2668 33158
rect 2724 33156 2748 33158
rect 2804 33156 2828 33158
rect 2884 33156 2890 33158
rect 2582 33136 2890 33156
rect 2778 32872 2834 32881
rect 2778 32807 2834 32816
rect 2792 32774 2820 32807
rect 2780 32768 2832 32774
rect 2780 32710 2832 32716
rect 2976 32570 3004 33458
rect 3056 33380 3108 33386
rect 3056 33322 3108 33328
rect 2964 32564 3016 32570
rect 2964 32506 3016 32512
rect 3068 32416 3096 33322
rect 2976 32388 3096 32416
rect 2582 32124 2890 32144
rect 2582 32122 2588 32124
rect 2644 32122 2668 32124
rect 2724 32122 2748 32124
rect 2804 32122 2828 32124
rect 2884 32122 2890 32124
rect 2644 32070 2646 32122
rect 2826 32070 2828 32122
rect 2582 32068 2588 32070
rect 2644 32068 2668 32070
rect 2724 32068 2748 32070
rect 2804 32068 2828 32070
rect 2884 32068 2890 32070
rect 2582 32048 2890 32068
rect 2504 32020 2556 32026
rect 2504 31962 2556 31968
rect 2596 31952 2648 31958
rect 2596 31894 2648 31900
rect 2504 31884 2556 31890
rect 2504 31826 2556 31832
rect 2516 31482 2544 31826
rect 2504 31476 2556 31482
rect 2504 31418 2556 31424
rect 2424 31300 2544 31328
rect 2412 31204 2464 31210
rect 2412 31146 2464 31152
rect 2318 30288 2374 30297
rect 2318 30223 2374 30232
rect 2320 30184 2372 30190
rect 2320 30126 2372 30132
rect 2332 26926 2360 30126
rect 2424 26926 2452 31146
rect 2516 28014 2544 31300
rect 2608 31210 2636 31894
rect 2688 31680 2740 31686
rect 2688 31622 2740 31628
rect 2700 31414 2728 31622
rect 2688 31408 2740 31414
rect 2688 31350 2740 31356
rect 2976 31346 3004 32388
rect 3054 32328 3110 32337
rect 3054 32263 3056 32272
rect 3108 32263 3110 32272
rect 3056 32234 3108 32240
rect 3056 31748 3108 31754
rect 3056 31690 3108 31696
rect 3068 31482 3096 31690
rect 3056 31476 3108 31482
rect 3056 31418 3108 31424
rect 2964 31340 3016 31346
rect 2964 31282 3016 31288
rect 2596 31204 2648 31210
rect 2596 31146 2648 31152
rect 2582 31036 2890 31056
rect 2582 31034 2588 31036
rect 2644 31034 2668 31036
rect 2724 31034 2748 31036
rect 2804 31034 2828 31036
rect 2884 31034 2890 31036
rect 2644 30982 2646 31034
rect 2826 30982 2828 31034
rect 2582 30980 2588 30982
rect 2644 30980 2668 30982
rect 2724 30980 2748 30982
rect 2804 30980 2828 30982
rect 2884 30980 2890 30982
rect 2582 30960 2890 30980
rect 2780 30592 2832 30598
rect 2778 30560 2780 30569
rect 2832 30560 2834 30569
rect 2778 30495 2834 30504
rect 2976 30190 3004 31282
rect 2964 30184 3016 30190
rect 2964 30126 3016 30132
rect 2582 29948 2890 29968
rect 2582 29946 2588 29948
rect 2644 29946 2668 29948
rect 2724 29946 2748 29948
rect 2804 29946 2828 29948
rect 2884 29946 2890 29948
rect 2644 29894 2646 29946
rect 2826 29894 2828 29946
rect 2582 29892 2588 29894
rect 2644 29892 2668 29894
rect 2724 29892 2748 29894
rect 2804 29892 2828 29894
rect 2884 29892 2890 29894
rect 2582 29872 2890 29892
rect 2778 29608 2834 29617
rect 2778 29543 2780 29552
rect 2832 29543 2834 29552
rect 2780 29514 2832 29520
rect 2976 29345 3004 30126
rect 3056 29504 3108 29510
rect 3056 29446 3108 29452
rect 2962 29336 3018 29345
rect 2962 29271 3018 29280
rect 2964 29164 3016 29170
rect 2964 29106 3016 29112
rect 2582 28860 2890 28880
rect 2582 28858 2588 28860
rect 2644 28858 2668 28860
rect 2724 28858 2748 28860
rect 2804 28858 2828 28860
rect 2884 28858 2890 28860
rect 2644 28806 2646 28858
rect 2826 28806 2828 28858
rect 2582 28804 2588 28806
rect 2644 28804 2668 28806
rect 2724 28804 2748 28806
rect 2804 28804 2828 28806
rect 2884 28804 2890 28806
rect 2582 28784 2890 28804
rect 2872 28688 2924 28694
rect 2976 28665 3004 29106
rect 3068 28694 3096 29446
rect 3160 29306 3188 37839
rect 3252 33658 3280 37998
rect 3528 37856 3556 41103
rect 3344 37828 3556 37856
rect 3344 36802 3372 37828
rect 3514 37768 3570 37777
rect 3514 37703 3516 37712
rect 3568 37703 3570 37712
rect 3516 37674 3568 37680
rect 3424 37664 3476 37670
rect 3424 37606 3476 37612
rect 3436 37369 3464 37606
rect 3422 37360 3478 37369
rect 3422 37295 3478 37304
rect 3344 36774 3556 36802
rect 3422 36680 3478 36689
rect 3422 36615 3424 36624
rect 3476 36615 3478 36624
rect 3424 36586 3476 36592
rect 3332 36576 3384 36582
rect 3332 36518 3384 36524
rect 3422 36544 3478 36553
rect 3240 33652 3292 33658
rect 3240 33594 3292 33600
rect 3240 33516 3292 33522
rect 3240 33458 3292 33464
rect 3148 29300 3200 29306
rect 3148 29242 3200 29248
rect 3148 29164 3200 29170
rect 3148 29106 3200 29112
rect 3056 28688 3108 28694
rect 2872 28630 2924 28636
rect 2962 28656 3018 28665
rect 2504 28008 2556 28014
rect 2504 27950 2556 27956
rect 2320 26920 2372 26926
rect 2320 26862 2372 26868
rect 2412 26920 2464 26926
rect 2412 26862 2464 26868
rect 2332 26314 2360 26862
rect 2320 26308 2372 26314
rect 2320 26250 2372 26256
rect 2320 26036 2372 26042
rect 2320 25978 2372 25984
rect 2332 22273 2360 25978
rect 2318 22264 2374 22273
rect 2318 22199 2374 22208
rect 2320 22160 2372 22166
rect 2320 22102 2372 22108
rect 2228 22092 2280 22098
rect 2228 22034 2280 22040
rect 2226 21992 2282 22001
rect 2226 21927 2282 21936
rect 2240 20466 2268 21927
rect 2332 21554 2360 22102
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 2320 21412 2372 21418
rect 2320 21354 2372 21360
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2240 18193 2268 18702
rect 2226 18184 2282 18193
rect 2226 18119 2282 18128
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2240 17066 2268 17614
rect 2228 17060 2280 17066
rect 2228 17002 2280 17008
rect 2240 15706 2268 17002
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2228 15564 2280 15570
rect 2228 15506 2280 15512
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 2240 15042 2268 15506
rect 2332 15450 2360 21354
rect 2424 21010 2452 26862
rect 2516 26042 2544 27950
rect 2884 27946 2912 28630
rect 3056 28630 3108 28636
rect 2962 28591 3018 28600
rect 3056 28552 3108 28558
rect 3056 28494 3108 28500
rect 2964 28416 3016 28422
rect 2964 28358 3016 28364
rect 2872 27940 2924 27946
rect 2872 27882 2924 27888
rect 2582 27772 2890 27792
rect 2582 27770 2588 27772
rect 2644 27770 2668 27772
rect 2724 27770 2748 27772
rect 2804 27770 2828 27772
rect 2884 27770 2890 27772
rect 2644 27718 2646 27770
rect 2826 27718 2828 27770
rect 2582 27716 2588 27718
rect 2644 27716 2668 27718
rect 2724 27716 2748 27718
rect 2804 27716 2828 27718
rect 2884 27716 2890 27718
rect 2582 27696 2890 27716
rect 2778 27628 2834 27637
rect 2778 27563 2834 27572
rect 2792 26874 2820 27563
rect 2976 27130 3004 28358
rect 3068 27606 3096 28494
rect 3160 28218 3188 29106
rect 3148 28212 3200 28218
rect 3148 28154 3200 28160
rect 3148 27940 3200 27946
rect 3148 27882 3200 27888
rect 3056 27600 3108 27606
rect 3056 27542 3108 27548
rect 2964 27124 3016 27130
rect 2964 27066 3016 27072
rect 3056 26988 3108 26994
rect 3056 26930 3108 26936
rect 2792 26846 3004 26874
rect 2582 26684 2890 26704
rect 2582 26682 2588 26684
rect 2644 26682 2668 26684
rect 2724 26682 2748 26684
rect 2804 26682 2828 26684
rect 2884 26682 2890 26684
rect 2644 26630 2646 26682
rect 2826 26630 2828 26682
rect 2582 26628 2588 26630
rect 2644 26628 2668 26630
rect 2724 26628 2748 26630
rect 2804 26628 2828 26630
rect 2884 26628 2890 26630
rect 2582 26608 2890 26628
rect 2596 26308 2648 26314
rect 2596 26250 2648 26256
rect 2504 26036 2556 26042
rect 2504 25978 2556 25984
rect 2608 25809 2636 26250
rect 2976 25906 3004 26846
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 2594 25800 2650 25809
rect 2594 25735 2650 25744
rect 2582 25596 2890 25616
rect 2582 25594 2588 25596
rect 2644 25594 2668 25596
rect 2724 25594 2748 25596
rect 2804 25594 2828 25596
rect 2884 25594 2890 25596
rect 2644 25542 2646 25594
rect 2826 25542 2828 25594
rect 2582 25540 2588 25542
rect 2644 25540 2668 25542
rect 2724 25540 2748 25542
rect 2804 25540 2828 25542
rect 2884 25540 2890 25542
rect 2582 25520 2890 25540
rect 2976 25294 3004 25842
rect 2964 25288 3016 25294
rect 2964 25230 3016 25236
rect 2504 25220 2556 25226
rect 2504 25162 2556 25168
rect 2516 23118 2544 25162
rect 2778 24848 2834 24857
rect 2778 24783 2780 24792
rect 2832 24783 2834 24792
rect 2780 24754 2832 24760
rect 2964 24744 3016 24750
rect 2964 24686 3016 24692
rect 2582 24508 2890 24528
rect 2582 24506 2588 24508
rect 2644 24506 2668 24508
rect 2724 24506 2748 24508
rect 2804 24506 2828 24508
rect 2884 24506 2890 24508
rect 2644 24454 2646 24506
rect 2826 24454 2828 24506
rect 2582 24452 2588 24454
rect 2644 24452 2668 24454
rect 2724 24452 2748 24454
rect 2804 24452 2828 24454
rect 2884 24452 2890 24454
rect 2582 24432 2890 24452
rect 2872 24336 2924 24342
rect 2872 24278 2924 24284
rect 2884 24018 2912 24278
rect 2976 24177 3004 24686
rect 3068 24342 3096 26930
rect 3160 24750 3188 27882
rect 3148 24744 3200 24750
rect 3148 24686 3200 24692
rect 3148 24608 3200 24614
rect 3148 24550 3200 24556
rect 3056 24336 3108 24342
rect 3056 24278 3108 24284
rect 2962 24168 3018 24177
rect 2962 24103 3018 24112
rect 3056 24132 3108 24138
rect 3056 24074 3108 24080
rect 2884 23990 3004 24018
rect 2780 23656 2832 23662
rect 2778 23624 2780 23633
rect 2832 23624 2834 23633
rect 2778 23559 2834 23568
rect 2582 23420 2890 23440
rect 2582 23418 2588 23420
rect 2644 23418 2668 23420
rect 2724 23418 2748 23420
rect 2804 23418 2828 23420
rect 2884 23418 2890 23420
rect 2644 23366 2646 23418
rect 2826 23366 2828 23418
rect 2582 23364 2588 23366
rect 2644 23364 2668 23366
rect 2724 23364 2748 23366
rect 2804 23364 2828 23366
rect 2884 23364 2890 23366
rect 2582 23344 2890 23364
rect 2976 23118 3004 23990
rect 3068 23322 3096 24074
rect 3056 23316 3108 23322
rect 3056 23258 3108 23264
rect 2504 23112 2556 23118
rect 2504 23054 2556 23060
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 2516 22234 2544 23054
rect 2582 22332 2890 22352
rect 2582 22330 2588 22332
rect 2644 22330 2668 22332
rect 2724 22330 2748 22332
rect 2804 22330 2828 22332
rect 2884 22330 2890 22332
rect 2644 22278 2646 22330
rect 2826 22278 2828 22330
rect 2582 22276 2588 22278
rect 2644 22276 2668 22278
rect 2724 22276 2748 22278
rect 2804 22276 2828 22278
rect 2884 22276 2890 22278
rect 2582 22256 2890 22276
rect 2504 22228 2556 22234
rect 2504 22170 2556 22176
rect 2688 22160 2740 22166
rect 2502 22128 2558 22137
rect 2688 22102 2740 22108
rect 2502 22063 2558 22072
rect 2596 22092 2648 22098
rect 2412 21004 2464 21010
rect 2412 20946 2464 20952
rect 2516 20058 2544 22063
rect 2596 22034 2648 22040
rect 2608 21418 2636 22034
rect 2700 21486 2728 22102
rect 2976 22030 3004 23054
rect 3054 22808 3110 22817
rect 3054 22743 3056 22752
rect 3108 22743 3110 22752
rect 3056 22714 3108 22720
rect 3160 22098 3188 24550
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 2964 22024 3016 22030
rect 2964 21966 3016 21972
rect 2976 21554 3004 21966
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 2688 21480 2740 21486
rect 2688 21422 2740 21428
rect 2976 21418 3004 21490
rect 2596 21412 2648 21418
rect 2596 21354 2648 21360
rect 2964 21412 3016 21418
rect 2964 21354 3016 21360
rect 2582 21244 2890 21264
rect 2582 21242 2588 21244
rect 2644 21242 2668 21244
rect 2724 21242 2748 21244
rect 2804 21242 2828 21244
rect 2884 21242 2890 21244
rect 2644 21190 2646 21242
rect 2826 21190 2828 21242
rect 2582 21188 2588 21190
rect 2644 21188 2668 21190
rect 2724 21188 2748 21190
rect 2804 21188 2828 21190
rect 2884 21188 2890 21190
rect 2582 21168 2890 21188
rect 2976 20942 3004 21354
rect 2964 20936 3016 20942
rect 2964 20878 3016 20884
rect 2582 20156 2890 20176
rect 2582 20154 2588 20156
rect 2644 20154 2668 20156
rect 2724 20154 2748 20156
rect 2804 20154 2828 20156
rect 2884 20154 2890 20156
rect 2644 20102 2646 20154
rect 2826 20102 2828 20154
rect 2582 20100 2588 20102
rect 2644 20100 2668 20102
rect 2724 20100 2748 20102
rect 2804 20100 2828 20102
rect 2884 20100 2890 20102
rect 2582 20080 2890 20100
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 2412 19984 2464 19990
rect 2412 19926 2464 19932
rect 2424 19514 2452 19926
rect 2976 19922 3004 20878
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 2884 19417 2912 19790
rect 2870 19408 2926 19417
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2780 19372 2832 19378
rect 2870 19343 2926 19352
rect 3148 19372 3200 19378
rect 2780 19314 2832 19320
rect 3148 19314 3200 19320
rect 2424 18358 2452 19314
rect 2792 19281 2820 19314
rect 2778 19272 2834 19281
rect 2778 19207 2834 19216
rect 2582 19068 2890 19088
rect 2582 19066 2588 19068
rect 2644 19066 2668 19068
rect 2724 19066 2748 19068
rect 2804 19066 2828 19068
rect 2884 19066 2890 19068
rect 2644 19014 2646 19066
rect 2826 19014 2828 19066
rect 2582 19012 2588 19014
rect 2644 19012 2668 19014
rect 2724 19012 2748 19014
rect 2804 19012 2828 19014
rect 2884 19012 2890 19014
rect 2582 18992 2890 19012
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2884 18601 2912 18702
rect 2870 18592 2926 18601
rect 2870 18527 2926 18536
rect 2412 18352 2464 18358
rect 2412 18294 2464 18300
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2582 17980 2890 18000
rect 2582 17978 2588 17980
rect 2644 17978 2668 17980
rect 2724 17978 2748 17980
rect 2804 17978 2828 17980
rect 2884 17978 2890 17980
rect 2644 17926 2646 17978
rect 2826 17926 2828 17978
rect 2582 17924 2588 17926
rect 2644 17924 2668 17926
rect 2724 17924 2748 17926
rect 2804 17924 2828 17926
rect 2884 17924 2890 17926
rect 2582 17904 2890 17924
rect 2976 17762 3004 18022
rect 2792 17734 3004 17762
rect 2792 17678 2820 17734
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2792 17066 2820 17614
rect 2976 17270 3004 17614
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 3068 17338 3096 17546
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2582 16892 2890 16912
rect 2582 16890 2588 16892
rect 2644 16890 2668 16892
rect 2724 16890 2748 16892
rect 2804 16890 2828 16892
rect 2884 16890 2890 16892
rect 2644 16838 2646 16890
rect 2826 16838 2828 16890
rect 2582 16836 2588 16838
rect 2644 16836 2668 16838
rect 2724 16836 2748 16838
rect 2804 16836 2828 16838
rect 2884 16836 2890 16838
rect 2582 16816 2890 16836
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2516 15978 2544 16390
rect 2792 16017 2820 16526
rect 2884 16250 2912 16594
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2778 16008 2834 16017
rect 2504 15972 2556 15978
rect 2778 15943 2834 15952
rect 2504 15914 2556 15920
rect 2582 15804 2890 15824
rect 2582 15802 2588 15804
rect 2644 15802 2668 15804
rect 2724 15802 2748 15804
rect 2804 15802 2828 15804
rect 2884 15802 2890 15804
rect 2644 15750 2646 15802
rect 2826 15750 2828 15802
rect 2582 15748 2588 15750
rect 2644 15748 2668 15750
rect 2724 15748 2748 15750
rect 2804 15748 2828 15750
rect 2884 15748 2890 15750
rect 2582 15728 2890 15748
rect 2872 15496 2924 15502
rect 2332 15422 2544 15450
rect 2872 15438 2924 15444
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2148 15014 2268 15042
rect 2148 14346 2176 15014
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 2042 13152 2098 13161
rect 2042 13087 2098 13096
rect 1964 12838 2084 12866
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1964 7954 1992 12718
rect 2056 11354 2084 12838
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1504 6854 1624 6882
rect 1504 5778 1532 6854
rect 1676 6792 1728 6798
rect 1582 6760 1638 6769
rect 1676 6734 1728 6740
rect 1582 6695 1638 6704
rect 1596 6662 1624 6695
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1400 5704 1452 5710
rect 1306 5672 1362 5681
rect 1400 5646 1452 5652
rect 1306 5607 1362 5616
rect 1320 5234 1348 5607
rect 1412 5273 1440 5646
rect 1398 5264 1454 5273
rect 1308 5228 1360 5234
rect 1398 5199 1454 5208
rect 1308 5170 1360 5176
rect 1400 4072 1452 4078
rect 1398 4040 1400 4049
rect 1452 4040 1454 4049
rect 1398 3975 1454 3984
rect 1688 2922 1716 6734
rect 2056 6390 2084 11154
rect 2148 10130 2176 14282
rect 2240 13938 2268 14758
rect 2332 14482 2360 15302
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2424 14074 2452 14962
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2228 13932 2280 13938
rect 2280 13892 2360 13920
rect 2228 13874 2280 13880
rect 2332 13394 2360 13892
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2424 12714 2452 13466
rect 2516 13326 2544 15422
rect 2884 14929 2912 15438
rect 2870 14920 2926 14929
rect 2870 14855 2926 14864
rect 2582 14716 2890 14736
rect 2582 14714 2588 14716
rect 2644 14714 2668 14716
rect 2724 14714 2748 14716
rect 2804 14714 2828 14716
rect 2884 14714 2890 14716
rect 2644 14662 2646 14714
rect 2826 14662 2828 14714
rect 2582 14660 2588 14662
rect 2644 14660 2668 14662
rect 2724 14660 2748 14662
rect 2804 14660 2828 14662
rect 2884 14660 2890 14662
rect 2582 14640 2890 14660
rect 2976 14618 3004 17206
rect 3160 15178 3188 19314
rect 3068 15150 3188 15178
rect 3068 14906 3096 15150
rect 3148 15088 3200 15094
rect 3146 15056 3148 15065
rect 3200 15056 3202 15065
rect 3146 14991 3202 15000
rect 3068 14878 3188 14906
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2688 14272 2740 14278
rect 2884 14260 2912 14486
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 2740 14232 2912 14260
rect 2688 14214 2740 14220
rect 2582 13628 2890 13648
rect 2582 13626 2588 13628
rect 2644 13626 2668 13628
rect 2724 13626 2748 13628
rect 2804 13626 2828 13628
rect 2884 13626 2890 13628
rect 2644 13574 2646 13626
rect 2826 13574 2828 13626
rect 2582 13572 2588 13574
rect 2644 13572 2668 13574
rect 2724 13572 2748 13574
rect 2804 13572 2828 13574
rect 2884 13572 2890 13574
rect 2582 13552 2890 13572
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2412 12708 2464 12714
rect 2412 12650 2464 12656
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2240 12442 2268 12582
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2240 11558 2268 12378
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2240 7562 2268 11290
rect 2148 7534 2268 7562
rect 2044 6384 2096 6390
rect 2044 6326 2096 6332
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1872 6225 1900 6258
rect 1858 6216 1914 6225
rect 1858 6151 1914 6160
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1780 4078 1808 4558
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1964 3534 1992 4558
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 2148 3194 2176 7534
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2240 7041 2268 7346
rect 2226 7032 2282 7041
rect 2226 6967 2282 6976
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2240 6633 2268 6666
rect 2226 6624 2282 6633
rect 2226 6559 2282 6568
rect 2332 5914 2360 11562
rect 2424 9042 2452 12650
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2424 5166 2452 8366
rect 2516 7478 2544 13262
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2608 12714 2636 12786
rect 2884 12714 2912 13330
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2596 12708 2648 12714
rect 2596 12650 2648 12656
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2582 12540 2890 12560
rect 2582 12538 2588 12540
rect 2644 12538 2668 12540
rect 2724 12538 2748 12540
rect 2804 12538 2828 12540
rect 2884 12538 2890 12540
rect 2644 12486 2646 12538
rect 2826 12486 2828 12538
rect 2582 12484 2588 12486
rect 2644 12484 2668 12486
rect 2724 12484 2748 12486
rect 2804 12484 2828 12486
rect 2884 12484 2890 12486
rect 2582 12464 2890 12484
rect 2976 12374 3004 13126
rect 3068 12986 3096 14282
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2582 11452 2890 11472
rect 2582 11450 2588 11452
rect 2644 11450 2668 11452
rect 2724 11450 2748 11452
rect 2804 11450 2828 11452
rect 2884 11450 2890 11452
rect 2644 11398 2646 11450
rect 2826 11398 2828 11450
rect 2582 11396 2588 11398
rect 2644 11396 2668 11398
rect 2724 11396 2748 11398
rect 2804 11396 2828 11398
rect 2884 11396 2890 11398
rect 2582 11376 2890 11396
rect 2582 10364 2890 10384
rect 2582 10362 2588 10364
rect 2644 10362 2668 10364
rect 2724 10362 2748 10364
rect 2804 10362 2828 10364
rect 2884 10362 2890 10364
rect 2644 10310 2646 10362
rect 2826 10310 2828 10362
rect 2582 10308 2588 10310
rect 2644 10308 2668 10310
rect 2724 10308 2748 10310
rect 2804 10308 2828 10310
rect 2884 10308 2890 10310
rect 2582 10288 2890 10308
rect 3068 10062 3096 12650
rect 3160 11898 3188 14878
rect 3252 13938 3280 33458
rect 3344 30938 3372 36518
rect 3422 36479 3478 36488
rect 3436 32230 3464 36479
rect 3528 35766 3556 36774
rect 3516 35760 3568 35766
rect 3516 35702 3568 35708
rect 3424 32224 3476 32230
rect 3424 32166 3476 32172
rect 3422 32056 3478 32065
rect 3422 31991 3478 32000
rect 3332 30932 3384 30938
rect 3332 30874 3384 30880
rect 3330 30832 3386 30841
rect 3330 30767 3386 30776
rect 3344 30122 3372 30767
rect 3332 30116 3384 30122
rect 3332 30058 3384 30064
rect 3332 28484 3384 28490
rect 3332 28426 3384 28432
rect 3344 28393 3372 28426
rect 3330 28384 3386 28393
rect 3330 28319 3386 28328
rect 3332 28212 3384 28218
rect 3332 28154 3384 28160
rect 3344 26518 3372 28154
rect 3332 26512 3384 26518
rect 3332 26454 3384 26460
rect 3332 26308 3384 26314
rect 3332 26250 3384 26256
rect 3344 25498 3372 26250
rect 3332 25492 3384 25498
rect 3332 25434 3384 25440
rect 3436 24818 3464 31991
rect 3528 26330 3556 35702
rect 3620 28218 3648 41239
rect 3712 37262 3740 46158
rect 3792 45960 3844 45966
rect 3988 45914 4016 46532
rect 3792 45902 3844 45908
rect 3804 45665 3832 45902
rect 3896 45886 4016 45914
rect 3790 45656 3846 45665
rect 3790 45591 3846 45600
rect 3792 45552 3844 45558
rect 3792 45494 3844 45500
rect 3804 44402 3832 45494
rect 3896 44742 3924 45886
rect 3976 45824 4028 45830
rect 3976 45766 4028 45772
rect 3988 45529 4016 45766
rect 3974 45520 4030 45529
rect 3974 45455 4030 45464
rect 3976 44804 4028 44810
rect 3976 44746 4028 44752
rect 3884 44736 3936 44742
rect 3884 44678 3936 44684
rect 3792 44396 3844 44402
rect 3792 44338 3844 44344
rect 3988 44334 4016 44746
rect 3884 44328 3936 44334
rect 3884 44270 3936 44276
rect 3976 44328 4028 44334
rect 3976 44270 4028 44276
rect 3792 44192 3844 44198
rect 3792 44134 3844 44140
rect 3804 43353 3832 44134
rect 3896 43897 3924 44270
rect 3882 43888 3938 43897
rect 3882 43823 3938 43832
rect 3884 43784 3936 43790
rect 3884 43726 3936 43732
rect 3790 43344 3846 43353
rect 3790 43279 3846 43288
rect 3792 43172 3844 43178
rect 3792 43114 3844 43120
rect 3804 42945 3832 43114
rect 3790 42936 3846 42945
rect 3790 42871 3846 42880
rect 3790 42800 3846 42809
rect 3790 42735 3846 42744
rect 3804 42702 3832 42735
rect 3792 42696 3844 42702
rect 3792 42638 3844 42644
rect 3790 42120 3846 42129
rect 3790 42055 3792 42064
rect 3844 42055 3846 42064
rect 3792 42026 3844 42032
rect 3790 41984 3846 41993
rect 3790 41919 3846 41928
rect 3804 41546 3832 41919
rect 3792 41540 3844 41546
rect 3792 41482 3844 41488
rect 3790 41440 3846 41449
rect 3790 41375 3846 41384
rect 3804 40730 3832 41375
rect 3896 41313 3924 43726
rect 3988 43217 4016 44270
rect 3974 43208 4030 43217
rect 3974 43143 4030 43152
rect 3976 43104 4028 43110
rect 3976 43046 4028 43052
rect 3988 42537 4016 43046
rect 3974 42528 4030 42537
rect 3974 42463 4030 42472
rect 3976 42220 4028 42226
rect 3976 42162 4028 42168
rect 3882 41304 3938 41313
rect 3882 41239 3938 41248
rect 3884 41200 3936 41206
rect 3884 41142 3936 41148
rect 3792 40724 3844 40730
rect 3792 40666 3844 40672
rect 3896 39624 3924 41142
rect 3988 40662 4016 42162
rect 4080 41614 4108 50798
rect 4172 50454 4200 50866
rect 4618 50824 4674 50833
rect 4618 50759 4674 50768
rect 4160 50448 4212 50454
rect 4160 50390 4212 50396
rect 4214 50076 4522 50096
rect 4214 50074 4220 50076
rect 4276 50074 4300 50076
rect 4356 50074 4380 50076
rect 4436 50074 4460 50076
rect 4516 50074 4522 50076
rect 4276 50022 4278 50074
rect 4458 50022 4460 50074
rect 4214 50020 4220 50022
rect 4276 50020 4300 50022
rect 4356 50020 4380 50022
rect 4436 50020 4460 50022
rect 4516 50020 4522 50022
rect 4214 50000 4522 50020
rect 4528 49360 4580 49366
rect 4526 49328 4528 49337
rect 4580 49328 4582 49337
rect 4526 49263 4582 49272
rect 4214 48988 4522 49008
rect 4214 48986 4220 48988
rect 4276 48986 4300 48988
rect 4356 48986 4380 48988
rect 4436 48986 4460 48988
rect 4516 48986 4522 48988
rect 4276 48934 4278 48986
rect 4458 48934 4460 48986
rect 4214 48932 4220 48934
rect 4276 48932 4300 48934
rect 4356 48932 4380 48934
rect 4436 48932 4460 48934
rect 4516 48932 4522 48934
rect 4214 48912 4522 48932
rect 4526 48512 4582 48521
rect 4526 48447 4582 48456
rect 4540 48346 4568 48447
rect 4528 48340 4580 48346
rect 4528 48282 4580 48288
rect 4526 48104 4582 48113
rect 4526 48039 4528 48048
rect 4580 48039 4582 48048
rect 4528 48010 4580 48016
rect 4214 47900 4522 47920
rect 4214 47898 4220 47900
rect 4276 47898 4300 47900
rect 4356 47898 4380 47900
rect 4436 47898 4460 47900
rect 4516 47898 4522 47900
rect 4276 47846 4278 47898
rect 4458 47846 4460 47898
rect 4214 47844 4220 47846
rect 4276 47844 4300 47846
rect 4356 47844 4380 47846
rect 4436 47844 4460 47846
rect 4516 47844 4522 47846
rect 4214 47824 4522 47844
rect 4632 47569 4660 50759
rect 4618 47560 4674 47569
rect 4618 47495 4674 47504
rect 4620 47184 4672 47190
rect 4620 47126 4672 47132
rect 4528 47048 4580 47054
rect 4526 47016 4528 47025
rect 4580 47016 4582 47025
rect 4526 46951 4582 46960
rect 4214 46812 4522 46832
rect 4214 46810 4220 46812
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4516 46810 4522 46812
rect 4276 46758 4278 46810
rect 4458 46758 4460 46810
rect 4214 46756 4220 46758
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4516 46756 4522 46758
rect 4214 46736 4522 46756
rect 4160 46504 4212 46510
rect 4160 46446 4212 46452
rect 4172 45898 4200 46446
rect 4632 46322 4660 47126
rect 4540 46294 4660 46322
rect 4540 46102 4568 46294
rect 4724 46186 4752 50918
rect 4804 50924 4856 50930
rect 4804 50866 4856 50872
rect 4802 50688 4858 50697
rect 4802 50623 4858 50632
rect 4632 46158 4752 46186
rect 4528 46096 4580 46102
rect 4528 46038 4580 46044
rect 4160 45892 4212 45898
rect 4160 45834 4212 45840
rect 4214 45724 4522 45744
rect 4214 45722 4220 45724
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4516 45722 4522 45724
rect 4276 45670 4278 45722
rect 4458 45670 4460 45722
rect 4214 45668 4220 45670
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4516 45668 4522 45670
rect 4214 45648 4522 45668
rect 4214 44636 4522 44656
rect 4214 44634 4220 44636
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4516 44634 4522 44636
rect 4276 44582 4278 44634
rect 4458 44582 4460 44634
rect 4214 44580 4220 44582
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4516 44580 4522 44582
rect 4214 44560 4522 44580
rect 4252 44396 4304 44402
rect 4252 44338 4304 44344
rect 4264 43790 4292 44338
rect 4252 43784 4304 43790
rect 4252 43726 4304 43732
rect 4214 43548 4522 43568
rect 4214 43546 4220 43548
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4516 43546 4522 43548
rect 4276 43494 4278 43546
rect 4458 43494 4460 43546
rect 4214 43492 4220 43494
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4516 43492 4522 43494
rect 4214 43472 4522 43492
rect 4158 43344 4214 43353
rect 4158 43279 4214 43288
rect 4172 43246 4200 43279
rect 4160 43240 4212 43246
rect 4160 43182 4212 43188
rect 4214 42460 4522 42480
rect 4214 42458 4220 42460
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4516 42458 4522 42460
rect 4276 42406 4278 42458
rect 4458 42406 4460 42458
rect 4214 42404 4220 42406
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4516 42404 4522 42406
rect 4214 42384 4522 42404
rect 4436 42288 4488 42294
rect 4436 42230 4488 42236
rect 4160 41676 4212 41682
rect 4160 41618 4212 41624
rect 4068 41608 4120 41614
rect 4068 41550 4120 41556
rect 4172 41460 4200 41618
rect 4448 41614 4476 42230
rect 4436 41608 4488 41614
rect 4436 41550 4488 41556
rect 4080 41432 4200 41460
rect 4080 41002 4108 41432
rect 4214 41372 4522 41392
rect 4214 41370 4220 41372
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4516 41370 4522 41372
rect 4276 41318 4278 41370
rect 4458 41318 4460 41370
rect 4214 41316 4220 41318
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4516 41316 4522 41318
rect 4214 41296 4522 41316
rect 4344 41200 4396 41206
rect 4344 41142 4396 41148
rect 4068 40996 4120 41002
rect 4068 40938 4120 40944
rect 4068 40724 4120 40730
rect 4068 40666 4120 40672
rect 3976 40656 4028 40662
rect 3976 40598 4028 40604
rect 3976 40384 4028 40390
rect 3976 40326 4028 40332
rect 3988 39817 4016 40326
rect 3974 39808 4030 39817
rect 3974 39743 4030 39752
rect 3896 39596 4016 39624
rect 3792 39568 3844 39574
rect 3792 39510 3844 39516
rect 3804 39137 3832 39510
rect 3882 39400 3938 39409
rect 3882 39335 3938 39344
rect 3790 39128 3846 39137
rect 3790 39063 3846 39072
rect 3792 39024 3844 39030
rect 3792 38966 3844 38972
rect 3804 37874 3832 38966
rect 3896 38457 3924 39335
rect 3882 38448 3938 38457
rect 3882 38383 3938 38392
rect 3988 38298 4016 39596
rect 3896 38270 4016 38298
rect 3792 37868 3844 37874
rect 3792 37810 3844 37816
rect 3790 37768 3846 37777
rect 3790 37703 3846 37712
rect 3700 37256 3752 37262
rect 3700 37198 3752 37204
rect 3700 37120 3752 37126
rect 3700 37062 3752 37068
rect 3712 35193 3740 37062
rect 3804 35698 3832 37703
rect 3792 35692 3844 35698
rect 3792 35634 3844 35640
rect 3790 35320 3846 35329
rect 3790 35255 3846 35264
rect 3698 35184 3754 35193
rect 3698 35119 3754 35128
rect 3700 35080 3752 35086
rect 3700 35022 3752 35028
rect 3712 32366 3740 35022
rect 3804 33930 3832 35255
rect 3792 33924 3844 33930
rect 3792 33866 3844 33872
rect 3790 33824 3846 33833
rect 3790 33759 3846 33768
rect 3804 33522 3832 33759
rect 3792 33516 3844 33522
rect 3792 33458 3844 33464
rect 3792 32904 3844 32910
rect 3792 32846 3844 32852
rect 3700 32360 3752 32366
rect 3700 32302 3752 32308
rect 3700 32224 3752 32230
rect 3700 32166 3752 32172
rect 3608 28212 3660 28218
rect 3608 28154 3660 28160
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3620 27169 3648 28018
rect 3606 27160 3662 27169
rect 3712 27130 3740 32166
rect 3804 30394 3832 32846
rect 3896 32502 3924 38270
rect 3976 35148 4028 35154
rect 3976 35090 4028 35096
rect 3988 34678 4016 35090
rect 3976 34672 4028 34678
rect 3976 34614 4028 34620
rect 3976 34536 4028 34542
rect 3976 34478 4028 34484
rect 3988 33862 4016 34478
rect 3976 33856 4028 33862
rect 3976 33798 4028 33804
rect 3884 32496 3936 32502
rect 3884 32438 3936 32444
rect 3988 32065 4016 33798
rect 3974 32056 4030 32065
rect 3974 31991 4030 32000
rect 3976 31952 4028 31958
rect 3976 31894 4028 31900
rect 3988 31793 4016 31894
rect 3974 31784 4030 31793
rect 3974 31719 4030 31728
rect 3884 31272 3936 31278
rect 3884 31214 3936 31220
rect 3792 30388 3844 30394
rect 3792 30330 3844 30336
rect 3792 30252 3844 30258
rect 3792 30194 3844 30200
rect 3606 27095 3662 27104
rect 3700 27124 3752 27130
rect 3700 27066 3752 27072
rect 3608 26988 3660 26994
rect 3608 26930 3660 26936
rect 3620 26489 3648 26930
rect 3606 26480 3662 26489
rect 3606 26415 3662 26424
rect 3528 26302 3648 26330
rect 3804 26314 3832 30194
rect 3896 28404 3924 31214
rect 4080 28694 4108 40666
rect 4356 40526 4384 41142
rect 4528 41132 4580 41138
rect 4528 41074 4580 41080
rect 4344 40520 4396 40526
rect 4344 40462 4396 40468
rect 4540 40458 4568 41074
rect 4528 40452 4580 40458
rect 4528 40394 4580 40400
rect 4214 40284 4522 40304
rect 4214 40282 4220 40284
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4516 40282 4522 40284
rect 4276 40230 4278 40282
rect 4458 40230 4460 40282
rect 4214 40228 4220 40230
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4516 40228 4522 40230
rect 4214 40208 4522 40228
rect 4344 40112 4396 40118
rect 4344 40054 4396 40060
rect 4526 40080 4582 40089
rect 4252 39840 4304 39846
rect 4252 39782 4304 39788
rect 4264 39409 4292 39782
rect 4356 39438 4384 40054
rect 4526 40015 4582 40024
rect 4344 39432 4396 39438
rect 4250 39400 4306 39409
rect 4344 39374 4396 39380
rect 4250 39335 4306 39344
rect 4540 39284 4568 40015
rect 4632 39438 4660 46158
rect 4712 46096 4764 46102
rect 4712 46038 4764 46044
rect 4724 40662 4752 46038
rect 4712 40656 4764 40662
rect 4712 40598 4764 40604
rect 4712 40452 4764 40458
rect 4712 40394 4764 40400
rect 4724 40118 4752 40394
rect 4712 40112 4764 40118
rect 4712 40054 4764 40060
rect 4710 39944 4766 39953
rect 4710 39879 4766 39888
rect 4620 39432 4672 39438
rect 4620 39374 4672 39380
rect 4540 39256 4660 39284
rect 4214 39196 4522 39216
rect 4214 39194 4220 39196
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4516 39194 4522 39196
rect 4276 39142 4278 39194
rect 4458 39142 4460 39194
rect 4214 39140 4220 39142
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4516 39140 4522 39142
rect 4214 39120 4522 39140
rect 4342 38992 4398 39001
rect 4342 38927 4398 38936
rect 4436 38956 4488 38962
rect 4160 38888 4212 38894
rect 4160 38830 4212 38836
rect 4172 38282 4200 38830
rect 4252 38820 4304 38826
rect 4252 38762 4304 38768
rect 4264 38486 4292 38762
rect 4252 38480 4304 38486
rect 4252 38422 4304 38428
rect 4356 38321 4384 38927
rect 4436 38898 4488 38904
rect 4448 38350 4476 38898
rect 4436 38344 4488 38350
rect 4342 38312 4398 38321
rect 4160 38276 4212 38282
rect 4436 38286 4488 38292
rect 4342 38247 4398 38256
rect 4160 38218 4212 38224
rect 4214 38108 4522 38128
rect 4214 38106 4220 38108
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4516 38106 4522 38108
rect 4276 38054 4278 38106
rect 4458 38054 4460 38106
rect 4214 38052 4220 38054
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4516 38052 4522 38054
rect 4214 38032 4522 38052
rect 4214 37020 4522 37040
rect 4214 37018 4220 37020
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4516 37018 4522 37020
rect 4276 36966 4278 37018
rect 4458 36966 4460 37018
rect 4214 36964 4220 36966
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4516 36964 4522 36966
rect 4214 36944 4522 36964
rect 4528 36848 4580 36854
rect 4526 36816 4528 36825
rect 4580 36816 4582 36825
rect 4526 36751 4582 36760
rect 4214 35932 4522 35952
rect 4214 35930 4220 35932
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4516 35930 4522 35932
rect 4276 35878 4278 35930
rect 4458 35878 4460 35930
rect 4214 35876 4220 35878
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4516 35876 4522 35878
rect 4214 35856 4522 35876
rect 4436 35760 4488 35766
rect 4632 35737 4660 39256
rect 4436 35702 4488 35708
rect 4618 35728 4674 35737
rect 4448 35154 4476 35702
rect 4618 35663 4674 35672
rect 4620 35624 4672 35630
rect 4620 35566 4672 35572
rect 4632 35222 4660 35566
rect 4620 35216 4672 35222
rect 4620 35158 4672 35164
rect 4436 35148 4488 35154
rect 4436 35090 4488 35096
rect 4214 34844 4522 34864
rect 4214 34842 4220 34844
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4516 34842 4522 34844
rect 4276 34790 4278 34842
rect 4458 34790 4460 34842
rect 4214 34788 4220 34790
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4516 34788 4522 34790
rect 4214 34768 4522 34788
rect 4160 34604 4212 34610
rect 4160 34546 4212 34552
rect 4172 33969 4200 34546
rect 4158 33960 4214 33969
rect 4158 33895 4214 33904
rect 4214 33756 4522 33776
rect 4214 33754 4220 33756
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4516 33754 4522 33756
rect 4276 33702 4278 33754
rect 4458 33702 4460 33754
rect 4214 33700 4220 33702
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4516 33700 4522 33702
rect 4214 33680 4522 33700
rect 4214 32668 4522 32688
rect 4214 32666 4220 32668
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4516 32666 4522 32668
rect 4276 32614 4278 32666
rect 4458 32614 4460 32666
rect 4214 32612 4220 32614
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4516 32612 4522 32614
rect 4214 32592 4522 32612
rect 4250 32464 4306 32473
rect 4250 32399 4306 32408
rect 4264 32026 4292 32399
rect 4724 32314 4752 39879
rect 4816 36009 4844 50623
rect 4908 46186 4936 65078
rect 5000 56166 5028 65962
rect 5080 59560 5132 59566
rect 5080 59502 5132 59508
rect 5092 58993 5120 59502
rect 5078 58984 5134 58993
rect 5078 58919 5134 58928
rect 5080 58540 5132 58546
rect 5080 58482 5132 58488
rect 4988 56160 5040 56166
rect 4988 56102 5040 56108
rect 4988 55888 5040 55894
rect 4988 55830 5040 55836
rect 5000 50969 5028 55830
rect 5092 51066 5120 58482
rect 5184 51066 5212 66710
rect 5080 51060 5132 51066
rect 5080 51002 5132 51008
rect 5172 51060 5224 51066
rect 5172 51002 5224 51008
rect 4986 50960 5042 50969
rect 4986 50895 5042 50904
rect 4988 50856 5040 50862
rect 4988 50798 5040 50804
rect 5172 50856 5224 50862
rect 5172 50798 5224 50804
rect 5000 46374 5028 50798
rect 5078 50688 5134 50697
rect 5078 50623 5134 50632
rect 4988 46368 5040 46374
rect 4988 46310 5040 46316
rect 4908 46158 5028 46186
rect 4896 44872 4948 44878
rect 4896 44814 4948 44820
rect 4908 44538 4936 44814
rect 4896 44532 4948 44538
rect 4896 44474 4948 44480
rect 4896 44396 4948 44402
rect 4896 44338 4948 44344
rect 4908 42294 4936 44338
rect 4896 42288 4948 42294
rect 4896 42230 4948 42236
rect 4894 42120 4950 42129
rect 4894 42055 4950 42064
rect 4802 36000 4858 36009
rect 4802 35935 4858 35944
rect 4908 35816 4936 42055
rect 5000 41857 5028 46158
rect 4986 41848 5042 41857
rect 4986 41783 5042 41792
rect 5092 41698 5120 50623
rect 5184 47190 5212 50798
rect 5172 47184 5224 47190
rect 5172 47126 5224 47132
rect 5172 46912 5224 46918
rect 5172 46854 5224 46860
rect 5184 44266 5212 46854
rect 5172 44260 5224 44266
rect 5172 44202 5224 44208
rect 5276 42226 5304 75958
rect 5846 75644 6154 75664
rect 5846 75642 5852 75644
rect 5908 75642 5932 75644
rect 5988 75642 6012 75644
rect 6068 75642 6092 75644
rect 6148 75642 6154 75644
rect 5908 75590 5910 75642
rect 6090 75590 6092 75642
rect 5846 75588 5852 75590
rect 5908 75588 5932 75590
rect 5988 75588 6012 75590
rect 6068 75588 6092 75590
rect 6148 75588 6154 75590
rect 5846 75568 6154 75588
rect 7478 75100 7786 75120
rect 7478 75098 7484 75100
rect 7540 75098 7564 75100
rect 7620 75098 7644 75100
rect 7700 75098 7724 75100
rect 7780 75098 7786 75100
rect 7540 75046 7542 75098
rect 7722 75046 7724 75098
rect 7478 75044 7484 75046
rect 7540 75044 7564 75046
rect 7620 75044 7644 75046
rect 7700 75044 7724 75046
rect 7780 75044 7786 75046
rect 7478 75024 7786 75044
rect 5846 74556 6154 74576
rect 5846 74554 5852 74556
rect 5908 74554 5932 74556
rect 5988 74554 6012 74556
rect 6068 74554 6092 74556
rect 6148 74554 6154 74556
rect 5908 74502 5910 74554
rect 6090 74502 6092 74554
rect 5846 74500 5852 74502
rect 5908 74500 5932 74502
rect 5988 74500 6012 74502
rect 6068 74500 6092 74502
rect 6148 74500 6154 74502
rect 5846 74480 6154 74500
rect 7478 74012 7786 74032
rect 7478 74010 7484 74012
rect 7540 74010 7564 74012
rect 7620 74010 7644 74012
rect 7700 74010 7724 74012
rect 7780 74010 7786 74012
rect 7540 73958 7542 74010
rect 7722 73958 7724 74010
rect 7478 73956 7484 73958
rect 7540 73956 7564 73958
rect 7620 73956 7644 73958
rect 7700 73956 7724 73958
rect 7780 73956 7786 73958
rect 7478 73936 7786 73956
rect 5846 73468 6154 73488
rect 5846 73466 5852 73468
rect 5908 73466 5932 73468
rect 5988 73466 6012 73468
rect 6068 73466 6092 73468
rect 6148 73466 6154 73468
rect 5908 73414 5910 73466
rect 6090 73414 6092 73466
rect 5846 73412 5852 73414
rect 5908 73412 5932 73414
rect 5988 73412 6012 73414
rect 6068 73412 6092 73414
rect 6148 73412 6154 73414
rect 5846 73392 6154 73412
rect 7478 72924 7786 72944
rect 7478 72922 7484 72924
rect 7540 72922 7564 72924
rect 7620 72922 7644 72924
rect 7700 72922 7724 72924
rect 7780 72922 7786 72924
rect 7540 72870 7542 72922
rect 7722 72870 7724 72922
rect 7478 72868 7484 72870
rect 7540 72868 7564 72870
rect 7620 72868 7644 72870
rect 7700 72868 7724 72870
rect 7780 72868 7786 72870
rect 7478 72848 7786 72868
rect 5540 72548 5592 72554
rect 5540 72490 5592 72496
rect 5448 67040 5500 67046
rect 5448 66982 5500 66988
rect 5460 66201 5488 66982
rect 5446 66192 5502 66201
rect 5446 66127 5502 66136
rect 5356 62416 5408 62422
rect 5356 62358 5408 62364
rect 5368 55894 5396 62358
rect 5448 56160 5500 56166
rect 5448 56102 5500 56108
rect 5356 55888 5408 55894
rect 5356 55830 5408 55836
rect 5356 53508 5408 53514
rect 5356 53450 5408 53456
rect 5368 52737 5396 53450
rect 5354 52728 5410 52737
rect 5354 52663 5410 52672
rect 5356 52556 5408 52562
rect 5356 52498 5408 52504
rect 5368 52193 5396 52498
rect 5354 52184 5410 52193
rect 5354 52119 5410 52128
rect 5356 52012 5408 52018
rect 5356 51954 5408 51960
rect 5368 51097 5396 51954
rect 5354 51088 5410 51097
rect 5354 51023 5410 51032
rect 5460 50946 5488 56102
rect 5368 50930 5488 50946
rect 5356 50924 5488 50930
rect 5408 50918 5488 50924
rect 5356 50866 5408 50872
rect 5448 50856 5500 50862
rect 5354 50824 5410 50833
rect 5448 50798 5500 50804
rect 5354 50759 5410 50768
rect 5264 42220 5316 42226
rect 5264 42162 5316 42168
rect 5000 41670 5120 41698
rect 5264 41676 5316 41682
rect 5000 40633 5028 41670
rect 5264 41618 5316 41624
rect 5080 41608 5132 41614
rect 5080 41550 5132 41556
rect 5092 41070 5120 41550
rect 5276 41313 5304 41618
rect 5262 41304 5318 41313
rect 5262 41239 5318 41248
rect 5368 41188 5396 50759
rect 5184 41160 5396 41188
rect 5080 41064 5132 41070
rect 5080 41006 5132 41012
rect 5080 40928 5132 40934
rect 5080 40870 5132 40876
rect 4986 40624 5042 40633
rect 4986 40559 5042 40568
rect 4988 40520 5040 40526
rect 4988 40462 5040 40468
rect 5000 36922 5028 40462
rect 4988 36916 5040 36922
rect 4988 36858 5040 36864
rect 4540 32286 4752 32314
rect 4816 35788 4936 35816
rect 4252 32020 4304 32026
rect 4252 31962 4304 31968
rect 4540 31793 4568 32286
rect 4712 32224 4764 32230
rect 4712 32166 4764 32172
rect 4620 31884 4672 31890
rect 4620 31826 4672 31832
rect 4526 31784 4582 31793
rect 4526 31719 4582 31728
rect 4214 31580 4522 31600
rect 4214 31578 4220 31580
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4516 31578 4522 31580
rect 4276 31526 4278 31578
rect 4458 31526 4460 31578
rect 4214 31524 4220 31526
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4516 31524 4522 31526
rect 4214 31504 4522 31524
rect 4526 31376 4582 31385
rect 4526 31311 4582 31320
rect 4540 30734 4568 31311
rect 4528 30728 4580 30734
rect 4528 30670 4580 30676
rect 4214 30492 4522 30512
rect 4214 30490 4220 30492
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4516 30490 4522 30492
rect 4276 30438 4278 30490
rect 4458 30438 4460 30490
rect 4214 30436 4220 30438
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4516 30436 4522 30438
rect 4214 30416 4522 30436
rect 4528 30320 4580 30326
rect 4528 30262 4580 30268
rect 4540 29594 4568 30262
rect 4632 30122 4660 31826
rect 4724 30870 4752 32166
rect 4816 31736 4844 35788
rect 4896 35692 4948 35698
rect 4896 35634 4948 35640
rect 4908 35290 4936 35634
rect 4896 35284 4948 35290
rect 4896 35226 4948 35232
rect 4988 35080 5040 35086
rect 4988 35022 5040 35028
rect 5000 32774 5028 35022
rect 4988 32768 5040 32774
rect 4988 32710 5040 32716
rect 4988 32428 5040 32434
rect 4988 32370 5040 32376
rect 4816 31708 4936 31736
rect 4908 31498 4936 31708
rect 4816 31470 4936 31498
rect 4712 30864 4764 30870
rect 4712 30806 4764 30812
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 4620 30116 4672 30122
rect 4620 30058 4672 30064
rect 4540 29566 4660 29594
rect 4214 29404 4522 29424
rect 4214 29402 4220 29404
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4516 29402 4522 29404
rect 4276 29350 4278 29402
rect 4458 29350 4460 29402
rect 4214 29348 4220 29350
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4516 29348 4522 29350
rect 4214 29328 4522 29348
rect 4068 28688 4120 28694
rect 4068 28630 4120 28636
rect 3896 28376 4108 28404
rect 3974 28248 4030 28257
rect 3974 28183 4030 28192
rect 3884 28076 3936 28082
rect 3884 28018 3936 28024
rect 3516 26240 3568 26246
rect 3514 26208 3516 26217
rect 3568 26208 3570 26217
rect 3620 26194 3648 26302
rect 3792 26308 3844 26314
rect 3792 26250 3844 26256
rect 3620 26166 3832 26194
rect 3514 26143 3570 26152
rect 3516 25832 3568 25838
rect 3516 25774 3568 25780
rect 3332 24812 3384 24818
rect 3332 24754 3384 24760
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3344 24721 3372 24754
rect 3330 24712 3386 24721
rect 3330 24647 3386 24656
rect 3332 24608 3384 24614
rect 3332 24550 3384 24556
rect 3422 24576 3478 24585
rect 3240 13932 3292 13938
rect 3240 13874 3292 13880
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3252 13025 3280 13262
rect 3238 13016 3294 13025
rect 3238 12951 3294 12960
rect 3240 12232 3292 12238
rect 3238 12200 3240 12209
rect 3292 12200 3294 12209
rect 3238 12135 3294 12144
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3344 11762 3372 24550
rect 3422 24511 3478 24520
rect 3436 22574 3464 24511
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3528 22094 3556 25774
rect 3700 25288 3752 25294
rect 3606 25256 3662 25265
rect 3700 25230 3752 25236
rect 3606 25191 3662 25200
rect 3620 23186 3648 25191
rect 3608 23180 3660 23186
rect 3608 23122 3660 23128
rect 3712 22710 3740 25230
rect 3700 22704 3752 22710
rect 3804 22681 3832 26166
rect 3896 26042 3924 28018
rect 3884 26036 3936 26042
rect 3884 25978 3936 25984
rect 3988 23730 4016 28183
rect 4080 27538 4108 28376
rect 4214 28316 4522 28336
rect 4214 28314 4220 28316
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4516 28314 4522 28316
rect 4276 28262 4278 28314
rect 4458 28262 4460 28314
rect 4214 28260 4220 28262
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4516 28260 4522 28262
rect 4214 28240 4522 28260
rect 4250 28112 4306 28121
rect 4250 28047 4306 28056
rect 4264 27577 4292 28047
rect 4436 27940 4488 27946
rect 4436 27882 4488 27888
rect 4250 27568 4306 27577
rect 4068 27532 4120 27538
rect 4250 27503 4306 27512
rect 4068 27474 4120 27480
rect 3976 23724 4028 23730
rect 3976 23666 4028 23672
rect 4080 23610 4108 27474
rect 4448 27441 4476 27882
rect 4632 27606 4660 29566
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 4434 27432 4490 27441
rect 4434 27367 4490 27376
rect 4620 27396 4672 27402
rect 4620 27338 4672 27344
rect 4214 27228 4522 27248
rect 4214 27226 4220 27228
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4516 27226 4522 27228
rect 4276 27174 4278 27226
rect 4458 27174 4460 27226
rect 4214 27172 4220 27174
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4516 27172 4522 27174
rect 4214 27152 4522 27172
rect 4214 26140 4522 26160
rect 4214 26138 4220 26140
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4516 26138 4522 26140
rect 4276 26086 4278 26138
rect 4458 26086 4460 26138
rect 4214 26084 4220 26086
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4516 26084 4522 26086
rect 4214 26064 4522 26084
rect 4526 25936 4582 25945
rect 4526 25871 4582 25880
rect 4540 25362 4568 25871
rect 4528 25356 4580 25362
rect 4528 25298 4580 25304
rect 4214 25052 4522 25072
rect 4214 25050 4220 25052
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4516 25050 4522 25052
rect 4276 24998 4278 25050
rect 4458 24998 4460 25050
rect 4214 24996 4220 24998
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4516 24996 4522 24998
rect 4214 24976 4522 24996
rect 4160 24812 4212 24818
rect 4160 24754 4212 24760
rect 4172 24274 4200 24754
rect 4632 24682 4660 27338
rect 4724 26518 4752 30670
rect 4816 26926 4844 31470
rect 5000 31362 5028 32370
rect 4908 31334 5028 31362
rect 4908 31210 4936 31334
rect 4986 31240 5042 31249
rect 4896 31204 4948 31210
rect 4986 31175 5042 31184
rect 4896 31146 4948 31152
rect 4896 30864 4948 30870
rect 4896 30806 4948 30812
rect 4804 26920 4856 26926
rect 4804 26862 4856 26868
rect 4908 26738 4936 30806
rect 5000 28218 5028 31175
rect 4988 28212 5040 28218
rect 4988 28154 5040 28160
rect 4988 26920 5040 26926
rect 4988 26862 5040 26868
rect 4816 26710 4936 26738
rect 4712 26512 4764 26518
rect 4712 26454 4764 26460
rect 4620 24676 4672 24682
rect 4620 24618 4672 24624
rect 4160 24268 4212 24274
rect 4160 24210 4212 24216
rect 4214 23964 4522 23984
rect 4214 23962 4220 23964
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4516 23962 4522 23964
rect 4276 23910 4278 23962
rect 4458 23910 4460 23962
rect 4214 23908 4220 23910
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4516 23908 4522 23910
rect 4214 23888 4522 23908
rect 3896 23582 4108 23610
rect 3700 22646 3752 22652
rect 3790 22672 3846 22681
rect 3608 22636 3660 22642
rect 3790 22607 3846 22616
rect 3608 22578 3660 22584
rect 3436 22066 3556 22094
rect 3436 21486 3464 22066
rect 3424 21480 3476 21486
rect 3424 21422 3476 21428
rect 3436 18970 3464 21422
rect 3620 21146 3648 22578
rect 3700 22432 3752 22438
rect 3700 22374 3752 22380
rect 3790 22400 3846 22409
rect 3712 22273 3740 22374
rect 3790 22335 3846 22344
rect 3698 22264 3754 22273
rect 3698 22199 3754 22208
rect 3608 21140 3660 21146
rect 3608 21082 3660 21088
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3620 19938 3648 20402
rect 3620 19910 3740 19938
rect 3424 18964 3476 18970
rect 3424 18906 3476 18912
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2870 9480 2926 9489
rect 2870 9415 2872 9424
rect 2924 9415 2926 9424
rect 2872 9386 2924 9392
rect 2582 9276 2890 9296
rect 2582 9274 2588 9276
rect 2644 9274 2668 9276
rect 2724 9274 2748 9276
rect 2804 9274 2828 9276
rect 2884 9274 2890 9276
rect 2644 9222 2646 9274
rect 2826 9222 2828 9274
rect 2582 9220 2588 9222
rect 2644 9220 2668 9222
rect 2724 9220 2748 9222
rect 2804 9220 2828 9222
rect 2884 9220 2890 9222
rect 2582 9200 2890 9220
rect 2962 9208 3018 9217
rect 2962 9143 2964 9152
rect 3016 9143 3018 9152
rect 2964 9114 3016 9120
rect 3068 9058 3096 9522
rect 2976 9030 3096 9058
rect 2976 8514 3004 9030
rect 3160 8974 3188 10610
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3068 8634 3096 8910
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2976 8486 3096 8514
rect 3252 8498 3280 9998
rect 2582 8188 2890 8208
rect 2582 8186 2588 8188
rect 2644 8186 2668 8188
rect 2724 8186 2748 8188
rect 2804 8186 2828 8188
rect 2884 8186 2890 8188
rect 2644 8134 2646 8186
rect 2826 8134 2828 8186
rect 2582 8132 2588 8134
rect 2644 8132 2668 8134
rect 2724 8132 2748 8134
rect 2804 8132 2828 8134
rect 2884 8132 2890 8134
rect 2582 8112 2890 8132
rect 3068 7886 3096 8486
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2582 7100 2890 7120
rect 2582 7098 2588 7100
rect 2644 7098 2668 7100
rect 2724 7098 2748 7100
rect 2804 7098 2828 7100
rect 2884 7098 2890 7100
rect 2644 7046 2646 7098
rect 2826 7046 2828 7098
rect 2582 7044 2588 7046
rect 2644 7044 2668 7046
rect 2724 7044 2748 7046
rect 2804 7044 2828 7046
rect 2884 7044 2890 7046
rect 2582 7024 2890 7044
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2582 6012 2890 6032
rect 2582 6010 2588 6012
rect 2644 6010 2668 6012
rect 2724 6010 2748 6012
rect 2804 6010 2828 6012
rect 2884 6010 2890 6012
rect 2644 5958 2646 6010
rect 2826 5958 2828 6010
rect 2582 5956 2588 5958
rect 2644 5956 2668 5958
rect 2724 5956 2748 5958
rect 2804 5956 2828 5958
rect 2884 5956 2890 5958
rect 2582 5936 2890 5956
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 1676 2916 1728 2922
rect 1676 2858 1728 2864
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 241 1440 2382
rect 2240 2310 2268 5102
rect 2582 4924 2890 4944
rect 2582 4922 2588 4924
rect 2644 4922 2668 4924
rect 2724 4922 2748 4924
rect 2804 4922 2828 4924
rect 2884 4922 2890 4924
rect 2644 4870 2646 4922
rect 2826 4870 2828 4922
rect 2582 4868 2588 4870
rect 2644 4868 2668 4870
rect 2724 4868 2748 4870
rect 2804 4868 2828 4870
rect 2884 4868 2890 4870
rect 2582 4848 2890 4868
rect 2976 4457 3004 6258
rect 2962 4448 3018 4457
rect 2962 4383 3018 4392
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2318 3224 2374 3233
rect 2318 3159 2374 3168
rect 2332 3058 2360 3159
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2424 2582 2452 4014
rect 2582 3836 2890 3856
rect 2582 3834 2588 3836
rect 2644 3834 2668 3836
rect 2724 3834 2748 3836
rect 2804 3834 2828 3836
rect 2884 3834 2890 3836
rect 2644 3782 2646 3834
rect 2826 3782 2828 3834
rect 2582 3780 2588 3782
rect 2644 3780 2668 3782
rect 2724 3780 2748 3782
rect 2804 3780 2828 3782
rect 2884 3780 2890 3782
rect 2582 3760 2890 3780
rect 2962 3632 3018 3641
rect 2962 3567 3018 3576
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2516 2990 2544 3470
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2700 3126 2728 3334
rect 2688 3120 2740 3126
rect 2688 3062 2740 3068
rect 2976 3058 3004 3567
rect 3068 3194 3096 7822
rect 3252 5710 3280 8434
rect 3344 6866 3372 11698
rect 3436 10266 3464 14962
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 3160 4570 3188 5238
rect 3252 4758 3280 5646
rect 3240 4752 3292 4758
rect 3344 4729 3372 6258
rect 3436 5778 3464 9930
rect 3528 7546 3556 13874
rect 3608 13796 3660 13802
rect 3608 13738 3660 13744
rect 3620 12322 3648 13738
rect 3712 12434 3740 19910
rect 3804 17814 3832 22335
rect 3896 20058 3924 23582
rect 4214 22876 4522 22896
rect 4214 22874 4220 22876
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4516 22874 4522 22876
rect 4276 22822 4278 22874
rect 4458 22822 4460 22874
rect 4214 22820 4220 22822
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4516 22820 4522 22822
rect 4214 22800 4522 22820
rect 3976 22704 4028 22710
rect 3976 22646 4028 22652
rect 3988 22030 4016 22646
rect 4160 22636 4212 22642
rect 4160 22578 4212 22584
rect 3976 22024 4028 22030
rect 4172 21978 4200 22578
rect 4620 22094 4672 22098
rect 4816 22094 4844 26710
rect 4896 26512 4948 26518
rect 4896 26454 4948 26460
rect 4908 24818 4936 26454
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4896 24676 4948 24682
rect 4896 24618 4948 24624
rect 4620 22092 4844 22094
rect 4672 22066 4844 22092
rect 4620 22034 4672 22040
rect 3976 21966 4028 21972
rect 3988 20466 4016 21966
rect 4080 21950 4200 21978
rect 4080 21690 4108 21950
rect 4214 21788 4522 21808
rect 4214 21786 4220 21788
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4516 21786 4522 21788
rect 4276 21734 4278 21786
rect 4458 21734 4460 21786
rect 4214 21732 4220 21734
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4516 21732 4522 21734
rect 4214 21712 4522 21732
rect 4908 21706 4936 24618
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 4724 21678 4936 21706
rect 4214 20700 4522 20720
rect 4214 20698 4220 20700
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4516 20698 4522 20700
rect 4276 20646 4278 20698
rect 4458 20646 4460 20698
rect 4214 20644 4220 20646
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4516 20644 4522 20646
rect 4214 20624 4522 20644
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 3976 19848 4028 19854
rect 3974 19816 3976 19825
rect 4028 19816 4030 19825
rect 3974 19751 4030 19760
rect 4214 19612 4522 19632
rect 4214 19610 4220 19612
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4516 19610 4522 19612
rect 4276 19558 4278 19610
rect 4458 19558 4460 19610
rect 4214 19556 4220 19558
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4516 19556 4522 19558
rect 4214 19536 4522 19556
rect 4214 18524 4522 18544
rect 4214 18522 4220 18524
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4516 18522 4522 18524
rect 4276 18470 4278 18522
rect 4458 18470 4460 18522
rect 4214 18468 4220 18470
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4516 18468 4522 18470
rect 4214 18448 4522 18468
rect 3792 17808 3844 17814
rect 3792 17750 3844 17756
rect 4214 17436 4522 17456
rect 4214 17434 4220 17436
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4516 17434 4522 17436
rect 4276 17382 4278 17434
rect 4458 17382 4460 17434
rect 4214 17380 4220 17382
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4516 17380 4522 17382
rect 4214 17360 4522 17380
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3792 16448 3844 16454
rect 3988 16425 4016 16526
rect 3792 16390 3844 16396
rect 3974 16416 4030 16425
rect 3804 16182 3832 16390
rect 3974 16351 4030 16360
rect 4214 16348 4522 16368
rect 4214 16346 4220 16348
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4516 16346 4522 16348
rect 4276 16294 4278 16346
rect 4458 16294 4460 16346
rect 4214 16292 4220 16294
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4516 16292 4522 16294
rect 4214 16272 4522 16292
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3804 15706 3832 15982
rect 3792 15700 3844 15706
rect 3792 15642 3844 15648
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3988 15201 4016 15438
rect 3974 15192 4030 15201
rect 3974 15127 4030 15136
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3804 13462 3832 14350
rect 3988 14249 4016 14350
rect 3974 14240 4030 14249
rect 3974 14175 4030 14184
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3792 13456 3844 13462
rect 3896 13433 3924 13874
rect 3974 13832 4030 13841
rect 3974 13767 4030 13776
rect 3792 13398 3844 13404
rect 3882 13424 3938 13433
rect 3882 13359 3938 13368
rect 3988 13326 4016 13767
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 4080 12434 4108 16050
rect 4214 15260 4522 15280
rect 4214 15258 4220 15260
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4516 15258 4522 15260
rect 4276 15206 4278 15258
rect 4458 15206 4460 15258
rect 4214 15204 4220 15206
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4516 15204 4522 15206
rect 4214 15184 4522 15204
rect 4214 14172 4522 14192
rect 4214 14170 4220 14172
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4516 14170 4522 14172
rect 4276 14118 4278 14170
rect 4458 14118 4460 14170
rect 4214 14116 4220 14118
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4516 14116 4522 14118
rect 4214 14096 4522 14116
rect 4214 13084 4522 13104
rect 4214 13082 4220 13084
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4516 13082 4522 13084
rect 4276 13030 4278 13082
rect 4458 13030 4460 13082
rect 4214 13028 4220 13030
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4516 13028 4522 13030
rect 4214 13008 4522 13028
rect 3712 12406 3924 12434
rect 3620 12294 3832 12322
rect 3608 12164 3660 12170
rect 3608 12106 3660 12112
rect 3620 9586 3648 12106
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3620 6186 3648 9522
rect 3712 8634 3740 9522
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3698 8528 3754 8537
rect 3698 8463 3754 8472
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3712 6066 3740 8463
rect 3528 6038 3740 6066
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3240 4694 3292 4700
rect 3330 4720 3386 4729
rect 3330 4655 3386 4664
rect 3240 4616 3292 4622
rect 3160 4564 3240 4570
rect 3160 4558 3292 4564
rect 3160 4542 3280 4558
rect 3160 4146 3188 4542
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2516 2650 2544 2926
rect 2582 2748 2890 2768
rect 2582 2746 2588 2748
rect 2644 2746 2668 2748
rect 2724 2746 2748 2748
rect 2804 2746 2828 2748
rect 2884 2746 2890 2748
rect 2644 2694 2646 2746
rect 2826 2694 2828 2746
rect 2582 2692 2588 2694
rect 2644 2692 2668 2694
rect 2724 2692 2748 2694
rect 2804 2692 2828 2694
rect 2884 2692 2890 2694
rect 2582 2672 2890 2692
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2412 2576 2464 2582
rect 2412 2518 2464 2524
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2228 2304 2280 2310
rect 2792 2281 2820 2450
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2228 2246 2280 2252
rect 2778 2272 2834 2281
rect 2778 2207 2834 2216
rect 2780 1080 2832 1086
rect 2778 1048 2780 1057
rect 2832 1048 2834 1057
rect 2778 983 2834 992
rect 2884 649 2912 2382
rect 3344 2378 3372 4422
rect 3436 2854 3464 5714
rect 3528 5370 3556 6038
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3528 3738 3556 5170
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3620 3534 3648 5578
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3712 5273 3740 5306
rect 3698 5264 3754 5273
rect 3698 5199 3754 5208
rect 3804 4486 3832 12294
rect 3896 5710 3924 12406
rect 3988 12406 4108 12434
rect 3988 10674 4016 12406
rect 4214 11996 4522 12016
rect 4214 11994 4220 11996
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4516 11994 4522 11996
rect 4276 11942 4278 11994
rect 4458 11942 4460 11994
rect 4214 11940 4220 11942
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4516 11940 4522 11942
rect 4214 11920 4522 11940
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3988 9081 4016 10610
rect 3974 9072 4030 9081
rect 3974 9007 4030 9016
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3988 6458 4016 8910
rect 4080 7410 4108 11018
rect 4214 10908 4522 10928
rect 4214 10906 4220 10908
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4516 10906 4522 10908
rect 4276 10854 4278 10906
rect 4458 10854 4460 10906
rect 4214 10852 4220 10854
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4516 10852 4522 10854
rect 4214 10832 4522 10852
rect 4632 10606 4660 17138
rect 4724 11150 4752 21678
rect 4804 21616 4856 21622
rect 4804 21558 4856 21564
rect 4816 17746 4844 21558
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4816 14822 4844 17682
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4908 14482 4936 15438
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 5000 13954 5028 26862
rect 5092 26790 5120 40870
rect 5184 35222 5212 41160
rect 5356 41064 5408 41070
rect 5356 41006 5408 41012
rect 5262 40896 5318 40905
rect 5262 40831 5318 40840
rect 5172 35216 5224 35222
rect 5172 35158 5224 35164
rect 5172 35080 5224 35086
rect 5172 35022 5224 35028
rect 5184 32298 5212 35022
rect 5172 32292 5224 32298
rect 5172 32234 5224 32240
rect 5170 32192 5226 32201
rect 5170 32127 5226 32136
rect 5184 28082 5212 32127
rect 5172 28076 5224 28082
rect 5172 28018 5224 28024
rect 5170 27976 5226 27985
rect 5170 27911 5226 27920
rect 5080 26784 5132 26790
rect 5080 26726 5132 26732
rect 5080 26580 5132 26586
rect 5080 26522 5132 26528
rect 5092 22710 5120 26522
rect 5080 22704 5132 22710
rect 5080 22646 5132 22652
rect 5184 16658 5212 27911
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 4816 13926 5028 13954
rect 4816 11354 4844 13926
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 5276 10538 5304 40831
rect 5368 31890 5396 41006
rect 5356 31884 5408 31890
rect 5356 31826 5408 31832
rect 5356 31340 5408 31346
rect 5356 31282 5408 31288
rect 5368 28218 5396 31282
rect 5460 28257 5488 50798
rect 5552 45830 5580 72490
rect 5846 72380 6154 72400
rect 5846 72378 5852 72380
rect 5908 72378 5932 72380
rect 5988 72378 6012 72380
rect 6068 72378 6092 72380
rect 6148 72378 6154 72380
rect 5908 72326 5910 72378
rect 6090 72326 6092 72378
rect 5846 72324 5852 72326
rect 5908 72324 5932 72326
rect 5988 72324 6012 72326
rect 6068 72324 6092 72326
rect 6148 72324 6154 72326
rect 5846 72304 6154 72324
rect 7478 71836 7786 71856
rect 7478 71834 7484 71836
rect 7540 71834 7564 71836
rect 7620 71834 7644 71836
rect 7700 71834 7724 71836
rect 7780 71834 7786 71836
rect 7540 71782 7542 71834
rect 7722 71782 7724 71834
rect 7478 71780 7484 71782
rect 7540 71780 7564 71782
rect 7620 71780 7644 71782
rect 7700 71780 7724 71782
rect 7780 71780 7786 71782
rect 7478 71760 7786 71780
rect 5632 71460 5684 71466
rect 5632 71402 5684 71408
rect 5644 46510 5672 71402
rect 5846 71292 6154 71312
rect 5846 71290 5852 71292
rect 5908 71290 5932 71292
rect 5988 71290 6012 71292
rect 6068 71290 6092 71292
rect 6148 71290 6154 71292
rect 5908 71238 5910 71290
rect 6090 71238 6092 71290
rect 5846 71236 5852 71238
rect 5908 71236 5932 71238
rect 5988 71236 6012 71238
rect 6068 71236 6092 71238
rect 6148 71236 6154 71238
rect 5846 71216 6154 71236
rect 7478 70748 7786 70768
rect 7478 70746 7484 70748
rect 7540 70746 7564 70748
rect 7620 70746 7644 70748
rect 7700 70746 7724 70748
rect 7780 70746 7786 70748
rect 7540 70694 7542 70746
rect 7722 70694 7724 70746
rect 7478 70692 7484 70694
rect 7540 70692 7564 70694
rect 7620 70692 7644 70694
rect 7700 70692 7724 70694
rect 7780 70692 7786 70694
rect 7478 70672 7786 70692
rect 5846 70204 6154 70224
rect 5846 70202 5852 70204
rect 5908 70202 5932 70204
rect 5988 70202 6012 70204
rect 6068 70202 6092 70204
rect 6148 70202 6154 70204
rect 5908 70150 5910 70202
rect 6090 70150 6092 70202
rect 5846 70148 5852 70150
rect 5908 70148 5932 70150
rect 5988 70148 6012 70150
rect 6068 70148 6092 70150
rect 6148 70148 6154 70150
rect 5846 70128 6154 70148
rect 7478 69660 7786 69680
rect 7478 69658 7484 69660
rect 7540 69658 7564 69660
rect 7620 69658 7644 69660
rect 7700 69658 7724 69660
rect 7780 69658 7786 69660
rect 7540 69606 7542 69658
rect 7722 69606 7724 69658
rect 7478 69604 7484 69606
rect 7540 69604 7564 69606
rect 7620 69604 7644 69606
rect 7700 69604 7724 69606
rect 7780 69604 7786 69606
rect 7478 69584 7786 69604
rect 5724 69284 5776 69290
rect 5724 69226 5776 69232
rect 5736 46578 5764 69226
rect 5846 69116 6154 69136
rect 5846 69114 5852 69116
rect 5908 69114 5932 69116
rect 5988 69114 6012 69116
rect 6068 69114 6092 69116
rect 6148 69114 6154 69116
rect 5908 69062 5910 69114
rect 6090 69062 6092 69114
rect 5846 69060 5852 69062
rect 5908 69060 5932 69062
rect 5988 69060 6012 69062
rect 6068 69060 6092 69062
rect 6148 69060 6154 69062
rect 5846 69040 6154 69060
rect 7478 68572 7786 68592
rect 7478 68570 7484 68572
rect 7540 68570 7564 68572
rect 7620 68570 7644 68572
rect 7700 68570 7724 68572
rect 7780 68570 7786 68572
rect 7540 68518 7542 68570
rect 7722 68518 7724 68570
rect 7478 68516 7484 68518
rect 7540 68516 7564 68518
rect 7620 68516 7644 68518
rect 7700 68516 7724 68518
rect 7780 68516 7786 68518
rect 7478 68496 7786 68516
rect 5846 68028 6154 68048
rect 5846 68026 5852 68028
rect 5908 68026 5932 68028
rect 5988 68026 6012 68028
rect 6068 68026 6092 68028
rect 6148 68026 6154 68028
rect 5908 67974 5910 68026
rect 6090 67974 6092 68026
rect 5846 67972 5852 67974
rect 5908 67972 5932 67974
rect 5988 67972 6012 67974
rect 6068 67972 6092 67974
rect 6148 67972 6154 67974
rect 5846 67952 6154 67972
rect 7478 67484 7786 67504
rect 7478 67482 7484 67484
rect 7540 67482 7564 67484
rect 7620 67482 7644 67484
rect 7700 67482 7724 67484
rect 7780 67482 7786 67484
rect 7540 67430 7542 67482
rect 7722 67430 7724 67482
rect 7478 67428 7484 67430
rect 7540 67428 7564 67430
rect 7620 67428 7644 67430
rect 7700 67428 7724 67430
rect 7780 67428 7786 67430
rect 7478 67408 7786 67428
rect 5846 66940 6154 66960
rect 5846 66938 5852 66940
rect 5908 66938 5932 66940
rect 5988 66938 6012 66940
rect 6068 66938 6092 66940
rect 6148 66938 6154 66940
rect 5908 66886 5910 66938
rect 6090 66886 6092 66938
rect 5846 66884 5852 66886
rect 5908 66884 5932 66886
rect 5988 66884 6012 66886
rect 6068 66884 6092 66886
rect 6148 66884 6154 66886
rect 5846 66864 6154 66884
rect 7478 66396 7786 66416
rect 7478 66394 7484 66396
rect 7540 66394 7564 66396
rect 7620 66394 7644 66396
rect 7700 66394 7724 66396
rect 7780 66394 7786 66396
rect 7540 66342 7542 66394
rect 7722 66342 7724 66394
rect 7478 66340 7484 66342
rect 7540 66340 7564 66342
rect 7620 66340 7644 66342
rect 7700 66340 7724 66342
rect 7780 66340 7786 66342
rect 7478 66320 7786 66340
rect 5846 65852 6154 65872
rect 5846 65850 5852 65852
rect 5908 65850 5932 65852
rect 5988 65850 6012 65852
rect 6068 65850 6092 65852
rect 6148 65850 6154 65852
rect 5908 65798 5910 65850
rect 6090 65798 6092 65850
rect 5846 65796 5852 65798
rect 5908 65796 5932 65798
rect 5988 65796 6012 65798
rect 6068 65796 6092 65798
rect 6148 65796 6154 65798
rect 5846 65776 6154 65796
rect 7852 65482 7880 77386
rect 8300 77376 8352 77382
rect 8300 77318 8352 77324
rect 8312 74798 8340 77318
rect 9416 77217 9444 77454
rect 9402 77208 9458 77217
rect 9402 77143 9458 77152
rect 9508 77042 9536 77959
rect 9600 77042 9628 78639
rect 9968 77518 9996 79455
rect 9956 77512 10008 77518
rect 9956 77454 10008 77460
rect 9496 77036 9548 77042
rect 9496 76978 9548 76984
rect 9588 77036 9640 77042
rect 9588 76978 9640 76984
rect 9772 76832 9824 76838
rect 9772 76774 9824 76780
rect 9110 76732 9418 76752
rect 9110 76730 9116 76732
rect 9172 76730 9196 76732
rect 9252 76730 9276 76732
rect 9332 76730 9356 76732
rect 9412 76730 9418 76732
rect 9172 76678 9174 76730
rect 9354 76678 9356 76730
rect 9110 76676 9116 76678
rect 9172 76676 9196 76678
rect 9252 76676 9276 76678
rect 9332 76676 9356 76678
rect 9412 76676 9418 76678
rect 9110 76656 9418 76676
rect 9110 75644 9418 75664
rect 9110 75642 9116 75644
rect 9172 75642 9196 75644
rect 9252 75642 9276 75644
rect 9332 75642 9356 75644
rect 9412 75642 9418 75644
rect 9172 75590 9174 75642
rect 9354 75590 9356 75642
rect 9110 75588 9116 75590
rect 9172 75588 9196 75590
rect 9252 75588 9276 75590
rect 9332 75588 9356 75590
rect 9412 75588 9418 75590
rect 9110 75568 9418 75588
rect 8300 74792 8352 74798
rect 8300 74734 8352 74740
rect 9110 74556 9418 74576
rect 9110 74554 9116 74556
rect 9172 74554 9196 74556
rect 9252 74554 9276 74556
rect 9332 74554 9356 74556
rect 9412 74554 9418 74556
rect 9172 74502 9174 74554
rect 9354 74502 9356 74554
rect 9110 74500 9116 74502
rect 9172 74500 9196 74502
rect 9252 74500 9276 74502
rect 9332 74500 9356 74502
rect 9412 74500 9418 74502
rect 9110 74480 9418 74500
rect 8300 73568 8352 73574
rect 8300 73510 8352 73516
rect 8312 72758 8340 73510
rect 9110 73468 9418 73488
rect 9110 73466 9116 73468
rect 9172 73466 9196 73468
rect 9252 73466 9276 73468
rect 9332 73466 9356 73468
rect 9412 73466 9418 73468
rect 9172 73414 9174 73466
rect 9354 73414 9356 73466
rect 9110 73412 9116 73414
rect 9172 73412 9196 73414
rect 9252 73412 9276 73414
rect 9332 73412 9356 73414
rect 9412 73412 9418 73414
rect 9110 73392 9418 73412
rect 8300 72752 8352 72758
rect 8300 72694 8352 72700
rect 9110 72380 9418 72400
rect 9110 72378 9116 72380
rect 9172 72378 9196 72380
rect 9252 72378 9276 72380
rect 9332 72378 9356 72380
rect 9412 72378 9418 72380
rect 9172 72326 9174 72378
rect 9354 72326 9356 72378
rect 9110 72324 9116 72326
rect 9172 72324 9196 72326
rect 9252 72324 9276 72326
rect 9332 72324 9356 72326
rect 9412 72324 9418 72326
rect 9110 72304 9418 72324
rect 9110 71292 9418 71312
rect 9110 71290 9116 71292
rect 9172 71290 9196 71292
rect 9252 71290 9276 71292
rect 9332 71290 9356 71292
rect 9412 71290 9418 71292
rect 9172 71238 9174 71290
rect 9354 71238 9356 71290
rect 9110 71236 9116 71238
rect 9172 71236 9196 71238
rect 9252 71236 9276 71238
rect 9332 71236 9356 71238
rect 9412 71236 9418 71238
rect 9110 71216 9418 71236
rect 9110 70204 9418 70224
rect 9110 70202 9116 70204
rect 9172 70202 9196 70204
rect 9252 70202 9276 70204
rect 9332 70202 9356 70204
rect 9412 70202 9418 70204
rect 9172 70150 9174 70202
rect 9354 70150 9356 70202
rect 9110 70148 9116 70150
rect 9172 70148 9196 70150
rect 9252 70148 9276 70150
rect 9332 70148 9356 70150
rect 9412 70148 9418 70150
rect 9110 70128 9418 70148
rect 9110 69116 9418 69136
rect 9110 69114 9116 69116
rect 9172 69114 9196 69116
rect 9252 69114 9276 69116
rect 9332 69114 9356 69116
rect 9412 69114 9418 69116
rect 9172 69062 9174 69114
rect 9354 69062 9356 69114
rect 9110 69060 9116 69062
rect 9172 69060 9196 69062
rect 9252 69060 9276 69062
rect 9332 69060 9356 69062
rect 9412 69060 9418 69062
rect 9110 69040 9418 69060
rect 8300 68128 8352 68134
rect 8300 68070 8352 68076
rect 8312 66842 8340 68070
rect 9110 68028 9418 68048
rect 9110 68026 9116 68028
rect 9172 68026 9196 68028
rect 9252 68026 9276 68028
rect 9332 68026 9356 68028
rect 9412 68026 9418 68028
rect 9172 67974 9174 68026
rect 9354 67974 9356 68026
rect 9110 67972 9116 67974
rect 9172 67972 9196 67974
rect 9252 67972 9276 67974
rect 9332 67972 9356 67974
rect 9412 67972 9418 67974
rect 9110 67952 9418 67972
rect 9110 66940 9418 66960
rect 9110 66938 9116 66940
rect 9172 66938 9196 66940
rect 9252 66938 9276 66940
rect 9332 66938 9356 66940
rect 9412 66938 9418 66940
rect 9172 66886 9174 66938
rect 9354 66886 9356 66938
rect 9110 66884 9116 66886
rect 9172 66884 9196 66886
rect 9252 66884 9276 66886
rect 9332 66884 9356 66886
rect 9412 66884 9418 66886
rect 9110 66864 9418 66884
rect 8300 66836 8352 66842
rect 8300 66778 8352 66784
rect 8300 66496 8352 66502
rect 8300 66438 8352 66444
rect 7840 65476 7892 65482
rect 7840 65418 7892 65424
rect 7478 65308 7786 65328
rect 7478 65306 7484 65308
rect 7540 65306 7564 65308
rect 7620 65306 7644 65308
rect 7700 65306 7724 65308
rect 7780 65306 7786 65308
rect 7540 65254 7542 65306
rect 7722 65254 7724 65306
rect 7478 65252 7484 65254
rect 7540 65252 7564 65254
rect 7620 65252 7644 65254
rect 7700 65252 7724 65254
rect 7780 65252 7786 65254
rect 7478 65232 7786 65252
rect 8312 65210 8340 66438
rect 9110 65852 9418 65872
rect 9110 65850 9116 65852
rect 9172 65850 9196 65852
rect 9252 65850 9276 65852
rect 9332 65850 9356 65852
rect 9412 65850 9418 65852
rect 9172 65798 9174 65850
rect 9354 65798 9356 65850
rect 9110 65796 9116 65798
rect 9172 65796 9196 65798
rect 9252 65796 9276 65798
rect 9332 65796 9356 65798
rect 9412 65796 9418 65798
rect 9110 65776 9418 65796
rect 8300 65204 8352 65210
rect 8300 65146 8352 65152
rect 8300 64932 8352 64938
rect 8300 64874 8352 64880
rect 5846 64764 6154 64784
rect 5846 64762 5852 64764
rect 5908 64762 5932 64764
rect 5988 64762 6012 64764
rect 6068 64762 6092 64764
rect 6148 64762 6154 64764
rect 5908 64710 5910 64762
rect 6090 64710 6092 64762
rect 5846 64708 5852 64710
rect 5908 64708 5932 64710
rect 5988 64708 6012 64710
rect 6068 64708 6092 64710
rect 6148 64708 6154 64710
rect 5846 64688 6154 64708
rect 8312 64530 8340 64874
rect 9110 64764 9418 64784
rect 9110 64762 9116 64764
rect 9172 64762 9196 64764
rect 9252 64762 9276 64764
rect 9332 64762 9356 64764
rect 9412 64762 9418 64764
rect 9172 64710 9174 64762
rect 9354 64710 9356 64762
rect 9110 64708 9116 64710
rect 9172 64708 9196 64710
rect 9252 64708 9276 64710
rect 9332 64708 9356 64710
rect 9412 64708 9418 64710
rect 9110 64688 9418 64708
rect 8300 64524 8352 64530
rect 8300 64466 8352 64472
rect 8300 64320 8352 64326
rect 8300 64262 8352 64268
rect 7478 64220 7786 64240
rect 7478 64218 7484 64220
rect 7540 64218 7564 64220
rect 7620 64218 7644 64220
rect 7700 64218 7724 64220
rect 7780 64218 7786 64220
rect 7540 64166 7542 64218
rect 7722 64166 7724 64218
rect 7478 64164 7484 64166
rect 7540 64164 7564 64166
rect 7620 64164 7644 64166
rect 7700 64164 7724 64166
rect 7780 64164 7786 64166
rect 7478 64144 7786 64164
rect 5846 63676 6154 63696
rect 5846 63674 5852 63676
rect 5908 63674 5932 63676
rect 5988 63674 6012 63676
rect 6068 63674 6092 63676
rect 6148 63674 6154 63676
rect 5908 63622 5910 63674
rect 6090 63622 6092 63674
rect 5846 63620 5852 63622
rect 5908 63620 5932 63622
rect 5988 63620 6012 63622
rect 6068 63620 6092 63622
rect 6148 63620 6154 63622
rect 5846 63600 6154 63620
rect 7478 63132 7786 63152
rect 7478 63130 7484 63132
rect 7540 63130 7564 63132
rect 7620 63130 7644 63132
rect 7700 63130 7724 63132
rect 7780 63130 7786 63132
rect 7540 63078 7542 63130
rect 7722 63078 7724 63130
rect 7478 63076 7484 63078
rect 7540 63076 7564 63078
rect 7620 63076 7644 63078
rect 7700 63076 7724 63078
rect 7780 63076 7786 63078
rect 7478 63056 7786 63076
rect 6184 62688 6236 62694
rect 6184 62630 6236 62636
rect 5846 62588 6154 62608
rect 5846 62586 5852 62588
rect 5908 62586 5932 62588
rect 5988 62586 6012 62588
rect 6068 62586 6092 62588
rect 6148 62586 6154 62588
rect 5908 62534 5910 62586
rect 6090 62534 6092 62586
rect 5846 62532 5852 62534
rect 5908 62532 5932 62534
rect 5988 62532 6012 62534
rect 6068 62532 6092 62534
rect 6148 62532 6154 62534
rect 5846 62512 6154 62532
rect 5846 61500 6154 61520
rect 5846 61498 5852 61500
rect 5908 61498 5932 61500
rect 5988 61498 6012 61500
rect 6068 61498 6092 61500
rect 6148 61498 6154 61500
rect 5908 61446 5910 61498
rect 6090 61446 6092 61498
rect 5846 61444 5852 61446
rect 5908 61444 5932 61446
rect 5988 61444 6012 61446
rect 6068 61444 6092 61446
rect 6148 61444 6154 61446
rect 5846 61424 6154 61444
rect 5846 60412 6154 60432
rect 5846 60410 5852 60412
rect 5908 60410 5932 60412
rect 5988 60410 6012 60412
rect 6068 60410 6092 60412
rect 6148 60410 6154 60412
rect 5908 60358 5910 60410
rect 6090 60358 6092 60410
rect 5846 60356 5852 60358
rect 5908 60356 5932 60358
rect 5988 60356 6012 60358
rect 6068 60356 6092 60358
rect 6148 60356 6154 60358
rect 5846 60336 6154 60356
rect 6196 60081 6224 62630
rect 8312 62354 8340 64262
rect 9110 63676 9418 63696
rect 9110 63674 9116 63676
rect 9172 63674 9196 63676
rect 9252 63674 9276 63676
rect 9332 63674 9356 63676
rect 9412 63674 9418 63676
rect 9172 63622 9174 63674
rect 9354 63622 9356 63674
rect 9110 63620 9116 63622
rect 9172 63620 9196 63622
rect 9252 63620 9276 63622
rect 9332 63620 9356 63622
rect 9412 63620 9418 63622
rect 9110 63600 9418 63620
rect 8484 63232 8536 63238
rect 8484 63174 8536 63180
rect 8300 62348 8352 62354
rect 8300 62290 8352 62296
rect 8300 62144 8352 62150
rect 8300 62086 8352 62092
rect 7478 62044 7786 62064
rect 7478 62042 7484 62044
rect 7540 62042 7564 62044
rect 7620 62042 7644 62044
rect 7700 62042 7724 62044
rect 7780 62042 7786 62044
rect 7540 61990 7542 62042
rect 7722 61990 7724 62042
rect 7478 61988 7484 61990
rect 7540 61988 7564 61990
rect 7620 61988 7644 61990
rect 7700 61988 7724 61990
rect 7780 61988 7786 61990
rect 7478 61968 7786 61988
rect 8312 61266 8340 62086
rect 8300 61260 8352 61266
rect 8300 61202 8352 61208
rect 7478 60956 7786 60976
rect 7478 60954 7484 60956
rect 7540 60954 7564 60956
rect 7620 60954 7644 60956
rect 7700 60954 7724 60956
rect 7780 60954 7786 60956
rect 7540 60902 7542 60954
rect 7722 60902 7724 60954
rect 7478 60900 7484 60902
rect 7540 60900 7564 60902
rect 7620 60900 7644 60902
rect 7700 60900 7724 60902
rect 7780 60900 7786 60902
rect 7478 60880 7786 60900
rect 6182 60072 6238 60081
rect 6182 60007 6238 60016
rect 7478 59868 7786 59888
rect 7478 59866 7484 59868
rect 7540 59866 7564 59868
rect 7620 59866 7644 59868
rect 7700 59866 7724 59868
rect 7780 59866 7786 59868
rect 7540 59814 7542 59866
rect 7722 59814 7724 59866
rect 7478 59812 7484 59814
rect 7540 59812 7564 59814
rect 7620 59812 7644 59814
rect 7700 59812 7724 59814
rect 7780 59812 7786 59814
rect 7478 59792 7786 59812
rect 8300 59424 8352 59430
rect 8300 59366 8352 59372
rect 5846 59324 6154 59344
rect 5846 59322 5852 59324
rect 5908 59322 5932 59324
rect 5988 59322 6012 59324
rect 6068 59322 6092 59324
rect 6148 59322 6154 59324
rect 5908 59270 5910 59322
rect 6090 59270 6092 59322
rect 5846 59268 5852 59270
rect 5908 59268 5932 59270
rect 5988 59268 6012 59270
rect 6068 59268 6092 59270
rect 6148 59268 6154 59270
rect 5846 59248 6154 59268
rect 7478 58780 7786 58800
rect 7478 58778 7484 58780
rect 7540 58778 7564 58780
rect 7620 58778 7644 58780
rect 7700 58778 7724 58780
rect 7780 58778 7786 58780
rect 7540 58726 7542 58778
rect 7722 58726 7724 58778
rect 7478 58724 7484 58726
rect 7540 58724 7564 58726
rect 7620 58724 7644 58726
rect 7700 58724 7724 58726
rect 7780 58724 7786 58726
rect 7478 58704 7786 58724
rect 5846 58236 6154 58256
rect 5846 58234 5852 58236
rect 5908 58234 5932 58236
rect 5988 58234 6012 58236
rect 6068 58234 6092 58236
rect 6148 58234 6154 58236
rect 5908 58182 5910 58234
rect 6090 58182 6092 58234
rect 5846 58180 5852 58182
rect 5908 58180 5932 58182
rect 5988 58180 6012 58182
rect 6068 58180 6092 58182
rect 6148 58180 6154 58182
rect 5846 58160 6154 58180
rect 7478 57692 7786 57712
rect 7478 57690 7484 57692
rect 7540 57690 7564 57692
rect 7620 57690 7644 57692
rect 7700 57690 7724 57692
rect 7780 57690 7786 57692
rect 7540 57638 7542 57690
rect 7722 57638 7724 57690
rect 7478 57636 7484 57638
rect 7540 57636 7564 57638
rect 7620 57636 7644 57638
rect 7700 57636 7724 57638
rect 7780 57636 7786 57638
rect 7478 57616 7786 57636
rect 6552 57452 6604 57458
rect 6552 57394 6604 57400
rect 5846 57148 6154 57168
rect 5846 57146 5852 57148
rect 5908 57146 5932 57148
rect 5988 57146 6012 57148
rect 6068 57146 6092 57148
rect 6148 57146 6154 57148
rect 5908 57094 5910 57146
rect 6090 57094 6092 57146
rect 5846 57092 5852 57094
rect 5908 57092 5932 57094
rect 5988 57092 6012 57094
rect 6068 57092 6092 57094
rect 6148 57092 6154 57094
rect 5846 57072 6154 57092
rect 6368 56296 6420 56302
rect 6368 56238 6420 56244
rect 6184 56160 6236 56166
rect 6184 56102 6236 56108
rect 5846 56060 6154 56080
rect 5846 56058 5852 56060
rect 5908 56058 5932 56060
rect 5988 56058 6012 56060
rect 6068 56058 6092 56060
rect 6148 56058 6154 56060
rect 5908 56006 5910 56058
rect 6090 56006 6092 56058
rect 5846 56004 5852 56006
rect 5908 56004 5932 56006
rect 5988 56004 6012 56006
rect 6068 56004 6092 56006
rect 6148 56004 6154 56006
rect 5846 55984 6154 56004
rect 5846 54972 6154 54992
rect 5846 54970 5852 54972
rect 5908 54970 5932 54972
rect 5988 54970 6012 54972
rect 6068 54970 6092 54972
rect 6148 54970 6154 54972
rect 5908 54918 5910 54970
rect 6090 54918 6092 54970
rect 5846 54916 5852 54918
rect 5908 54916 5932 54918
rect 5988 54916 6012 54918
rect 6068 54916 6092 54918
rect 6148 54916 6154 54918
rect 5846 54896 6154 54916
rect 6196 54602 6224 56102
rect 6276 54664 6328 54670
rect 6276 54606 6328 54612
rect 6184 54596 6236 54602
rect 6184 54538 6236 54544
rect 5846 53884 6154 53904
rect 5846 53882 5852 53884
rect 5908 53882 5932 53884
rect 5988 53882 6012 53884
rect 6068 53882 6092 53884
rect 6148 53882 6154 53884
rect 5908 53830 5910 53882
rect 6090 53830 6092 53882
rect 5846 53828 5852 53830
rect 5908 53828 5932 53830
rect 5988 53828 6012 53830
rect 6068 53828 6092 53830
rect 6148 53828 6154 53830
rect 5846 53808 6154 53828
rect 5846 52796 6154 52816
rect 5846 52794 5852 52796
rect 5908 52794 5932 52796
rect 5988 52794 6012 52796
rect 6068 52794 6092 52796
rect 6148 52794 6154 52796
rect 5908 52742 5910 52794
rect 6090 52742 6092 52794
rect 5846 52740 5852 52742
rect 5908 52740 5932 52742
rect 5988 52740 6012 52742
rect 6068 52740 6092 52742
rect 6148 52740 6154 52742
rect 5846 52720 6154 52740
rect 5846 51708 6154 51728
rect 5846 51706 5852 51708
rect 5908 51706 5932 51708
rect 5988 51706 6012 51708
rect 6068 51706 6092 51708
rect 6148 51706 6154 51708
rect 5908 51654 5910 51706
rect 6090 51654 6092 51706
rect 5846 51652 5852 51654
rect 5908 51652 5932 51654
rect 5988 51652 6012 51654
rect 6068 51652 6092 51654
rect 6148 51652 6154 51654
rect 5846 51632 6154 51652
rect 6184 50788 6236 50794
rect 6184 50730 6236 50736
rect 5846 50620 6154 50640
rect 5846 50618 5852 50620
rect 5908 50618 5932 50620
rect 5988 50618 6012 50620
rect 6068 50618 6092 50620
rect 6148 50618 6154 50620
rect 5908 50566 5910 50618
rect 6090 50566 6092 50618
rect 5846 50564 5852 50566
rect 5908 50564 5932 50566
rect 5988 50564 6012 50566
rect 6068 50564 6092 50566
rect 6148 50564 6154 50566
rect 5846 50544 6154 50564
rect 5846 49532 6154 49552
rect 5846 49530 5852 49532
rect 5908 49530 5932 49532
rect 5988 49530 6012 49532
rect 6068 49530 6092 49532
rect 6148 49530 6154 49532
rect 5908 49478 5910 49530
rect 6090 49478 6092 49530
rect 5846 49476 5852 49478
rect 5908 49476 5932 49478
rect 5988 49476 6012 49478
rect 6068 49476 6092 49478
rect 6148 49476 6154 49478
rect 5846 49456 6154 49476
rect 5846 48444 6154 48464
rect 5846 48442 5852 48444
rect 5908 48442 5932 48444
rect 5988 48442 6012 48444
rect 6068 48442 6092 48444
rect 6148 48442 6154 48444
rect 5908 48390 5910 48442
rect 6090 48390 6092 48442
rect 5846 48388 5852 48390
rect 5908 48388 5932 48390
rect 5988 48388 6012 48390
rect 6068 48388 6092 48390
rect 6148 48388 6154 48390
rect 5846 48368 6154 48388
rect 6196 48278 6224 50730
rect 6184 48272 6236 48278
rect 6184 48214 6236 48220
rect 6184 48068 6236 48074
rect 6184 48010 6236 48016
rect 5846 47356 6154 47376
rect 5846 47354 5852 47356
rect 5908 47354 5932 47356
rect 5988 47354 6012 47356
rect 6068 47354 6092 47356
rect 6148 47354 6154 47356
rect 5908 47302 5910 47354
rect 6090 47302 6092 47354
rect 5846 47300 5852 47302
rect 5908 47300 5932 47302
rect 5988 47300 6012 47302
rect 6068 47300 6092 47302
rect 6148 47300 6154 47302
rect 5846 47280 6154 47300
rect 6196 47122 6224 48010
rect 5816 47116 5868 47122
rect 5816 47058 5868 47064
rect 6184 47116 6236 47122
rect 6184 47058 6236 47064
rect 5724 46572 5776 46578
rect 5724 46514 5776 46520
rect 5632 46504 5684 46510
rect 5632 46446 5684 46452
rect 5828 46356 5856 47058
rect 6184 46504 6236 46510
rect 6184 46446 6236 46452
rect 5644 46328 5856 46356
rect 5540 45824 5592 45830
rect 5540 45766 5592 45772
rect 5538 45656 5594 45665
rect 5538 45591 5594 45600
rect 5552 41414 5580 45591
rect 5644 44402 5672 46328
rect 5846 46268 6154 46288
rect 5846 46266 5852 46268
rect 5908 46266 5932 46268
rect 5988 46266 6012 46268
rect 6068 46266 6092 46268
rect 6148 46266 6154 46268
rect 5908 46214 5910 46266
rect 6090 46214 6092 46266
rect 5846 46212 5852 46214
rect 5908 46212 5932 46214
rect 5988 46212 6012 46214
rect 6068 46212 6092 46214
rect 6148 46212 6154 46214
rect 5846 46192 6154 46212
rect 5724 45824 5776 45830
rect 5724 45766 5776 45772
rect 5632 44396 5684 44402
rect 5632 44338 5684 44344
rect 5632 42220 5684 42226
rect 5632 42162 5684 42168
rect 5644 41818 5672 42162
rect 5632 41812 5684 41818
rect 5632 41754 5684 41760
rect 5552 41386 5672 41414
rect 5644 41070 5672 41386
rect 5632 41064 5684 41070
rect 5632 41006 5684 41012
rect 5632 40656 5684 40662
rect 5632 40598 5684 40604
rect 5540 39432 5592 39438
rect 5540 39374 5592 39380
rect 5552 38554 5580 39374
rect 5644 39030 5672 40598
rect 5736 40050 5764 45766
rect 5846 45180 6154 45200
rect 5846 45178 5852 45180
rect 5908 45178 5932 45180
rect 5988 45178 6012 45180
rect 6068 45178 6092 45180
rect 6148 45178 6154 45180
rect 5908 45126 5910 45178
rect 6090 45126 6092 45178
rect 5846 45124 5852 45126
rect 5908 45124 5932 45126
rect 5988 45124 6012 45126
rect 6068 45124 6092 45126
rect 6148 45124 6154 45126
rect 5846 45104 6154 45124
rect 5846 44092 6154 44112
rect 5846 44090 5852 44092
rect 5908 44090 5932 44092
rect 5988 44090 6012 44092
rect 6068 44090 6092 44092
rect 6148 44090 6154 44092
rect 5908 44038 5910 44090
rect 6090 44038 6092 44090
rect 5846 44036 5852 44038
rect 5908 44036 5932 44038
rect 5988 44036 6012 44038
rect 6068 44036 6092 44038
rect 6148 44036 6154 44038
rect 5846 44016 6154 44036
rect 5846 43004 6154 43024
rect 5846 43002 5852 43004
rect 5908 43002 5932 43004
rect 5988 43002 6012 43004
rect 6068 43002 6092 43004
rect 6148 43002 6154 43004
rect 5908 42950 5910 43002
rect 6090 42950 6092 43002
rect 5846 42948 5852 42950
rect 5908 42948 5932 42950
rect 5988 42948 6012 42950
rect 6068 42948 6092 42950
rect 6148 42948 6154 42950
rect 5846 42928 6154 42948
rect 5846 41916 6154 41936
rect 5846 41914 5852 41916
rect 5908 41914 5932 41916
rect 5988 41914 6012 41916
rect 6068 41914 6092 41916
rect 6148 41914 6154 41916
rect 5908 41862 5910 41914
rect 6090 41862 6092 41914
rect 5846 41860 5852 41862
rect 5908 41860 5932 41862
rect 5988 41860 6012 41862
rect 6068 41860 6092 41862
rect 6148 41860 6154 41862
rect 5846 41840 6154 41860
rect 6196 41274 6224 46446
rect 6184 41268 6236 41274
rect 6184 41210 6236 41216
rect 6184 41132 6236 41138
rect 6184 41074 6236 41080
rect 5846 40828 6154 40848
rect 5846 40826 5852 40828
rect 5908 40826 5932 40828
rect 5988 40826 6012 40828
rect 6068 40826 6092 40828
rect 6148 40826 6154 40828
rect 5908 40774 5910 40826
rect 6090 40774 6092 40826
rect 5846 40772 5852 40774
rect 5908 40772 5932 40774
rect 5988 40772 6012 40774
rect 6068 40772 6092 40774
rect 6148 40772 6154 40774
rect 5846 40752 6154 40772
rect 5724 40044 5776 40050
rect 5724 39986 5776 39992
rect 5846 39740 6154 39760
rect 5846 39738 5852 39740
rect 5908 39738 5932 39740
rect 5988 39738 6012 39740
rect 6068 39738 6092 39740
rect 6148 39738 6154 39740
rect 5908 39686 5910 39738
rect 6090 39686 6092 39738
rect 5846 39684 5852 39686
rect 5908 39684 5932 39686
rect 5988 39684 6012 39686
rect 6068 39684 6092 39686
rect 6148 39684 6154 39686
rect 5846 39664 6154 39684
rect 6196 39642 6224 41074
rect 6184 39636 6236 39642
rect 6184 39578 6236 39584
rect 5724 39500 5776 39506
rect 5724 39442 5776 39448
rect 5632 39024 5684 39030
rect 5632 38966 5684 38972
rect 5736 38962 5764 39442
rect 5724 38956 5776 38962
rect 5724 38898 5776 38904
rect 5846 38652 6154 38672
rect 5846 38650 5852 38652
rect 5908 38650 5932 38652
rect 5988 38650 6012 38652
rect 6068 38650 6092 38652
rect 6148 38650 6154 38652
rect 5908 38598 5910 38650
rect 6090 38598 6092 38650
rect 5846 38596 5852 38598
rect 5908 38596 5932 38598
rect 5988 38596 6012 38598
rect 6068 38596 6092 38598
rect 6148 38596 6154 38598
rect 5846 38576 6154 38596
rect 5540 38548 5592 38554
rect 5540 38490 5592 38496
rect 5540 38344 5592 38350
rect 5540 38286 5592 38292
rect 5552 36786 5580 38286
rect 5846 37564 6154 37584
rect 5846 37562 5852 37564
rect 5908 37562 5932 37564
rect 5988 37562 6012 37564
rect 6068 37562 6092 37564
rect 6148 37562 6154 37564
rect 5908 37510 5910 37562
rect 6090 37510 6092 37562
rect 5846 37508 5852 37510
rect 5908 37508 5932 37510
rect 5988 37508 6012 37510
rect 6068 37508 6092 37510
rect 6148 37508 6154 37510
rect 5846 37488 6154 37508
rect 5632 37324 5684 37330
rect 5632 37266 5684 37272
rect 5540 36780 5592 36786
rect 5540 36722 5592 36728
rect 5540 36168 5592 36174
rect 5540 36110 5592 36116
rect 5552 35834 5580 36110
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 5540 33516 5592 33522
rect 5540 33458 5592 33464
rect 5552 31657 5580 33458
rect 5644 32201 5672 37266
rect 5724 36780 5776 36786
rect 5724 36722 5776 36728
rect 5736 35766 5764 36722
rect 5846 36476 6154 36496
rect 5846 36474 5852 36476
rect 5908 36474 5932 36476
rect 5988 36474 6012 36476
rect 6068 36474 6092 36476
rect 6148 36474 6154 36476
rect 5908 36422 5910 36474
rect 6090 36422 6092 36474
rect 5846 36420 5852 36422
rect 5908 36420 5932 36422
rect 5988 36420 6012 36422
rect 6068 36420 6092 36422
rect 6148 36420 6154 36422
rect 5846 36400 6154 36420
rect 5724 35760 5776 35766
rect 5724 35702 5776 35708
rect 5846 35388 6154 35408
rect 5846 35386 5852 35388
rect 5908 35386 5932 35388
rect 5988 35386 6012 35388
rect 6068 35386 6092 35388
rect 6148 35386 6154 35388
rect 5908 35334 5910 35386
rect 6090 35334 6092 35386
rect 5846 35332 5852 35334
rect 5908 35332 5932 35334
rect 5988 35332 6012 35334
rect 6068 35332 6092 35334
rect 6148 35332 6154 35334
rect 5846 35312 6154 35332
rect 5846 34300 6154 34320
rect 5846 34298 5852 34300
rect 5908 34298 5932 34300
rect 5988 34298 6012 34300
rect 6068 34298 6092 34300
rect 6148 34298 6154 34300
rect 5908 34246 5910 34298
rect 6090 34246 6092 34298
rect 5846 34244 5852 34246
rect 5908 34244 5932 34246
rect 5988 34244 6012 34246
rect 6068 34244 6092 34246
rect 6148 34244 6154 34246
rect 5846 34224 6154 34244
rect 5846 33212 6154 33232
rect 5846 33210 5852 33212
rect 5908 33210 5932 33212
rect 5988 33210 6012 33212
rect 6068 33210 6092 33212
rect 6148 33210 6154 33212
rect 5908 33158 5910 33210
rect 6090 33158 6092 33210
rect 5846 33156 5852 33158
rect 5908 33156 5932 33158
rect 5988 33156 6012 33158
rect 6068 33156 6092 33158
rect 6148 33156 6154 33158
rect 5846 33136 6154 33156
rect 5724 32768 5776 32774
rect 5724 32710 5776 32716
rect 5630 32192 5686 32201
rect 5630 32127 5686 32136
rect 5632 31884 5684 31890
rect 5632 31826 5684 31832
rect 5538 31648 5594 31657
rect 5538 31583 5594 31592
rect 5644 31346 5672 31826
rect 5632 31340 5684 31346
rect 5632 31282 5684 31288
rect 5538 31104 5594 31113
rect 5538 31039 5594 31048
rect 5446 28248 5502 28257
rect 5356 28212 5408 28218
rect 5446 28183 5502 28192
rect 5356 28154 5408 28160
rect 5448 28144 5500 28150
rect 5448 28086 5500 28092
rect 5356 28076 5408 28082
rect 5356 28018 5408 28024
rect 5368 16794 5396 28018
rect 5460 26874 5488 28086
rect 5552 27010 5580 31039
rect 5736 30326 5764 32710
rect 5846 32124 6154 32144
rect 5846 32122 5852 32124
rect 5908 32122 5932 32124
rect 5988 32122 6012 32124
rect 6068 32122 6092 32124
rect 6148 32122 6154 32124
rect 5908 32070 5910 32122
rect 6090 32070 6092 32122
rect 5846 32068 5852 32070
rect 5908 32068 5932 32070
rect 5988 32068 6012 32070
rect 6068 32068 6092 32070
rect 6148 32068 6154 32070
rect 5846 32048 6154 32068
rect 5846 31036 6154 31056
rect 5846 31034 5852 31036
rect 5908 31034 5932 31036
rect 5988 31034 6012 31036
rect 6068 31034 6092 31036
rect 6148 31034 6154 31036
rect 5908 30982 5910 31034
rect 6090 30982 6092 31034
rect 5846 30980 5852 30982
rect 5908 30980 5932 30982
rect 5988 30980 6012 30982
rect 6068 30980 6092 30982
rect 6148 30980 6154 30982
rect 5846 30960 6154 30980
rect 5724 30320 5776 30326
rect 5724 30262 5776 30268
rect 5632 30252 5684 30258
rect 5632 30194 5684 30200
rect 5644 27946 5672 30194
rect 5846 29948 6154 29968
rect 5846 29946 5852 29948
rect 5908 29946 5932 29948
rect 5988 29946 6012 29948
rect 6068 29946 6092 29948
rect 6148 29946 6154 29948
rect 5908 29894 5910 29946
rect 6090 29894 6092 29946
rect 5846 29892 5852 29894
rect 5908 29892 5932 29894
rect 5988 29892 6012 29894
rect 6068 29892 6092 29894
rect 6148 29892 6154 29894
rect 5846 29872 6154 29892
rect 5846 28860 6154 28880
rect 5846 28858 5852 28860
rect 5908 28858 5932 28860
rect 5988 28858 6012 28860
rect 6068 28858 6092 28860
rect 6148 28858 6154 28860
rect 5908 28806 5910 28858
rect 6090 28806 6092 28858
rect 5846 28804 5852 28806
rect 5908 28804 5932 28806
rect 5988 28804 6012 28806
rect 6068 28804 6092 28806
rect 6148 28804 6154 28806
rect 5846 28784 6154 28804
rect 5632 27940 5684 27946
rect 5632 27882 5684 27888
rect 5846 27772 6154 27792
rect 5846 27770 5852 27772
rect 5908 27770 5932 27772
rect 5988 27770 6012 27772
rect 6068 27770 6092 27772
rect 6148 27770 6154 27772
rect 5908 27718 5910 27770
rect 6090 27718 6092 27770
rect 5846 27716 5852 27718
rect 5908 27716 5932 27718
rect 5988 27716 6012 27718
rect 6068 27716 6092 27718
rect 6148 27716 6154 27718
rect 5846 27696 6154 27716
rect 5552 26982 5672 27010
rect 5460 26846 5580 26874
rect 5448 26784 5500 26790
rect 5448 26726 5500 26732
rect 5460 19378 5488 26726
rect 5552 26586 5580 26846
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 5644 26518 5672 26982
rect 5846 26684 6154 26704
rect 5846 26682 5852 26684
rect 5908 26682 5932 26684
rect 5988 26682 6012 26684
rect 6068 26682 6092 26684
rect 6148 26682 6154 26684
rect 5908 26630 5910 26682
rect 6090 26630 6092 26682
rect 5846 26628 5852 26630
rect 5908 26628 5932 26630
rect 5988 26628 6012 26630
rect 6068 26628 6092 26630
rect 6148 26628 6154 26630
rect 5846 26608 6154 26628
rect 5632 26512 5684 26518
rect 5632 26454 5684 26460
rect 6288 26450 6316 54606
rect 6380 28626 6408 56238
rect 6460 55684 6512 55690
rect 6460 55626 6512 55632
rect 6472 28762 6500 55626
rect 6564 49881 6592 57394
rect 8312 56914 8340 59366
rect 8496 59090 8524 63174
rect 9110 62588 9418 62608
rect 9110 62586 9116 62588
rect 9172 62586 9196 62588
rect 9252 62586 9276 62588
rect 9332 62586 9356 62588
rect 9412 62586 9418 62588
rect 9172 62534 9174 62586
rect 9354 62534 9356 62586
rect 9110 62532 9116 62534
rect 9172 62532 9196 62534
rect 9252 62532 9276 62534
rect 9332 62532 9356 62534
rect 9412 62532 9418 62534
rect 9110 62512 9418 62532
rect 9110 61500 9418 61520
rect 9110 61498 9116 61500
rect 9172 61498 9196 61500
rect 9252 61498 9276 61500
rect 9332 61498 9356 61500
rect 9412 61498 9418 61500
rect 9172 61446 9174 61498
rect 9354 61446 9356 61498
rect 9110 61444 9116 61446
rect 9172 61444 9196 61446
rect 9252 61444 9276 61446
rect 9332 61444 9356 61446
rect 9412 61444 9418 61446
rect 9110 61424 9418 61444
rect 9110 60412 9418 60432
rect 9110 60410 9116 60412
rect 9172 60410 9196 60412
rect 9252 60410 9276 60412
rect 9332 60410 9356 60412
rect 9412 60410 9418 60412
rect 9172 60358 9174 60410
rect 9354 60358 9356 60410
rect 9110 60356 9116 60358
rect 9172 60356 9196 60358
rect 9252 60356 9276 60358
rect 9332 60356 9356 60358
rect 9412 60356 9418 60358
rect 9110 60336 9418 60356
rect 9110 59324 9418 59344
rect 9110 59322 9116 59324
rect 9172 59322 9196 59324
rect 9252 59322 9276 59324
rect 9332 59322 9356 59324
rect 9412 59322 9418 59324
rect 9172 59270 9174 59322
rect 9354 59270 9356 59322
rect 9110 59268 9116 59270
rect 9172 59268 9196 59270
rect 9252 59268 9276 59270
rect 9332 59268 9356 59270
rect 9412 59268 9418 59270
rect 9110 59248 9418 59268
rect 8484 59084 8536 59090
rect 8484 59026 8536 59032
rect 9496 58472 9548 58478
rect 9496 58414 9548 58420
rect 9110 58236 9418 58256
rect 9110 58234 9116 58236
rect 9172 58234 9196 58236
rect 9252 58234 9276 58236
rect 9332 58234 9356 58236
rect 9412 58234 9418 58236
rect 9172 58182 9174 58234
rect 9354 58182 9356 58234
rect 9110 58180 9116 58182
rect 9172 58180 9196 58182
rect 9252 58180 9276 58182
rect 9332 58180 9356 58182
rect 9412 58180 9418 58182
rect 9110 58160 9418 58180
rect 9508 58041 9536 58414
rect 9494 58032 9550 58041
rect 9494 57967 9550 57976
rect 9496 57384 9548 57390
rect 9496 57326 9548 57332
rect 9508 57225 9536 57326
rect 9494 57216 9550 57225
rect 9110 57148 9418 57168
rect 9494 57151 9550 57160
rect 9110 57146 9116 57148
rect 9172 57146 9196 57148
rect 9252 57146 9276 57148
rect 9332 57146 9356 57148
rect 9412 57146 9418 57148
rect 9172 57094 9174 57146
rect 9354 57094 9356 57146
rect 9110 57092 9116 57094
rect 9172 57092 9196 57094
rect 9252 57092 9276 57094
rect 9332 57092 9356 57094
rect 9412 57092 9418 57094
rect 9110 57072 9418 57092
rect 8300 56908 8352 56914
rect 8300 56850 8352 56856
rect 8484 56908 8536 56914
rect 8484 56850 8536 56856
rect 7478 56604 7786 56624
rect 7478 56602 7484 56604
rect 7540 56602 7564 56604
rect 7620 56602 7644 56604
rect 7700 56602 7724 56604
rect 7780 56602 7786 56604
rect 7540 56550 7542 56602
rect 7722 56550 7724 56602
rect 7478 56548 7484 56550
rect 7540 56548 7564 56550
rect 7620 56548 7644 56550
rect 7700 56548 7724 56550
rect 7780 56548 7786 56550
rect 7478 56528 7786 56548
rect 6828 55616 6880 55622
rect 6828 55558 6880 55564
rect 8300 55616 8352 55622
rect 8300 55558 8352 55564
rect 6840 54670 6868 55558
rect 7478 55516 7786 55536
rect 7478 55514 7484 55516
rect 7540 55514 7564 55516
rect 7620 55514 7644 55516
rect 7700 55514 7724 55516
rect 7780 55514 7786 55516
rect 7540 55462 7542 55514
rect 7722 55462 7724 55514
rect 7478 55460 7484 55462
rect 7540 55460 7564 55462
rect 7620 55460 7644 55462
rect 7700 55460 7724 55462
rect 7780 55460 7786 55462
rect 7478 55440 7786 55460
rect 6828 54664 6880 54670
rect 6828 54606 6880 54612
rect 7478 54428 7786 54448
rect 7478 54426 7484 54428
rect 7540 54426 7564 54428
rect 7620 54426 7644 54428
rect 7700 54426 7724 54428
rect 7780 54426 7786 54428
rect 7540 54374 7542 54426
rect 7722 54374 7724 54426
rect 7478 54372 7484 54374
rect 7540 54372 7564 54374
rect 7620 54372 7644 54374
rect 7700 54372 7724 54374
rect 7780 54372 7786 54374
rect 7478 54352 7786 54372
rect 8312 54262 8340 55558
rect 8300 54256 8352 54262
rect 8300 54198 8352 54204
rect 7478 53340 7786 53360
rect 7478 53338 7484 53340
rect 7540 53338 7564 53340
rect 7620 53338 7644 53340
rect 7700 53338 7724 53340
rect 7780 53338 7786 53340
rect 7540 53286 7542 53338
rect 7722 53286 7724 53338
rect 7478 53284 7484 53286
rect 7540 53284 7564 53286
rect 7620 53284 7644 53286
rect 7700 53284 7724 53286
rect 7780 53284 7786 53286
rect 7478 53264 7786 53284
rect 6828 53168 6880 53174
rect 6828 53110 6880 53116
rect 6644 51264 6696 51270
rect 6644 51206 6696 51212
rect 6656 50862 6684 51206
rect 6644 50856 6696 50862
rect 6644 50798 6696 50804
rect 6550 49872 6606 49881
rect 6550 49807 6606 49816
rect 6552 49224 6604 49230
rect 6552 49166 6604 49172
rect 6564 48550 6592 49166
rect 6736 49156 6788 49162
rect 6736 49098 6788 49104
rect 6552 48544 6604 48550
rect 6552 48486 6604 48492
rect 6552 46572 6604 46578
rect 6552 46514 6604 46520
rect 6564 40746 6592 46514
rect 6644 46368 6696 46374
rect 6644 46310 6696 46316
rect 6656 41154 6684 46310
rect 6748 41313 6776 49098
rect 6734 41304 6790 41313
rect 6734 41239 6790 41248
rect 6656 41126 6776 41154
rect 6564 40718 6684 40746
rect 6656 40118 6684 40718
rect 6644 40112 6696 40118
rect 6644 40054 6696 40060
rect 6552 40044 6604 40050
rect 6552 39986 6604 39992
rect 6564 39098 6592 39986
rect 6552 39092 6604 39098
rect 6552 39034 6604 39040
rect 6748 37874 6776 41126
rect 6736 37868 6788 37874
rect 6736 37810 6788 37816
rect 6840 36378 6868 53110
rect 7478 52252 7786 52272
rect 7478 52250 7484 52252
rect 7540 52250 7564 52252
rect 7620 52250 7644 52252
rect 7700 52250 7724 52252
rect 7780 52250 7786 52252
rect 7540 52198 7542 52250
rect 7722 52198 7724 52250
rect 7478 52196 7484 52198
rect 7540 52196 7564 52198
rect 7620 52196 7644 52198
rect 7700 52196 7724 52198
rect 7780 52196 7786 52198
rect 7478 52176 7786 52196
rect 6920 51944 6972 51950
rect 6920 51886 6972 51892
rect 6828 36372 6880 36378
rect 6828 36314 6880 36320
rect 6932 29646 6960 51886
rect 7478 51164 7786 51184
rect 7478 51162 7484 51164
rect 7540 51162 7564 51164
rect 7620 51162 7644 51164
rect 7700 51162 7724 51164
rect 7780 51162 7786 51164
rect 7540 51110 7542 51162
rect 7722 51110 7724 51162
rect 7478 51108 7484 51110
rect 7540 51108 7564 51110
rect 7620 51108 7644 51110
rect 7700 51108 7724 51110
rect 7780 51108 7786 51110
rect 7478 51088 7786 51108
rect 8496 50386 8524 56850
rect 9312 56840 9364 56846
rect 9312 56782 9364 56788
rect 9324 56409 9352 56782
rect 9310 56400 9366 56409
rect 9310 56335 9366 56344
rect 9110 56060 9418 56080
rect 9110 56058 9116 56060
rect 9172 56058 9196 56060
rect 9252 56058 9276 56060
rect 9332 56058 9356 56060
rect 9412 56058 9418 56060
rect 9172 56006 9174 56058
rect 9354 56006 9356 56058
rect 9110 56004 9116 56006
rect 9172 56004 9196 56006
rect 9252 56004 9276 56006
rect 9332 56004 9356 56006
rect 9412 56004 9418 56006
rect 9110 55984 9418 56004
rect 9588 55752 9640 55758
rect 9588 55694 9640 55700
rect 9110 54972 9418 54992
rect 9110 54970 9116 54972
rect 9172 54970 9196 54972
rect 9252 54970 9276 54972
rect 9332 54970 9356 54972
rect 9412 54970 9418 54972
rect 9172 54918 9174 54970
rect 9354 54918 9356 54970
rect 9110 54916 9116 54918
rect 9172 54916 9196 54918
rect 9252 54916 9276 54918
rect 9332 54916 9356 54918
rect 9412 54916 9418 54918
rect 9110 54896 9418 54916
rect 9600 54913 9628 55694
rect 9586 54904 9642 54913
rect 9586 54839 9642 54848
rect 9680 54528 9732 54534
rect 9680 54470 9732 54476
rect 9110 53884 9418 53904
rect 9110 53882 9116 53884
rect 9172 53882 9196 53884
rect 9252 53882 9276 53884
rect 9332 53882 9356 53884
rect 9412 53882 9418 53884
rect 9172 53830 9174 53882
rect 9354 53830 9356 53882
rect 9110 53828 9116 53830
rect 9172 53828 9196 53830
rect 9252 53828 9276 53830
rect 9332 53828 9356 53830
rect 9412 53828 9418 53830
rect 9110 53808 9418 53828
rect 9692 53582 9720 54470
rect 9680 53576 9732 53582
rect 9680 53518 9732 53524
rect 9110 52796 9418 52816
rect 9110 52794 9116 52796
rect 9172 52794 9196 52796
rect 9252 52794 9276 52796
rect 9332 52794 9356 52796
rect 9412 52794 9418 52796
rect 9172 52742 9174 52794
rect 9354 52742 9356 52794
rect 9110 52740 9116 52742
rect 9172 52740 9196 52742
rect 9252 52740 9276 52742
rect 9332 52740 9356 52742
rect 9412 52740 9418 52742
rect 9110 52720 9418 52740
rect 9110 51708 9418 51728
rect 9110 51706 9116 51708
rect 9172 51706 9196 51708
rect 9252 51706 9276 51708
rect 9332 51706 9356 51708
rect 9412 51706 9418 51708
rect 9172 51654 9174 51706
rect 9354 51654 9356 51706
rect 9110 51652 9116 51654
rect 9172 51652 9196 51654
rect 9252 51652 9276 51654
rect 9332 51652 9356 51654
rect 9412 51652 9418 51654
rect 9110 51632 9418 51652
rect 9680 51400 9732 51406
rect 9680 51342 9732 51348
rect 9110 50620 9418 50640
rect 9110 50618 9116 50620
rect 9172 50618 9196 50620
rect 9252 50618 9276 50620
rect 9332 50618 9356 50620
rect 9412 50618 9418 50620
rect 9172 50566 9174 50618
rect 9354 50566 9356 50618
rect 9110 50564 9116 50566
rect 9172 50564 9196 50566
rect 9252 50564 9276 50566
rect 9332 50564 9356 50566
rect 9412 50564 9418 50566
rect 9110 50544 9418 50564
rect 8484 50380 8536 50386
rect 8484 50322 8536 50328
rect 7104 50312 7156 50318
rect 7104 50254 7156 50260
rect 7012 46572 7064 46578
rect 7012 46514 7064 46520
rect 7024 45082 7052 46514
rect 7012 45076 7064 45082
rect 7012 45018 7064 45024
rect 7116 37330 7144 50254
rect 7478 50076 7786 50096
rect 7478 50074 7484 50076
rect 7540 50074 7564 50076
rect 7620 50074 7644 50076
rect 7700 50074 7724 50076
rect 7780 50074 7786 50076
rect 7540 50022 7542 50074
rect 7722 50022 7724 50074
rect 7478 50020 7484 50022
rect 7540 50020 7564 50022
rect 7620 50020 7644 50022
rect 7700 50020 7724 50022
rect 7780 50020 7786 50022
rect 7478 50000 7786 50020
rect 9588 49972 9640 49978
rect 9588 49914 9640 49920
rect 9110 49532 9418 49552
rect 9110 49530 9116 49532
rect 9172 49530 9196 49532
rect 9252 49530 9276 49532
rect 9332 49530 9356 49532
rect 9412 49530 9418 49532
rect 9172 49478 9174 49530
rect 9354 49478 9356 49530
rect 9110 49476 9116 49478
rect 9172 49476 9196 49478
rect 9252 49476 9276 49478
rect 9332 49476 9356 49478
rect 9412 49476 9418 49478
rect 9110 49456 9418 49476
rect 9600 49473 9628 49914
rect 9586 49464 9642 49473
rect 9692 49434 9720 51342
rect 9586 49399 9642 49408
rect 9680 49428 9732 49434
rect 9680 49370 9732 49376
rect 9496 49224 9548 49230
rect 9496 49166 9548 49172
rect 7478 48988 7786 49008
rect 7478 48986 7484 48988
rect 7540 48986 7564 48988
rect 7620 48986 7644 48988
rect 7700 48986 7724 48988
rect 7780 48986 7786 48988
rect 7540 48934 7542 48986
rect 7722 48934 7724 48986
rect 7478 48932 7484 48934
rect 7540 48932 7564 48934
rect 7620 48932 7644 48934
rect 7700 48932 7724 48934
rect 7780 48932 7786 48934
rect 7478 48912 7786 48932
rect 9110 48444 9418 48464
rect 9110 48442 9116 48444
rect 9172 48442 9196 48444
rect 9252 48442 9276 48444
rect 9332 48442 9356 48444
rect 9412 48442 9418 48444
rect 9172 48390 9174 48442
rect 9354 48390 9356 48442
rect 9110 48388 9116 48390
rect 9172 48388 9196 48390
rect 9252 48388 9276 48390
rect 9332 48388 9356 48390
rect 9412 48388 9418 48390
rect 9110 48368 9418 48388
rect 9508 48278 9536 49166
rect 7196 48272 7248 48278
rect 7196 48214 7248 48220
rect 9496 48272 9548 48278
rect 9496 48214 9548 48220
rect 7104 37324 7156 37330
rect 7104 37266 7156 37272
rect 6920 29640 6972 29646
rect 6920 29582 6972 29588
rect 6460 28756 6512 28762
rect 6460 28698 6512 28704
rect 6368 28620 6420 28626
rect 6368 28562 6420 28568
rect 7208 28014 7236 48214
rect 7478 47900 7786 47920
rect 7478 47898 7484 47900
rect 7540 47898 7564 47900
rect 7620 47898 7644 47900
rect 7700 47898 7724 47900
rect 7780 47898 7786 47900
rect 7540 47846 7542 47898
rect 7722 47846 7724 47898
rect 7478 47844 7484 47846
rect 7540 47844 7564 47846
rect 7620 47844 7644 47846
rect 7700 47844 7724 47846
rect 7780 47844 7786 47846
rect 7478 47824 7786 47844
rect 7472 47660 7524 47666
rect 7472 47602 7524 47608
rect 7484 47258 7512 47602
rect 9110 47356 9418 47376
rect 9110 47354 9116 47356
rect 9172 47354 9196 47356
rect 9252 47354 9276 47356
rect 9332 47354 9356 47356
rect 9412 47354 9418 47356
rect 9172 47302 9174 47354
rect 9354 47302 9356 47354
rect 9110 47300 9116 47302
rect 9172 47300 9196 47302
rect 9252 47300 9276 47302
rect 9332 47300 9356 47302
rect 9412 47300 9418 47302
rect 9110 47280 9418 47300
rect 7288 47252 7340 47258
rect 7288 47194 7340 47200
rect 7472 47252 7524 47258
rect 7472 47194 7524 47200
rect 7300 40934 7328 47194
rect 7478 46812 7786 46832
rect 7478 46810 7484 46812
rect 7540 46810 7564 46812
rect 7620 46810 7644 46812
rect 7700 46810 7724 46812
rect 7780 46810 7786 46812
rect 7540 46758 7542 46810
rect 7722 46758 7724 46810
rect 7478 46756 7484 46758
rect 7540 46756 7564 46758
rect 7620 46756 7644 46758
rect 7700 46756 7724 46758
rect 7780 46756 7786 46758
rect 7478 46736 7786 46756
rect 9110 46268 9418 46288
rect 9110 46266 9116 46268
rect 9172 46266 9196 46268
rect 9252 46266 9276 46268
rect 9332 46266 9356 46268
rect 9412 46266 9418 46268
rect 9172 46214 9174 46266
rect 9354 46214 9356 46266
rect 9110 46212 9116 46214
rect 9172 46212 9196 46214
rect 9252 46212 9276 46214
rect 9332 46212 9356 46214
rect 9412 46212 9418 46214
rect 9110 46192 9418 46212
rect 7478 45724 7786 45744
rect 7478 45722 7484 45724
rect 7540 45722 7564 45724
rect 7620 45722 7644 45724
rect 7700 45722 7724 45724
rect 7780 45722 7786 45724
rect 7540 45670 7542 45722
rect 7722 45670 7724 45722
rect 7478 45668 7484 45670
rect 7540 45668 7564 45670
rect 7620 45668 7644 45670
rect 7700 45668 7724 45670
rect 7780 45668 7786 45670
rect 7478 45648 7786 45668
rect 9110 45180 9418 45200
rect 9110 45178 9116 45180
rect 9172 45178 9196 45180
rect 9252 45178 9276 45180
rect 9332 45178 9356 45180
rect 9412 45178 9418 45180
rect 9172 45126 9174 45178
rect 9354 45126 9356 45178
rect 9110 45124 9116 45126
rect 9172 45124 9196 45126
rect 9252 45124 9276 45126
rect 9332 45124 9356 45126
rect 9412 45124 9418 45126
rect 9110 45104 9418 45124
rect 8300 44872 8352 44878
rect 8300 44814 8352 44820
rect 7478 44636 7786 44656
rect 7478 44634 7484 44636
rect 7540 44634 7564 44636
rect 7620 44634 7644 44636
rect 7700 44634 7724 44636
rect 7780 44634 7786 44636
rect 7540 44582 7542 44634
rect 7722 44582 7724 44634
rect 7478 44580 7484 44582
rect 7540 44580 7564 44582
rect 7620 44580 7644 44582
rect 7700 44580 7724 44582
rect 7780 44580 7786 44582
rect 7478 44560 7786 44580
rect 7478 43548 7786 43568
rect 7478 43546 7484 43548
rect 7540 43546 7564 43548
rect 7620 43546 7644 43548
rect 7700 43546 7724 43548
rect 7780 43546 7786 43548
rect 7540 43494 7542 43546
rect 7722 43494 7724 43546
rect 7478 43492 7484 43494
rect 7540 43492 7564 43494
rect 7620 43492 7644 43494
rect 7700 43492 7724 43494
rect 7780 43492 7786 43494
rect 7478 43472 7786 43492
rect 7478 42460 7786 42480
rect 7478 42458 7484 42460
rect 7540 42458 7564 42460
rect 7620 42458 7644 42460
rect 7700 42458 7724 42460
rect 7780 42458 7786 42460
rect 7540 42406 7542 42458
rect 7722 42406 7724 42458
rect 7478 42404 7484 42406
rect 7540 42404 7564 42406
rect 7620 42404 7644 42406
rect 7700 42404 7724 42406
rect 7780 42404 7786 42406
rect 7478 42384 7786 42404
rect 8312 42090 8340 44814
rect 9496 44396 9548 44402
rect 9496 44338 9548 44344
rect 9110 44092 9418 44112
rect 9110 44090 9116 44092
rect 9172 44090 9196 44092
rect 9252 44090 9276 44092
rect 9332 44090 9356 44092
rect 9412 44090 9418 44092
rect 9172 44038 9174 44090
rect 9354 44038 9356 44090
rect 9110 44036 9116 44038
rect 9172 44036 9196 44038
rect 9252 44036 9276 44038
rect 9332 44036 9356 44038
rect 9412 44036 9418 44038
rect 9110 44016 9418 44036
rect 9508 43994 9536 44338
rect 9496 43988 9548 43994
rect 9496 43930 9548 43936
rect 9784 43926 9812 76774
rect 10140 76424 10192 76430
rect 10138 76392 10140 76401
rect 10192 76392 10194 76401
rect 10138 76327 10194 76336
rect 10140 75948 10192 75954
rect 10140 75890 10192 75896
rect 10152 75721 10180 75890
rect 10138 75712 10194 75721
rect 10138 75647 10194 75656
rect 10140 75336 10192 75342
rect 10140 75278 10192 75284
rect 10152 74905 10180 75278
rect 10138 74896 10194 74905
rect 10138 74831 10194 74840
rect 10140 74248 10192 74254
rect 10140 74190 10192 74196
rect 10152 74089 10180 74190
rect 10138 74080 10194 74089
rect 10138 74015 10194 74024
rect 10140 73772 10192 73778
rect 10140 73714 10192 73720
rect 10152 73409 10180 73714
rect 10138 73400 10194 73409
rect 10138 73335 10194 73344
rect 10140 72684 10192 72690
rect 10140 72626 10192 72632
rect 9956 72616 10008 72622
rect 10152 72593 10180 72626
rect 9956 72558 10008 72564
rect 10138 72584 10194 72593
rect 9968 72282 9996 72558
rect 10138 72519 10194 72528
rect 9956 72276 10008 72282
rect 9956 72218 10008 72224
rect 10140 72072 10192 72078
rect 10140 72014 10192 72020
rect 10152 71777 10180 72014
rect 10138 71768 10194 71777
rect 10138 71703 10194 71712
rect 10140 71596 10192 71602
rect 10140 71538 10192 71544
rect 10152 71097 10180 71538
rect 10138 71088 10194 71097
rect 10138 71023 10194 71032
rect 10140 70508 10192 70514
rect 10140 70450 10192 70456
rect 10152 70281 10180 70450
rect 10138 70272 10194 70281
rect 10138 70207 10194 70216
rect 10140 69896 10192 69902
rect 10140 69838 10192 69844
rect 9956 69760 10008 69766
rect 9956 69702 10008 69708
rect 9968 69358 9996 69702
rect 10152 69465 10180 69838
rect 10138 69456 10194 69465
rect 10138 69391 10194 69400
rect 9956 69352 10008 69358
rect 9956 69294 10008 69300
rect 10140 68808 10192 68814
rect 10138 68776 10140 68785
rect 10192 68776 10194 68785
rect 10138 68711 10194 68720
rect 10140 68332 10192 68338
rect 10140 68274 10192 68280
rect 10152 67969 10180 68274
rect 10138 67960 10194 67969
rect 10138 67895 10194 67904
rect 10140 67244 10192 67250
rect 10140 67186 10192 67192
rect 10152 67153 10180 67186
rect 10138 67144 10194 67153
rect 10138 67079 10194 67088
rect 10140 66632 10192 66638
rect 10140 66574 10192 66580
rect 10152 66473 10180 66574
rect 10138 66464 10194 66473
rect 10138 66399 10194 66408
rect 10140 66156 10192 66162
rect 10140 66098 10192 66104
rect 9956 65952 10008 65958
rect 9956 65894 10008 65900
rect 9968 65618 9996 65894
rect 10152 65657 10180 66098
rect 10138 65648 10194 65657
rect 9956 65612 10008 65618
rect 10138 65583 10194 65592
rect 9956 65554 10008 65560
rect 10140 65068 10192 65074
rect 10140 65010 10192 65016
rect 10152 64841 10180 65010
rect 10138 64832 10194 64841
rect 10138 64767 10194 64776
rect 10140 64456 10192 64462
rect 10140 64398 10192 64404
rect 10152 64161 10180 64398
rect 10138 64152 10194 64161
rect 10138 64087 10194 64096
rect 10140 63368 10192 63374
rect 10138 63336 10140 63345
rect 10192 63336 10194 63345
rect 10138 63271 10194 63280
rect 10140 62892 10192 62898
rect 10140 62834 10192 62840
rect 10152 62529 10180 62834
rect 10138 62520 10194 62529
rect 10138 62455 10194 62464
rect 10140 62280 10192 62286
rect 10140 62222 10192 62228
rect 9956 61872 10008 61878
rect 10152 61849 10180 62222
rect 9956 61814 10008 61820
rect 10138 61840 10194 61849
rect 9968 61402 9996 61814
rect 10138 61775 10194 61784
rect 9956 61396 10008 61402
rect 9956 61338 10008 61344
rect 10140 61192 10192 61198
rect 10140 61134 10192 61140
rect 10152 61033 10180 61134
rect 10138 61024 10194 61033
rect 10138 60959 10194 60968
rect 10140 60716 10192 60722
rect 10140 60658 10192 60664
rect 9956 60512 10008 60518
rect 9956 60454 10008 60460
rect 9968 59566 9996 60454
rect 10152 60353 10180 60658
rect 10138 60344 10194 60353
rect 10138 60279 10194 60288
rect 10140 59628 10192 59634
rect 10140 59570 10192 59576
rect 9956 59560 10008 59566
rect 10152 59537 10180 59570
rect 9956 59502 10008 59508
rect 10138 59528 10194 59537
rect 10138 59463 10194 59472
rect 10140 59016 10192 59022
rect 10140 58958 10192 58964
rect 9956 58880 10008 58886
rect 9956 58822 10008 58828
rect 9968 57322 9996 58822
rect 10152 58721 10180 58958
rect 10138 58712 10194 58721
rect 10138 58647 10194 58656
rect 9956 57316 10008 57322
rect 9956 57258 10008 57264
rect 10140 56364 10192 56370
rect 10140 56306 10192 56312
rect 10152 55729 10180 56306
rect 10138 55720 10194 55729
rect 10138 55655 10194 55664
rect 10140 55412 10192 55418
rect 10140 55354 10192 55360
rect 9864 55072 9916 55078
rect 9864 55014 9916 55020
rect 9876 54194 9904 55014
rect 10152 54670 10180 55354
rect 10140 54664 10192 54670
rect 10140 54606 10192 54612
rect 9956 54528 10008 54534
rect 9956 54470 10008 54476
rect 9864 54188 9916 54194
rect 9864 54130 9916 54136
rect 9968 53106 9996 54470
rect 10046 54088 10102 54097
rect 10046 54023 10048 54032
rect 10100 54023 10102 54032
rect 10048 53994 10100 54000
rect 10048 53440 10100 53446
rect 10046 53408 10048 53417
rect 10100 53408 10102 53417
rect 10046 53343 10102 53352
rect 9956 53100 10008 53106
rect 9956 53042 10008 53048
rect 10048 52896 10100 52902
rect 10048 52838 10100 52844
rect 10060 52601 10088 52838
rect 10046 52592 10102 52601
rect 10046 52527 10102 52536
rect 9864 52012 9916 52018
rect 9864 51954 9916 51960
rect 9876 51066 9904 51954
rect 10048 51808 10100 51814
rect 10046 51776 10048 51785
rect 10100 51776 10102 51785
rect 10046 51711 10102 51720
rect 10048 51264 10100 51270
rect 10048 51206 10100 51212
rect 10060 51105 10088 51206
rect 10046 51096 10102 51105
rect 9864 51060 9916 51066
rect 10046 51031 10102 51040
rect 9864 51002 9916 51008
rect 9864 50312 9916 50318
rect 9864 50254 9916 50260
rect 10046 50280 10102 50289
rect 9876 48890 9904 50254
rect 10046 50215 10102 50224
rect 10060 50182 10088 50215
rect 10048 50176 10100 50182
rect 10048 50118 10100 50124
rect 9956 49836 10008 49842
rect 9956 49778 10008 49784
rect 9864 48884 9916 48890
rect 9864 48826 9916 48832
rect 9968 47258 9996 49778
rect 10048 49088 10100 49094
rect 10048 49030 10100 49036
rect 10060 48793 10088 49030
rect 10046 48784 10102 48793
rect 10046 48719 10102 48728
rect 10140 48748 10192 48754
rect 10140 48690 10192 48696
rect 10048 48000 10100 48006
rect 10046 47968 10048 47977
rect 10100 47968 10102 47977
rect 10046 47903 10102 47912
rect 10048 47456 10100 47462
rect 10048 47398 10100 47404
rect 9956 47252 10008 47258
rect 9956 47194 10008 47200
rect 10060 47161 10088 47398
rect 10046 47152 10102 47161
rect 10046 47087 10102 47096
rect 10152 46714 10180 48690
rect 10140 46708 10192 46714
rect 10140 46650 10192 46656
rect 10046 46472 10102 46481
rect 10046 46407 10048 46416
rect 10100 46407 10102 46416
rect 10048 46378 10100 46384
rect 9864 45960 9916 45966
rect 9864 45902 9916 45908
rect 9772 43920 9824 43926
rect 9772 43862 9824 43868
rect 9110 43004 9418 43024
rect 9110 43002 9116 43004
rect 9172 43002 9196 43004
rect 9252 43002 9276 43004
rect 9332 43002 9356 43004
rect 9412 43002 9418 43004
rect 9172 42950 9174 43002
rect 9354 42950 9356 43002
rect 9110 42948 9116 42950
rect 9172 42948 9196 42950
rect 9252 42948 9276 42950
rect 9332 42948 9356 42950
rect 9412 42948 9418 42950
rect 9110 42928 9418 42948
rect 9772 42696 9824 42702
rect 9772 42638 9824 42644
rect 9496 42220 9548 42226
rect 9496 42162 9548 42168
rect 8300 42084 8352 42090
rect 8300 42026 8352 42032
rect 9110 41916 9418 41936
rect 9110 41914 9116 41916
rect 9172 41914 9196 41916
rect 9252 41914 9276 41916
rect 9332 41914 9356 41916
rect 9412 41914 9418 41916
rect 9172 41862 9174 41914
rect 9354 41862 9356 41914
rect 9110 41860 9116 41862
rect 9172 41860 9196 41862
rect 9252 41860 9276 41862
rect 9332 41860 9356 41862
rect 9412 41860 9418 41862
rect 9110 41840 9418 41860
rect 7478 41372 7786 41392
rect 7478 41370 7484 41372
rect 7540 41370 7564 41372
rect 7620 41370 7644 41372
rect 7700 41370 7724 41372
rect 7780 41370 7786 41372
rect 7540 41318 7542 41370
rect 7722 41318 7724 41370
rect 7478 41316 7484 41318
rect 7540 41316 7564 41318
rect 7620 41316 7644 41318
rect 7700 41316 7724 41318
rect 7780 41316 7786 41318
rect 7478 41296 7786 41316
rect 7288 40928 7340 40934
rect 7288 40870 7340 40876
rect 9110 40828 9418 40848
rect 9110 40826 9116 40828
rect 9172 40826 9196 40828
rect 9252 40826 9276 40828
rect 9332 40826 9356 40828
rect 9412 40826 9418 40828
rect 9172 40774 9174 40826
rect 9354 40774 9356 40826
rect 9110 40772 9116 40774
rect 9172 40772 9196 40774
rect 9252 40772 9276 40774
rect 9332 40772 9356 40774
rect 9412 40772 9418 40774
rect 9110 40752 9418 40772
rect 9508 40730 9536 42162
rect 9496 40724 9548 40730
rect 9496 40666 9548 40672
rect 7478 40284 7786 40304
rect 7478 40282 7484 40284
rect 7540 40282 7564 40284
rect 7620 40282 7644 40284
rect 7700 40282 7724 40284
rect 7780 40282 7786 40284
rect 7540 40230 7542 40282
rect 7722 40230 7724 40282
rect 7478 40228 7484 40230
rect 7540 40228 7564 40230
rect 7620 40228 7644 40230
rect 7700 40228 7724 40230
rect 7780 40228 7786 40230
rect 7478 40208 7786 40228
rect 9110 39740 9418 39760
rect 9110 39738 9116 39740
rect 9172 39738 9196 39740
rect 9252 39738 9276 39740
rect 9332 39738 9356 39740
rect 9412 39738 9418 39740
rect 9172 39686 9174 39738
rect 9354 39686 9356 39738
rect 9110 39684 9116 39686
rect 9172 39684 9196 39686
rect 9252 39684 9276 39686
rect 9332 39684 9356 39686
rect 9412 39684 9418 39686
rect 9110 39664 9418 39684
rect 9784 39642 9812 42638
rect 9876 41002 9904 45902
rect 10048 45824 10100 45830
rect 10048 45766 10100 45772
rect 10060 45665 10088 45766
rect 10046 45656 10102 45665
rect 10046 45591 10102 45600
rect 10046 44840 10102 44849
rect 10046 44775 10102 44784
rect 10060 44742 10088 44775
rect 10048 44736 10100 44742
rect 10048 44678 10100 44684
rect 10048 44192 10100 44198
rect 10046 44160 10048 44169
rect 10100 44160 10102 44169
rect 10046 44095 10102 44104
rect 9956 43784 10008 43790
rect 9956 43726 10008 43732
rect 9968 43450 9996 43726
rect 10048 43648 10100 43654
rect 10048 43590 10100 43596
rect 9956 43444 10008 43450
rect 9956 43386 10008 43392
rect 10060 43353 10088 43590
rect 10046 43344 10102 43353
rect 10046 43279 10102 43288
rect 10140 43308 10192 43314
rect 10140 43250 10192 43256
rect 10048 42560 10100 42566
rect 10046 42528 10048 42537
rect 10100 42528 10102 42537
rect 10046 42463 10102 42472
rect 10152 42362 10180 43250
rect 10140 42356 10192 42362
rect 10140 42298 10192 42304
rect 10048 42016 10100 42022
rect 10048 41958 10100 41964
rect 10060 41857 10088 41958
rect 10046 41848 10102 41857
rect 10046 41783 10102 41792
rect 10046 41032 10102 41041
rect 9864 40996 9916 41002
rect 10046 40967 10048 40976
rect 9864 40938 9916 40944
rect 10100 40967 10102 40976
rect 10048 40938 10100 40944
rect 9864 40520 9916 40526
rect 9864 40462 9916 40468
rect 9876 40186 9904 40462
rect 10048 40384 10100 40390
rect 10046 40352 10048 40361
rect 10100 40352 10102 40361
rect 10046 40287 10102 40296
rect 9864 40180 9916 40186
rect 9864 40122 9916 40128
rect 9864 40044 9916 40050
rect 9864 39986 9916 39992
rect 9772 39636 9824 39642
rect 9772 39578 9824 39584
rect 7478 39196 7786 39216
rect 7478 39194 7484 39196
rect 7540 39194 7564 39196
rect 7620 39194 7644 39196
rect 7700 39194 7724 39196
rect 7780 39194 7786 39196
rect 7540 39142 7542 39194
rect 7722 39142 7724 39194
rect 7478 39140 7484 39142
rect 7540 39140 7564 39142
rect 7620 39140 7644 39142
rect 7700 39140 7724 39142
rect 7780 39140 7786 39142
rect 7478 39120 7786 39140
rect 9680 38956 9732 38962
rect 9680 38898 9732 38904
rect 9110 38652 9418 38672
rect 9110 38650 9116 38652
rect 9172 38650 9196 38652
rect 9252 38650 9276 38652
rect 9332 38650 9356 38652
rect 9412 38650 9418 38652
rect 9172 38598 9174 38650
rect 9354 38598 9356 38650
rect 9110 38596 9116 38598
rect 9172 38596 9196 38598
rect 9252 38596 9276 38598
rect 9332 38596 9356 38598
rect 9412 38596 9418 38598
rect 9110 38576 9418 38596
rect 7478 38108 7786 38128
rect 7478 38106 7484 38108
rect 7540 38106 7564 38108
rect 7620 38106 7644 38108
rect 7700 38106 7724 38108
rect 7780 38106 7786 38108
rect 7540 38054 7542 38106
rect 7722 38054 7724 38106
rect 7478 38052 7484 38054
rect 7540 38052 7564 38054
rect 7620 38052 7644 38054
rect 7700 38052 7724 38054
rect 7780 38052 7786 38054
rect 7478 38032 7786 38052
rect 9110 37564 9418 37584
rect 9110 37562 9116 37564
rect 9172 37562 9196 37564
rect 9252 37562 9276 37564
rect 9332 37562 9356 37564
rect 9412 37562 9418 37564
rect 9172 37510 9174 37562
rect 9354 37510 9356 37562
rect 9110 37508 9116 37510
rect 9172 37508 9196 37510
rect 9252 37508 9276 37510
rect 9332 37508 9356 37510
rect 9412 37508 9418 37510
rect 9110 37488 9418 37508
rect 7478 37020 7786 37040
rect 7478 37018 7484 37020
rect 7540 37018 7564 37020
rect 7620 37018 7644 37020
rect 7700 37018 7724 37020
rect 7780 37018 7786 37020
rect 7540 36966 7542 37018
rect 7722 36966 7724 37018
rect 7478 36964 7484 36966
rect 7540 36964 7564 36966
rect 7620 36964 7644 36966
rect 7700 36964 7724 36966
rect 7780 36964 7786 36966
rect 7478 36944 7786 36964
rect 9110 36476 9418 36496
rect 9110 36474 9116 36476
rect 9172 36474 9196 36476
rect 9252 36474 9276 36476
rect 9332 36474 9356 36476
rect 9412 36474 9418 36476
rect 9172 36422 9174 36474
rect 9354 36422 9356 36474
rect 9110 36420 9116 36422
rect 9172 36420 9196 36422
rect 9252 36420 9276 36422
rect 9332 36420 9356 36422
rect 9412 36420 9418 36422
rect 9110 36400 9418 36420
rect 9692 36378 9720 38898
rect 9876 38010 9904 39986
rect 10048 39840 10100 39846
rect 10048 39782 10100 39788
rect 10060 39545 10088 39782
rect 10046 39536 10102 39545
rect 10046 39471 10102 39480
rect 10048 38752 10100 38758
rect 10046 38720 10048 38729
rect 10100 38720 10102 38729
rect 10046 38655 10102 38664
rect 9956 38344 10008 38350
rect 9956 38286 10008 38292
rect 9864 38004 9916 38010
rect 9864 37946 9916 37952
rect 9864 37256 9916 37262
rect 9864 37198 9916 37204
rect 9680 36372 9732 36378
rect 9680 36314 9732 36320
rect 9772 36168 9824 36174
rect 9772 36110 9824 36116
rect 7478 35932 7786 35952
rect 7478 35930 7484 35932
rect 7540 35930 7564 35932
rect 7620 35930 7644 35932
rect 7700 35930 7724 35932
rect 7780 35930 7786 35932
rect 7540 35878 7542 35930
rect 7722 35878 7724 35930
rect 7478 35876 7484 35878
rect 7540 35876 7564 35878
rect 7620 35876 7644 35878
rect 7700 35876 7724 35878
rect 7780 35876 7786 35878
rect 7478 35856 7786 35876
rect 9110 35388 9418 35408
rect 9110 35386 9116 35388
rect 9172 35386 9196 35388
rect 9252 35386 9276 35388
rect 9332 35386 9356 35388
rect 9412 35386 9418 35388
rect 9172 35334 9174 35386
rect 9354 35334 9356 35386
rect 9110 35332 9116 35334
rect 9172 35332 9196 35334
rect 9252 35332 9276 35334
rect 9332 35332 9356 35334
rect 9412 35332 9418 35334
rect 9110 35312 9418 35332
rect 7478 34844 7786 34864
rect 7478 34842 7484 34844
rect 7540 34842 7564 34844
rect 7620 34842 7644 34844
rect 7700 34842 7724 34844
rect 7780 34842 7786 34844
rect 7540 34790 7542 34842
rect 7722 34790 7724 34842
rect 7478 34788 7484 34790
rect 7540 34788 7564 34790
rect 7620 34788 7644 34790
rect 7700 34788 7724 34790
rect 7780 34788 7786 34790
rect 7478 34768 7786 34788
rect 9588 34740 9640 34746
rect 9588 34682 9640 34688
rect 9110 34300 9418 34320
rect 9110 34298 9116 34300
rect 9172 34298 9196 34300
rect 9252 34298 9276 34300
rect 9332 34298 9356 34300
rect 9412 34298 9418 34300
rect 9172 34246 9174 34298
rect 9354 34246 9356 34298
rect 9110 34244 9116 34246
rect 9172 34244 9196 34246
rect 9252 34244 9276 34246
rect 9332 34244 9356 34246
rect 9412 34244 9418 34246
rect 9110 34224 9418 34244
rect 9600 34105 9628 34682
rect 9680 34604 9732 34610
rect 9680 34546 9732 34552
rect 9586 34096 9642 34105
rect 9586 34031 9642 34040
rect 7478 33756 7786 33776
rect 7478 33754 7484 33756
rect 7540 33754 7564 33756
rect 7620 33754 7644 33756
rect 7700 33754 7724 33756
rect 7780 33754 7786 33756
rect 7540 33702 7542 33754
rect 7722 33702 7724 33754
rect 7478 33700 7484 33702
rect 7540 33700 7564 33702
rect 7620 33700 7644 33702
rect 7700 33700 7724 33702
rect 7780 33700 7786 33702
rect 7478 33680 7786 33700
rect 9110 33212 9418 33232
rect 9110 33210 9116 33212
rect 9172 33210 9196 33212
rect 9252 33210 9276 33212
rect 9332 33210 9356 33212
rect 9412 33210 9418 33212
rect 9172 33158 9174 33210
rect 9354 33158 9356 33210
rect 9110 33156 9116 33158
rect 9172 33156 9196 33158
rect 9252 33156 9276 33158
rect 9332 33156 9356 33158
rect 9412 33156 9418 33158
rect 9110 33136 9418 33156
rect 9692 33114 9720 34546
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 7478 32668 7786 32688
rect 7478 32666 7484 32668
rect 7540 32666 7564 32668
rect 7620 32666 7644 32668
rect 7700 32666 7724 32668
rect 7780 32666 7786 32668
rect 7540 32614 7542 32666
rect 7722 32614 7724 32666
rect 7478 32612 7484 32614
rect 7540 32612 7564 32614
rect 7620 32612 7644 32614
rect 7700 32612 7724 32614
rect 7780 32612 7786 32614
rect 7478 32592 7786 32612
rect 9110 32124 9418 32144
rect 9110 32122 9116 32124
rect 9172 32122 9196 32124
rect 9252 32122 9276 32124
rect 9332 32122 9356 32124
rect 9412 32122 9418 32124
rect 9172 32070 9174 32122
rect 9354 32070 9356 32122
rect 9110 32068 9116 32070
rect 9172 32068 9196 32070
rect 9252 32068 9276 32070
rect 9332 32068 9356 32070
rect 9412 32068 9418 32070
rect 9110 32048 9418 32068
rect 9784 32026 9812 36110
rect 9876 34202 9904 37198
rect 9968 35834 9996 38286
rect 10048 38208 10100 38214
rect 10048 38150 10100 38156
rect 10060 38049 10088 38150
rect 10046 38040 10102 38049
rect 10046 37975 10102 37984
rect 10232 37868 10284 37874
rect 10232 37810 10284 37816
rect 10046 37224 10102 37233
rect 10046 37159 10102 37168
rect 10060 37126 10088 37159
rect 10048 37120 10100 37126
rect 10048 37062 10100 37068
rect 10140 36780 10192 36786
rect 10140 36722 10192 36728
rect 10048 36576 10100 36582
rect 10048 36518 10100 36524
rect 10060 36417 10088 36518
rect 10046 36408 10102 36417
rect 10046 36343 10102 36352
rect 10048 36032 10100 36038
rect 10048 35974 10100 35980
rect 9956 35828 10008 35834
rect 9956 35770 10008 35776
rect 10060 35737 10088 35974
rect 10046 35728 10102 35737
rect 10046 35663 10102 35672
rect 10048 34944 10100 34950
rect 10046 34912 10048 34921
rect 10100 34912 10102 34921
rect 10046 34847 10102 34856
rect 9864 34196 9916 34202
rect 9864 34138 9916 34144
rect 10152 34134 10180 36722
rect 10244 34678 10272 37810
rect 10232 34672 10284 34678
rect 10232 34614 10284 34620
rect 10140 34128 10192 34134
rect 10140 34070 10192 34076
rect 10140 33992 10192 33998
rect 10140 33934 10192 33940
rect 10152 33658 10180 33934
rect 10140 33652 10192 33658
rect 10140 33594 10192 33600
rect 10046 33416 10102 33425
rect 10046 33351 10048 33360
rect 10100 33351 10102 33360
rect 10048 33322 10100 33328
rect 9864 32904 9916 32910
rect 9864 32846 9916 32852
rect 9876 32570 9904 32846
rect 10048 32768 10100 32774
rect 10048 32710 10100 32716
rect 10060 32609 10088 32710
rect 10046 32600 10102 32609
rect 9864 32564 9916 32570
rect 10046 32535 10102 32544
rect 9864 32506 9916 32512
rect 9772 32020 9824 32026
rect 9772 31962 9824 31968
rect 10048 31952 10100 31958
rect 10048 31894 10100 31900
rect 10060 31793 10088 31894
rect 10046 31784 10102 31793
rect 10046 31719 10102 31728
rect 7478 31580 7786 31600
rect 7478 31578 7484 31580
rect 7540 31578 7564 31580
rect 7620 31578 7644 31580
rect 7700 31578 7724 31580
rect 7780 31578 7786 31580
rect 7540 31526 7542 31578
rect 7722 31526 7724 31578
rect 7478 31524 7484 31526
rect 7540 31524 7564 31526
rect 7620 31524 7644 31526
rect 7700 31524 7724 31526
rect 7780 31524 7786 31526
rect 7478 31504 7786 31524
rect 9864 31340 9916 31346
rect 9864 31282 9916 31288
rect 9110 31036 9418 31056
rect 9110 31034 9116 31036
rect 9172 31034 9196 31036
rect 9252 31034 9276 31036
rect 9332 31034 9356 31036
rect 9412 31034 9418 31036
rect 9172 30982 9174 31034
rect 9354 30982 9356 31034
rect 9110 30980 9116 30982
rect 9172 30980 9196 30982
rect 9252 30980 9276 30982
rect 9332 30980 9356 30982
rect 9412 30980 9418 30982
rect 9110 30960 9418 30980
rect 8300 30728 8352 30734
rect 8300 30670 8352 30676
rect 7478 30492 7786 30512
rect 7478 30490 7484 30492
rect 7540 30490 7564 30492
rect 7620 30490 7644 30492
rect 7700 30490 7724 30492
rect 7780 30490 7786 30492
rect 7540 30438 7542 30490
rect 7722 30438 7724 30490
rect 7478 30436 7484 30438
rect 7540 30436 7564 30438
rect 7620 30436 7644 30438
rect 7700 30436 7724 30438
rect 7780 30436 7786 30438
rect 7478 30416 7786 30436
rect 8312 29850 8340 30670
rect 9876 30054 9904 31282
rect 10048 31136 10100 31142
rect 10046 31104 10048 31113
rect 10100 31104 10102 31113
rect 10046 31039 10102 31048
rect 10048 30592 10100 30598
rect 10048 30534 10100 30540
rect 10060 30297 10088 30534
rect 10046 30288 10102 30297
rect 10046 30223 10102 30232
rect 9864 30048 9916 30054
rect 9864 29990 9916 29996
rect 9110 29948 9418 29968
rect 9110 29946 9116 29948
rect 9172 29946 9196 29948
rect 9252 29946 9276 29948
rect 9332 29946 9356 29948
rect 9412 29946 9418 29948
rect 9172 29894 9174 29946
rect 9354 29894 9356 29946
rect 9110 29892 9116 29894
rect 9172 29892 9196 29894
rect 9252 29892 9276 29894
rect 9332 29892 9356 29894
rect 9412 29892 9418 29894
rect 9110 29872 9418 29892
rect 8300 29844 8352 29850
rect 8300 29786 8352 29792
rect 7840 29640 7892 29646
rect 7840 29582 7892 29588
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 7478 29404 7786 29424
rect 7478 29402 7484 29404
rect 7540 29402 7564 29404
rect 7620 29402 7644 29404
rect 7700 29402 7724 29404
rect 7780 29402 7786 29404
rect 7540 29350 7542 29402
rect 7722 29350 7724 29402
rect 7478 29348 7484 29350
rect 7540 29348 7564 29350
rect 7620 29348 7644 29350
rect 7700 29348 7724 29350
rect 7780 29348 7786 29350
rect 7478 29328 7786 29348
rect 7478 28316 7786 28336
rect 7478 28314 7484 28316
rect 7540 28314 7564 28316
rect 7620 28314 7644 28316
rect 7700 28314 7724 28316
rect 7780 28314 7786 28316
rect 7540 28262 7542 28314
rect 7722 28262 7724 28314
rect 7478 28260 7484 28262
rect 7540 28260 7564 28262
rect 7620 28260 7644 28262
rect 7700 28260 7724 28262
rect 7780 28260 7786 28262
rect 7478 28240 7786 28260
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 7478 27228 7786 27248
rect 7478 27226 7484 27228
rect 7540 27226 7564 27228
rect 7620 27226 7644 27228
rect 7700 27226 7724 27228
rect 7780 27226 7786 27228
rect 7540 27174 7542 27226
rect 7722 27174 7724 27226
rect 7478 27172 7484 27174
rect 7540 27172 7564 27174
rect 7620 27172 7644 27174
rect 7700 27172 7724 27174
rect 7780 27172 7786 27174
rect 7478 27152 7786 27172
rect 6276 26444 6328 26450
rect 6276 26386 6328 26392
rect 7478 26140 7786 26160
rect 7478 26138 7484 26140
rect 7540 26138 7564 26140
rect 7620 26138 7644 26140
rect 7700 26138 7724 26140
rect 7780 26138 7786 26140
rect 7540 26086 7542 26138
rect 7722 26086 7724 26138
rect 7478 26084 7484 26086
rect 7540 26084 7564 26086
rect 7620 26084 7644 26086
rect 7700 26084 7724 26086
rect 7780 26084 7786 26086
rect 7478 26064 7786 26084
rect 5846 25596 6154 25616
rect 5846 25594 5852 25596
rect 5908 25594 5932 25596
rect 5988 25594 6012 25596
rect 6068 25594 6092 25596
rect 6148 25594 6154 25596
rect 5908 25542 5910 25594
rect 6090 25542 6092 25594
rect 5846 25540 5852 25542
rect 5908 25540 5932 25542
rect 5988 25540 6012 25542
rect 6068 25540 6092 25542
rect 6148 25540 6154 25542
rect 5846 25520 6154 25540
rect 7478 25052 7786 25072
rect 7478 25050 7484 25052
rect 7540 25050 7564 25052
rect 7620 25050 7644 25052
rect 7700 25050 7724 25052
rect 7780 25050 7786 25052
rect 7540 24998 7542 25050
rect 7722 24998 7724 25050
rect 7478 24996 7484 24998
rect 7540 24996 7564 24998
rect 7620 24996 7644 24998
rect 7700 24996 7724 24998
rect 7780 24996 7786 24998
rect 7478 24976 7786 24996
rect 5846 24508 6154 24528
rect 5846 24506 5852 24508
rect 5908 24506 5932 24508
rect 5988 24506 6012 24508
rect 6068 24506 6092 24508
rect 6148 24506 6154 24508
rect 5908 24454 5910 24506
rect 6090 24454 6092 24506
rect 5846 24452 5852 24454
rect 5908 24452 5932 24454
rect 5988 24452 6012 24454
rect 6068 24452 6092 24454
rect 6148 24452 6154 24454
rect 5846 24432 6154 24452
rect 7478 23964 7786 23984
rect 7478 23962 7484 23964
rect 7540 23962 7564 23964
rect 7620 23962 7644 23964
rect 7700 23962 7724 23964
rect 7780 23962 7786 23964
rect 7540 23910 7542 23962
rect 7722 23910 7724 23962
rect 7478 23908 7484 23910
rect 7540 23908 7564 23910
rect 7620 23908 7644 23910
rect 7700 23908 7724 23910
rect 7780 23908 7786 23910
rect 7478 23888 7786 23908
rect 5846 23420 6154 23440
rect 5846 23418 5852 23420
rect 5908 23418 5932 23420
rect 5988 23418 6012 23420
rect 6068 23418 6092 23420
rect 6148 23418 6154 23420
rect 5908 23366 5910 23418
rect 6090 23366 6092 23418
rect 5846 23364 5852 23366
rect 5908 23364 5932 23366
rect 5988 23364 6012 23366
rect 6068 23364 6092 23366
rect 6148 23364 6154 23366
rect 5846 23344 6154 23364
rect 7478 22876 7786 22896
rect 7478 22874 7484 22876
rect 7540 22874 7564 22876
rect 7620 22874 7644 22876
rect 7700 22874 7724 22876
rect 7780 22874 7786 22876
rect 7540 22822 7542 22874
rect 7722 22822 7724 22874
rect 7478 22820 7484 22822
rect 7540 22820 7564 22822
rect 7620 22820 7644 22822
rect 7700 22820 7724 22822
rect 7780 22820 7786 22822
rect 7478 22800 7786 22820
rect 5846 22332 6154 22352
rect 5846 22330 5852 22332
rect 5908 22330 5932 22332
rect 5988 22330 6012 22332
rect 6068 22330 6092 22332
rect 6148 22330 6154 22332
rect 5908 22278 5910 22330
rect 6090 22278 6092 22330
rect 5846 22276 5852 22278
rect 5908 22276 5932 22278
rect 5988 22276 6012 22278
rect 6068 22276 6092 22278
rect 6148 22276 6154 22278
rect 5846 22256 6154 22276
rect 7478 21788 7786 21808
rect 7478 21786 7484 21788
rect 7540 21786 7564 21788
rect 7620 21786 7644 21788
rect 7700 21786 7724 21788
rect 7780 21786 7786 21788
rect 7540 21734 7542 21786
rect 7722 21734 7724 21786
rect 7478 21732 7484 21734
rect 7540 21732 7564 21734
rect 7620 21732 7644 21734
rect 7700 21732 7724 21734
rect 7780 21732 7786 21734
rect 7478 21712 7786 21732
rect 5846 21244 6154 21264
rect 5846 21242 5852 21244
rect 5908 21242 5932 21244
rect 5988 21242 6012 21244
rect 6068 21242 6092 21244
rect 6148 21242 6154 21244
rect 5908 21190 5910 21242
rect 6090 21190 6092 21242
rect 5846 21188 5852 21190
rect 5908 21188 5932 21190
rect 5988 21188 6012 21190
rect 6068 21188 6092 21190
rect 6148 21188 6154 21190
rect 5846 21168 6154 21188
rect 7478 20700 7786 20720
rect 7478 20698 7484 20700
rect 7540 20698 7564 20700
rect 7620 20698 7644 20700
rect 7700 20698 7724 20700
rect 7780 20698 7786 20700
rect 7540 20646 7542 20698
rect 7722 20646 7724 20698
rect 7478 20644 7484 20646
rect 7540 20644 7564 20646
rect 7620 20644 7644 20646
rect 7700 20644 7724 20646
rect 7780 20644 7786 20646
rect 7478 20624 7786 20644
rect 7852 20602 7880 29582
rect 10152 29481 10180 29582
rect 10138 29472 10194 29481
rect 10138 29407 10194 29416
rect 10140 29028 10192 29034
rect 10140 28970 10192 28976
rect 9110 28860 9418 28880
rect 9110 28858 9116 28860
rect 9172 28858 9196 28860
rect 9252 28858 9276 28860
rect 9332 28858 9356 28860
rect 9412 28858 9418 28860
rect 9172 28806 9174 28858
rect 9354 28806 9356 28858
rect 9110 28804 9116 28806
rect 9172 28804 9196 28806
rect 9252 28804 9276 28806
rect 9332 28804 9356 28806
rect 9412 28804 9418 28806
rect 9110 28784 9418 28804
rect 10152 28801 10180 28970
rect 10138 28792 10194 28801
rect 10138 28727 10194 28736
rect 9956 28008 10008 28014
rect 9954 27976 9956 27985
rect 10008 27976 10010 27985
rect 9954 27911 10010 27920
rect 9110 27772 9418 27792
rect 9110 27770 9116 27772
rect 9172 27770 9196 27772
rect 9252 27770 9276 27772
rect 9332 27770 9356 27772
rect 9412 27770 9418 27772
rect 9172 27718 9174 27770
rect 9354 27718 9356 27770
rect 9110 27716 9116 27718
rect 9172 27716 9196 27718
rect 9252 27716 9276 27718
rect 9332 27716 9356 27718
rect 9412 27716 9418 27718
rect 9110 27696 9418 27716
rect 9956 27328 10008 27334
rect 9956 27270 10008 27276
rect 9968 27169 9996 27270
rect 9954 27160 10010 27169
rect 9954 27095 10010 27104
rect 10140 26784 10192 26790
rect 10140 26726 10192 26732
rect 9110 26684 9418 26704
rect 9110 26682 9116 26684
rect 9172 26682 9196 26684
rect 9252 26682 9276 26684
rect 9332 26682 9356 26684
rect 9412 26682 9418 26684
rect 9172 26630 9174 26682
rect 9354 26630 9356 26682
rect 9110 26628 9116 26630
rect 9172 26628 9196 26630
rect 9252 26628 9276 26630
rect 9332 26628 9356 26630
rect 9412 26628 9418 26630
rect 9110 26608 9418 26628
rect 10152 26489 10180 26726
rect 10138 26480 10194 26489
rect 10138 26415 10194 26424
rect 10140 25696 10192 25702
rect 10138 25664 10140 25673
rect 10192 25664 10194 25673
rect 9110 25596 9418 25616
rect 10138 25599 10194 25608
rect 9110 25594 9116 25596
rect 9172 25594 9196 25596
rect 9252 25594 9276 25596
rect 9332 25594 9356 25596
rect 9412 25594 9418 25596
rect 9172 25542 9174 25594
rect 9354 25542 9356 25594
rect 9110 25540 9116 25542
rect 9172 25540 9196 25542
rect 9252 25540 9276 25542
rect 9332 25540 9356 25542
rect 9412 25540 9418 25542
rect 9110 25520 9418 25540
rect 10140 25288 10192 25294
rect 10140 25230 10192 25236
rect 10152 24857 10180 25230
rect 10138 24848 10194 24857
rect 10138 24783 10194 24792
rect 9110 24508 9418 24528
rect 9110 24506 9116 24508
rect 9172 24506 9196 24508
rect 9252 24506 9276 24508
rect 9332 24506 9356 24508
rect 9412 24506 9418 24508
rect 9172 24454 9174 24506
rect 9354 24454 9356 24506
rect 9110 24452 9116 24454
rect 9172 24452 9196 24454
rect 9252 24452 9276 24454
rect 9332 24452 9356 24454
rect 9412 24452 9418 24454
rect 9110 24432 9418 24452
rect 10140 24200 10192 24206
rect 10138 24168 10140 24177
rect 10192 24168 10194 24177
rect 10138 24103 10194 24112
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 9110 23420 9418 23440
rect 9110 23418 9116 23420
rect 9172 23418 9196 23420
rect 9252 23418 9276 23420
rect 9332 23418 9356 23420
rect 9412 23418 9418 23420
rect 9172 23366 9174 23418
rect 9354 23366 9356 23418
rect 9110 23364 9116 23366
rect 9172 23364 9196 23366
rect 9252 23364 9276 23366
rect 9332 23364 9356 23366
rect 9412 23364 9418 23366
rect 9110 23344 9418 23364
rect 10152 23361 10180 23462
rect 10138 23352 10194 23361
rect 10138 23287 10194 23296
rect 10138 22536 10194 22545
rect 10138 22471 10140 22480
rect 10192 22471 10194 22480
rect 10140 22442 10192 22448
rect 9110 22332 9418 22352
rect 9110 22330 9116 22332
rect 9172 22330 9196 22332
rect 9252 22330 9276 22332
rect 9332 22330 9356 22332
rect 9412 22330 9418 22332
rect 9172 22278 9174 22330
rect 9354 22278 9356 22330
rect 9110 22276 9116 22278
rect 9172 22276 9196 22278
rect 9252 22276 9276 22278
rect 9332 22276 9356 22278
rect 9412 22276 9418 22278
rect 9110 22256 9418 22276
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 10152 21865 10180 22102
rect 10138 21856 10194 21865
rect 10138 21791 10194 21800
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 9110 21244 9418 21264
rect 9110 21242 9116 21244
rect 9172 21242 9196 21244
rect 9252 21242 9276 21244
rect 9332 21242 9356 21244
rect 9412 21242 9418 21244
rect 9172 21190 9174 21242
rect 9354 21190 9356 21242
rect 9110 21188 9116 21190
rect 9172 21188 9196 21190
rect 9252 21188 9276 21190
rect 9332 21188 9356 21190
rect 9412 21188 9418 21190
rect 9110 21168 9418 21188
rect 10152 21049 10180 21286
rect 10138 21040 10194 21049
rect 10138 20975 10194 20984
rect 7840 20596 7892 20602
rect 7840 20538 7892 20544
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 5846 20156 6154 20176
rect 5846 20154 5852 20156
rect 5908 20154 5932 20156
rect 5988 20154 6012 20156
rect 6068 20154 6092 20156
rect 6148 20154 6154 20156
rect 5908 20102 5910 20154
rect 6090 20102 6092 20154
rect 5846 20100 5852 20102
rect 5908 20100 5932 20102
rect 5988 20100 6012 20102
rect 6068 20100 6092 20102
rect 6148 20100 6154 20102
rect 5846 20080 6154 20100
rect 9110 20156 9418 20176
rect 9110 20154 9116 20156
rect 9172 20154 9196 20156
rect 9252 20154 9276 20156
rect 9332 20154 9356 20156
rect 9412 20154 9418 20156
rect 9172 20102 9174 20154
rect 9354 20102 9356 20154
rect 9110 20100 9116 20102
rect 9172 20100 9196 20102
rect 9252 20100 9276 20102
rect 9332 20100 9356 20102
rect 9412 20100 9418 20102
rect 9110 20080 9418 20100
rect 7478 19612 7786 19632
rect 7478 19610 7484 19612
rect 7540 19610 7564 19612
rect 7620 19610 7644 19612
rect 7700 19610 7724 19612
rect 7780 19610 7786 19612
rect 7540 19558 7542 19610
rect 7722 19558 7724 19610
rect 7478 19556 7484 19558
rect 7540 19556 7564 19558
rect 7620 19556 7644 19558
rect 7700 19556 7724 19558
rect 7780 19556 7786 19558
rect 7478 19536 7786 19556
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5846 19068 6154 19088
rect 5846 19066 5852 19068
rect 5908 19066 5932 19068
rect 5988 19066 6012 19068
rect 6068 19066 6092 19068
rect 6148 19066 6154 19068
rect 5908 19014 5910 19066
rect 6090 19014 6092 19066
rect 5846 19012 5852 19014
rect 5908 19012 5932 19014
rect 5988 19012 6012 19014
rect 6068 19012 6092 19014
rect 6148 19012 6154 19014
rect 5846 18992 6154 19012
rect 9110 19068 9418 19088
rect 9110 19066 9116 19068
rect 9172 19066 9196 19068
rect 9252 19066 9276 19068
rect 9332 19066 9356 19068
rect 9412 19066 9418 19068
rect 9172 19014 9174 19066
rect 9354 19014 9356 19066
rect 9110 19012 9116 19014
rect 9172 19012 9196 19014
rect 9252 19012 9276 19014
rect 9332 19012 9356 19014
rect 9412 19012 9418 19014
rect 9110 18992 9418 19012
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 7478 18524 7786 18544
rect 7478 18522 7484 18524
rect 7540 18522 7564 18524
rect 7620 18522 7644 18524
rect 7700 18522 7724 18524
rect 7780 18522 7786 18524
rect 7540 18470 7542 18522
rect 7722 18470 7724 18522
rect 7478 18468 7484 18470
rect 7540 18468 7564 18470
rect 7620 18468 7644 18470
rect 7700 18468 7724 18470
rect 7780 18468 7786 18470
rect 7478 18448 7786 18468
rect 9232 18426 9260 18702
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5460 17202 5488 18294
rect 5846 17980 6154 18000
rect 5846 17978 5852 17980
rect 5908 17978 5932 17980
rect 5988 17978 6012 17980
rect 6068 17978 6092 17980
rect 6148 17978 6154 17980
rect 5908 17926 5910 17978
rect 6090 17926 6092 17978
rect 5846 17924 5852 17926
rect 5908 17924 5932 17926
rect 5988 17924 6012 17926
rect 6068 17924 6092 17926
rect 6148 17924 6154 17926
rect 5846 17904 6154 17924
rect 9110 17980 9418 18000
rect 9110 17978 9116 17980
rect 9172 17978 9196 17980
rect 9252 17978 9276 17980
rect 9332 17978 9356 17980
rect 9412 17978 9418 17980
rect 9172 17926 9174 17978
rect 9354 17926 9356 17978
rect 9110 17924 9116 17926
rect 9172 17924 9196 17926
rect 9252 17924 9276 17926
rect 9332 17924 9356 17926
rect 9412 17924 9418 17926
rect 9110 17904 9418 17924
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 7478 17436 7786 17456
rect 7478 17434 7484 17436
rect 7540 17434 7564 17436
rect 7620 17434 7644 17436
rect 7700 17434 7724 17436
rect 7780 17434 7786 17436
rect 7540 17382 7542 17434
rect 7722 17382 7724 17434
rect 7478 17380 7484 17382
rect 7540 17380 7564 17382
rect 7620 17380 7644 17382
rect 7700 17380 7724 17382
rect 7780 17380 7786 17382
rect 7478 17360 7786 17380
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5846 16892 6154 16912
rect 5846 16890 5852 16892
rect 5908 16890 5932 16892
rect 5988 16890 6012 16892
rect 6068 16890 6092 16892
rect 6148 16890 6154 16892
rect 5908 16838 5910 16890
rect 6090 16838 6092 16890
rect 5846 16836 5852 16838
rect 5908 16836 5932 16838
rect 5988 16836 6012 16838
rect 6068 16836 6092 16838
rect 6148 16836 6154 16838
rect 5846 16816 6154 16836
rect 9110 16892 9418 16912
rect 9110 16890 9116 16892
rect 9172 16890 9196 16892
rect 9252 16890 9276 16892
rect 9332 16890 9356 16892
rect 9412 16890 9418 16892
rect 9172 16838 9174 16890
rect 9354 16838 9356 16890
rect 9110 16836 9116 16838
rect 9172 16836 9196 16838
rect 9252 16836 9276 16838
rect 9332 16836 9356 16838
rect 9412 16836 9418 16838
rect 9110 16816 9418 16836
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 7478 16348 7786 16368
rect 7478 16346 7484 16348
rect 7540 16346 7564 16348
rect 7620 16346 7644 16348
rect 7700 16346 7724 16348
rect 7780 16346 7786 16348
rect 7540 16294 7542 16346
rect 7722 16294 7724 16346
rect 7478 16292 7484 16294
rect 7540 16292 7564 16294
rect 7620 16292 7644 16294
rect 7700 16292 7724 16294
rect 7780 16292 7786 16294
rect 7478 16272 7786 16292
rect 9508 16250 9536 17614
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 5846 15804 6154 15824
rect 5846 15802 5852 15804
rect 5908 15802 5932 15804
rect 5988 15802 6012 15804
rect 6068 15802 6092 15804
rect 6148 15802 6154 15804
rect 5908 15750 5910 15802
rect 6090 15750 6092 15802
rect 5846 15748 5852 15750
rect 5908 15748 5932 15750
rect 5988 15748 6012 15750
rect 6068 15748 6092 15750
rect 6148 15748 6154 15750
rect 5846 15728 6154 15748
rect 6196 15570 6224 16050
rect 9110 15804 9418 15824
rect 9110 15802 9116 15804
rect 9172 15802 9196 15804
rect 9252 15802 9276 15804
rect 9332 15802 9356 15804
rect 9412 15802 9418 15804
rect 9172 15750 9174 15802
rect 9354 15750 9356 15802
rect 9110 15748 9116 15750
rect 9172 15748 9196 15750
rect 9252 15748 9276 15750
rect 9332 15748 9356 15750
rect 9412 15748 9418 15750
rect 9110 15728 9418 15748
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 7478 15260 7786 15280
rect 7478 15258 7484 15260
rect 7540 15258 7564 15260
rect 7620 15258 7644 15260
rect 7700 15258 7724 15260
rect 7780 15258 7786 15260
rect 7540 15206 7542 15258
rect 7722 15206 7724 15258
rect 7478 15204 7484 15206
rect 7540 15204 7564 15206
rect 7620 15204 7644 15206
rect 7700 15204 7724 15206
rect 7780 15204 7786 15206
rect 7478 15184 7786 15204
rect 5846 14716 6154 14736
rect 5846 14714 5852 14716
rect 5908 14714 5932 14716
rect 5988 14714 6012 14716
rect 6068 14714 6092 14716
rect 6148 14714 6154 14716
rect 5908 14662 5910 14714
rect 6090 14662 6092 14714
rect 5846 14660 5852 14662
rect 5908 14660 5932 14662
rect 5988 14660 6012 14662
rect 6068 14660 6092 14662
rect 6148 14660 6154 14662
rect 5846 14640 6154 14660
rect 9110 14716 9418 14736
rect 9110 14714 9116 14716
rect 9172 14714 9196 14716
rect 9252 14714 9276 14716
rect 9332 14714 9356 14716
rect 9412 14714 9418 14716
rect 9172 14662 9174 14714
rect 9354 14662 9356 14714
rect 9110 14660 9116 14662
rect 9172 14660 9196 14662
rect 9252 14660 9276 14662
rect 9332 14660 9356 14662
rect 9412 14660 9418 14662
rect 9110 14640 9418 14660
rect 7478 14172 7786 14192
rect 7478 14170 7484 14172
rect 7540 14170 7564 14172
rect 7620 14170 7644 14172
rect 7700 14170 7724 14172
rect 7780 14170 7786 14172
rect 7540 14118 7542 14170
rect 7722 14118 7724 14170
rect 7478 14116 7484 14118
rect 7540 14116 7564 14118
rect 7620 14116 7644 14118
rect 7700 14116 7724 14118
rect 7780 14116 7786 14118
rect 7478 14096 7786 14116
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 5846 13628 6154 13648
rect 5846 13626 5852 13628
rect 5908 13626 5932 13628
rect 5988 13626 6012 13628
rect 6068 13626 6092 13628
rect 6148 13626 6154 13628
rect 5908 13574 5910 13626
rect 6090 13574 6092 13626
rect 5846 13572 5852 13574
rect 5908 13572 5932 13574
rect 5988 13572 6012 13574
rect 6068 13572 6092 13574
rect 6148 13572 6154 13574
rect 5846 13552 6154 13572
rect 9110 13628 9418 13648
rect 9110 13626 9116 13628
rect 9172 13626 9196 13628
rect 9252 13626 9276 13628
rect 9332 13626 9356 13628
rect 9412 13626 9418 13628
rect 9172 13574 9174 13626
rect 9354 13574 9356 13626
rect 9110 13572 9116 13574
rect 9172 13572 9196 13574
rect 9252 13572 9276 13574
rect 9332 13572 9356 13574
rect 9412 13572 9418 13574
rect 9110 13552 9418 13572
rect 9600 13433 9628 14010
rect 9586 13424 9642 13433
rect 9586 13359 9642 13368
rect 9692 13190 9720 16050
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 7478 13084 7786 13104
rect 7478 13082 7484 13084
rect 7540 13082 7564 13084
rect 7620 13082 7644 13084
rect 7700 13082 7724 13084
rect 7780 13082 7786 13084
rect 7540 13030 7542 13082
rect 7722 13030 7724 13082
rect 7478 13028 7484 13030
rect 7540 13028 7564 13030
rect 7620 13028 7644 13030
rect 7700 13028 7724 13030
rect 7780 13028 7786 13030
rect 7478 13008 7786 13028
rect 9784 12986 9812 20402
rect 10046 20360 10102 20369
rect 10046 20295 10048 20304
rect 10100 20295 10102 20304
rect 10048 20266 10100 20272
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9876 19514 9904 19790
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10060 19553 10088 19654
rect 10046 19544 10102 19553
rect 9864 19508 9916 19514
rect 10046 19479 10102 19488
rect 9864 19450 9916 19456
rect 10046 18728 10102 18737
rect 10046 18663 10102 18672
rect 10060 18630 10088 18663
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9876 17338 9904 18226
rect 10048 18080 10100 18086
rect 10046 18048 10048 18057
rect 10100 18048 10102 18057
rect 10046 17983 10102 17992
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 10060 17241 10088 17478
rect 10046 17232 10102 17241
rect 10046 17167 10102 17176
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9968 15706 9996 16526
rect 10048 16448 10100 16454
rect 10046 16416 10048 16425
rect 10100 16416 10102 16425
rect 10046 16351 10102 16360
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10060 15745 10088 15846
rect 10046 15736 10102 15745
rect 9956 15700 10008 15706
rect 10046 15671 10102 15680
rect 9956 15642 10008 15648
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9876 13530 9904 14350
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9876 12850 9904 13194
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 5846 12540 6154 12560
rect 5846 12538 5852 12540
rect 5908 12538 5932 12540
rect 5988 12538 6012 12540
rect 6068 12538 6092 12540
rect 6148 12538 6154 12540
rect 5908 12486 5910 12538
rect 6090 12486 6092 12538
rect 5846 12484 5852 12486
rect 5908 12484 5932 12486
rect 5988 12484 6012 12486
rect 6068 12484 6092 12486
rect 6148 12484 6154 12486
rect 5846 12464 6154 12484
rect 9110 12540 9418 12560
rect 9110 12538 9116 12540
rect 9172 12538 9196 12540
rect 9252 12538 9276 12540
rect 9332 12538 9356 12540
rect 9412 12538 9418 12540
rect 9172 12486 9174 12538
rect 9354 12486 9356 12538
rect 9110 12484 9116 12486
rect 9172 12484 9196 12486
rect 9252 12484 9276 12486
rect 9332 12484 9356 12486
rect 9412 12484 9418 12486
rect 9110 12464 9418 12484
rect 9968 12442 9996 14962
rect 10046 14920 10102 14929
rect 10046 14855 10048 14864
rect 10100 14855 10102 14864
rect 10048 14826 10100 14832
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 14113 10088 14214
rect 10046 14104 10102 14113
rect 10046 14039 10102 14048
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10152 12782 10180 13262
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10048 12640 10100 12646
rect 10046 12608 10048 12617
rect 10100 12608 10102 12617
rect 10046 12543 10102 12552
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 7478 11996 7786 12016
rect 7478 11994 7484 11996
rect 7540 11994 7564 11996
rect 7620 11994 7644 11996
rect 7700 11994 7724 11996
rect 7780 11994 7786 11996
rect 7540 11942 7542 11994
rect 7722 11942 7724 11994
rect 7478 11940 7484 11942
rect 7540 11940 7564 11942
rect 7620 11940 7644 11942
rect 7700 11940 7724 11942
rect 7780 11940 7786 11942
rect 7478 11920 7786 11940
rect 9876 11898 9904 12174
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 10060 11801 10088 12038
rect 10046 11792 10102 11801
rect 10046 11727 10102 11736
rect 5846 11452 6154 11472
rect 5846 11450 5852 11452
rect 5908 11450 5932 11452
rect 5988 11450 6012 11452
rect 6068 11450 6092 11452
rect 6148 11450 6154 11452
rect 5908 11398 5910 11450
rect 6090 11398 6092 11450
rect 5846 11396 5852 11398
rect 5908 11396 5932 11398
rect 5988 11396 6012 11398
rect 6068 11396 6092 11398
rect 6148 11396 6154 11398
rect 5846 11376 6154 11396
rect 9110 11452 9418 11472
rect 9110 11450 9116 11452
rect 9172 11450 9196 11452
rect 9252 11450 9276 11452
rect 9332 11450 9356 11452
rect 9412 11450 9418 11452
rect 9172 11398 9174 11450
rect 9354 11398 9356 11450
rect 9110 11396 9116 11398
rect 9172 11396 9196 11398
rect 9252 11396 9276 11398
rect 9332 11396 9356 11398
rect 9412 11396 9418 11398
rect 9110 11376 9418 11396
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10060 11121 10088 11222
rect 10046 11112 10102 11121
rect 10046 11047 10102 11056
rect 7478 10908 7786 10928
rect 7478 10906 7484 10908
rect 7540 10906 7564 10908
rect 7620 10906 7644 10908
rect 7700 10906 7724 10908
rect 7780 10906 7786 10908
rect 7540 10854 7542 10906
rect 7722 10854 7724 10906
rect 7478 10852 7484 10854
rect 7540 10852 7564 10854
rect 7620 10852 7644 10854
rect 7700 10852 7724 10854
rect 7780 10852 7786 10854
rect 7478 10832 7786 10852
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 5846 10364 6154 10384
rect 5846 10362 5852 10364
rect 5908 10362 5932 10364
rect 5988 10362 6012 10364
rect 6068 10362 6092 10364
rect 6148 10362 6154 10364
rect 5908 10310 5910 10362
rect 6090 10310 6092 10362
rect 5846 10308 5852 10310
rect 5908 10308 5932 10310
rect 5988 10308 6012 10310
rect 6068 10308 6092 10310
rect 6148 10308 6154 10310
rect 5846 10288 6154 10308
rect 9110 10364 9418 10384
rect 9110 10362 9116 10364
rect 9172 10362 9196 10364
rect 9252 10362 9276 10364
rect 9332 10362 9356 10364
rect 9412 10362 9418 10364
rect 9172 10310 9174 10362
rect 9354 10310 9356 10362
rect 9110 10308 9116 10310
rect 9172 10308 9196 10310
rect 9252 10308 9276 10310
rect 9332 10308 9356 10310
rect 9412 10308 9418 10310
rect 9110 10288 9418 10308
rect 10060 10305 10088 10406
rect 10046 10296 10102 10305
rect 10046 10231 10102 10240
rect 4214 9820 4522 9840
rect 4214 9818 4220 9820
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4516 9818 4522 9820
rect 4276 9766 4278 9818
rect 4458 9766 4460 9818
rect 4214 9764 4220 9766
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4516 9764 4522 9766
rect 4214 9744 4522 9764
rect 7478 9820 7786 9840
rect 7478 9818 7484 9820
rect 7540 9818 7564 9820
rect 7620 9818 7644 9820
rect 7700 9818 7724 9820
rect 7780 9818 7786 9820
rect 7540 9766 7542 9818
rect 7722 9766 7724 9818
rect 7478 9764 7484 9766
rect 7540 9764 7564 9766
rect 7620 9764 7644 9766
rect 7700 9764 7724 9766
rect 7780 9764 7786 9766
rect 7478 9744 7786 9764
rect 10046 9480 10102 9489
rect 10046 9415 10048 9424
rect 10100 9415 10102 9424
rect 10048 9386 10100 9392
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 5846 9276 6154 9296
rect 5846 9274 5852 9276
rect 5908 9274 5932 9276
rect 5988 9274 6012 9276
rect 6068 9274 6092 9276
rect 6148 9274 6154 9276
rect 5908 9222 5910 9274
rect 6090 9222 6092 9274
rect 5846 9220 5852 9222
rect 5908 9220 5932 9222
rect 5988 9220 6012 9222
rect 6068 9220 6092 9222
rect 6148 9220 6154 9222
rect 5846 9200 6154 9220
rect 9110 9276 9418 9296
rect 9110 9274 9116 9276
rect 9172 9274 9196 9276
rect 9252 9274 9276 9276
rect 9332 9274 9356 9276
rect 9412 9274 9418 9276
rect 9172 9222 9174 9274
rect 9354 9222 9356 9274
rect 9110 9220 9116 9222
rect 9172 9220 9196 9222
rect 9252 9220 9276 9222
rect 9332 9220 9356 9222
rect 9412 9220 9418 9222
rect 9110 9200 9418 9220
rect 9876 8974 9904 9318
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9864 8832 9916 8838
rect 10048 8832 10100 8838
rect 9864 8774 9916 8780
rect 10046 8800 10048 8809
rect 10100 8800 10102 8809
rect 4214 8732 4522 8752
rect 4214 8730 4220 8732
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4516 8730 4522 8732
rect 4276 8678 4278 8730
rect 4458 8678 4460 8730
rect 4214 8676 4220 8678
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4516 8676 4522 8678
rect 4214 8656 4522 8676
rect 7478 8732 7786 8752
rect 7478 8730 7484 8732
rect 7540 8730 7564 8732
rect 7620 8730 7644 8732
rect 7700 8730 7724 8732
rect 7780 8730 7786 8732
rect 7540 8678 7542 8730
rect 7722 8678 7724 8730
rect 7478 8676 7484 8678
rect 7540 8676 7564 8678
rect 7620 8676 7644 8678
rect 7700 8676 7724 8678
rect 7780 8676 7786 8678
rect 7478 8656 7786 8676
rect 9876 8498 9904 8774
rect 10046 8735 10102 8744
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 5846 8188 6154 8208
rect 5846 8186 5852 8188
rect 5908 8186 5932 8188
rect 5988 8186 6012 8188
rect 6068 8186 6092 8188
rect 6148 8186 6154 8188
rect 5908 8134 5910 8186
rect 6090 8134 6092 8186
rect 5846 8132 5852 8134
rect 5908 8132 5932 8134
rect 5988 8132 6012 8134
rect 6068 8132 6092 8134
rect 6148 8132 6154 8134
rect 5846 8112 6154 8132
rect 9110 8188 9418 8208
rect 9110 8186 9116 8188
rect 9172 8186 9196 8188
rect 9252 8186 9276 8188
rect 9332 8186 9356 8188
rect 9412 8186 9418 8188
rect 9172 8134 9174 8186
rect 9354 8134 9356 8186
rect 9110 8132 9116 8134
rect 9172 8132 9196 8134
rect 9252 8132 9276 8134
rect 9332 8132 9356 8134
rect 9412 8132 9418 8134
rect 9110 8112 9418 8132
rect 10060 7993 10088 8298
rect 10046 7984 10102 7993
rect 10046 7919 10102 7928
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 4214 7644 4522 7664
rect 4214 7642 4220 7644
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4516 7642 4522 7644
rect 4276 7590 4278 7642
rect 4458 7590 4460 7642
rect 4214 7588 4220 7590
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4516 7588 4522 7590
rect 4214 7568 4522 7588
rect 7478 7644 7786 7664
rect 7478 7642 7484 7644
rect 7540 7642 7564 7644
rect 7620 7642 7644 7644
rect 7700 7642 7724 7644
rect 7780 7642 7786 7644
rect 7540 7590 7542 7642
rect 7722 7590 7724 7642
rect 7478 7588 7484 7590
rect 7540 7588 7564 7590
rect 7620 7588 7644 7590
rect 7700 7588 7724 7590
rect 7780 7588 7786 7590
rect 7478 7568 7786 7588
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3896 5302 3924 5646
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3974 4856 4030 4865
rect 3974 4791 3976 4800
rect 4028 4791 4030 4800
rect 3976 4762 4028 4768
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 4080 4146 4108 7346
rect 5846 7100 6154 7120
rect 5846 7098 5852 7100
rect 5908 7098 5932 7100
rect 5988 7098 6012 7100
rect 6068 7098 6092 7100
rect 6148 7098 6154 7100
rect 5908 7046 5910 7098
rect 6090 7046 6092 7098
rect 5846 7044 5852 7046
rect 5908 7044 5932 7046
rect 5988 7044 6012 7046
rect 6068 7044 6092 7046
rect 6148 7044 6154 7046
rect 5846 7024 6154 7044
rect 9110 7100 9418 7120
rect 9110 7098 9116 7100
rect 9172 7098 9196 7100
rect 9252 7098 9276 7100
rect 9332 7098 9356 7100
rect 9412 7098 9418 7100
rect 9172 7046 9174 7098
rect 9354 7046 9356 7098
rect 9110 7044 9116 7046
rect 9172 7044 9196 7046
rect 9252 7044 9276 7046
rect 9332 7044 9356 7046
rect 9412 7044 9418 7046
rect 9110 7024 9418 7044
rect 9876 6798 9904 7686
rect 10048 7200 10100 7206
rect 10046 7168 10048 7177
rect 10100 7168 10102 7177
rect 10046 7103 10102 7112
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 4214 6556 4522 6576
rect 4214 6554 4220 6556
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4516 6554 4522 6556
rect 4276 6502 4278 6554
rect 4458 6502 4460 6554
rect 4214 6500 4220 6502
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4516 6500 4522 6502
rect 4214 6480 4522 6500
rect 7478 6556 7786 6576
rect 7478 6554 7484 6556
rect 7540 6554 7564 6556
rect 7620 6554 7644 6556
rect 7700 6554 7724 6556
rect 7780 6554 7786 6556
rect 7540 6502 7542 6554
rect 7722 6502 7724 6554
rect 7478 6500 7484 6502
rect 7540 6500 7564 6502
rect 7620 6500 7644 6502
rect 7700 6500 7724 6502
rect 7780 6500 7786 6502
rect 7478 6480 7786 6500
rect 5846 6012 6154 6032
rect 5846 6010 5852 6012
rect 5908 6010 5932 6012
rect 5988 6010 6012 6012
rect 6068 6010 6092 6012
rect 6148 6010 6154 6012
rect 5908 5958 5910 6010
rect 6090 5958 6092 6010
rect 5846 5956 5852 5958
rect 5908 5956 5932 5958
rect 5988 5956 6012 5958
rect 6068 5956 6092 5958
rect 6148 5956 6154 5958
rect 5846 5936 6154 5956
rect 9110 6012 9418 6032
rect 9110 6010 9116 6012
rect 9172 6010 9196 6012
rect 9252 6010 9276 6012
rect 9332 6010 9356 6012
rect 9412 6010 9418 6012
rect 9172 5958 9174 6010
rect 9354 5958 9356 6010
rect 9110 5956 9116 5958
rect 9172 5956 9196 5958
rect 9252 5956 9276 5958
rect 9332 5956 9356 5958
rect 9412 5956 9418 5958
rect 9110 5936 9418 5956
rect 9876 5710 9904 6598
rect 10060 6497 10088 6598
rect 10046 6488 10102 6497
rect 10046 6423 10102 6432
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 10046 5672 10102 5681
rect 10046 5607 10102 5616
rect 10060 5574 10088 5607
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 4214 5468 4522 5488
rect 4214 5466 4220 5468
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4516 5466 4522 5468
rect 4276 5414 4278 5466
rect 4458 5414 4460 5466
rect 4214 5412 4220 5414
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4516 5412 4522 5414
rect 4214 5392 4522 5412
rect 6840 5234 6868 5510
rect 7478 5468 7786 5488
rect 7478 5466 7484 5468
rect 7540 5466 7564 5468
rect 7620 5466 7644 5468
rect 7700 5466 7724 5468
rect 7780 5466 7786 5468
rect 7540 5414 7542 5466
rect 7722 5414 7724 5466
rect 7478 5412 7484 5414
rect 7540 5412 7564 5414
rect 7620 5412 7644 5414
rect 7700 5412 7724 5414
rect 7780 5412 7786 5414
rect 7478 5392 7786 5412
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4214 4380 4522 4400
rect 4214 4378 4220 4380
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4516 4378 4522 4380
rect 4276 4326 4278 4378
rect 4458 4326 4460 4378
rect 4214 4324 4220 4326
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4516 4324 4522 4326
rect 4214 4304 4522 4324
rect 4632 4146 4660 4490
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3620 3194 3648 3470
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3804 3058 3832 3878
rect 3988 3534 4016 4082
rect 4724 4078 4752 4558
rect 5184 4146 5212 5034
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 5846 4924 6154 4944
rect 5846 4922 5852 4924
rect 5908 4922 5932 4924
rect 5988 4922 6012 4924
rect 6068 4922 6092 4924
rect 6148 4922 6154 4924
rect 5908 4870 5910 4922
rect 6090 4870 6092 4922
rect 5846 4868 5852 4870
rect 5908 4868 5932 4870
rect 5988 4868 6012 4870
rect 6068 4868 6092 4870
rect 6148 4868 6154 4870
rect 5846 4848 6154 4868
rect 9110 4924 9418 4944
rect 9110 4922 9116 4924
rect 9172 4922 9196 4924
rect 9252 4922 9276 4924
rect 9332 4922 9356 4924
rect 9412 4922 9418 4924
rect 9172 4870 9174 4922
rect 9354 4870 9356 4922
rect 9110 4868 9116 4870
rect 9172 4868 9196 4870
rect 9252 4868 9276 4870
rect 9332 4868 9356 4870
rect 9412 4868 9418 4870
rect 9110 4848 9418 4868
rect 10060 4865 10088 4966
rect 10046 4856 10102 4865
rect 10046 4791 10102 4800
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 7478 4380 7786 4400
rect 7478 4378 7484 4380
rect 7540 4378 7564 4380
rect 7620 4378 7644 4380
rect 7700 4378 7724 4380
rect 7780 4378 7786 4380
rect 7540 4326 7542 4378
rect 7722 4326 7724 4378
rect 7478 4324 7484 4326
rect 7540 4324 7564 4326
rect 7620 4324 7644 4326
rect 7700 4324 7724 4326
rect 7780 4324 7786 4326
rect 7478 4304 7786 4324
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 4172 3602 4200 3946
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 4214 3292 4522 3312
rect 4214 3290 4220 3292
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4516 3290 4522 3292
rect 4276 3238 4278 3290
rect 4458 3238 4460 3290
rect 4214 3236 4220 3238
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4516 3236 4522 3238
rect 4214 3216 4522 3236
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 4066 2544 4122 2553
rect 4172 2530 4200 2926
rect 4122 2502 4200 2530
rect 4448 2514 4476 2994
rect 4632 2650 4660 3538
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4436 2508 4488 2514
rect 4066 2479 4122 2488
rect 4436 2450 4488 2456
rect 5644 2446 5672 3946
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 5846 3836 6154 3856
rect 5846 3834 5852 3836
rect 5908 3834 5932 3836
rect 5988 3834 6012 3836
rect 6068 3834 6092 3836
rect 6148 3834 6154 3836
rect 5908 3782 5910 3834
rect 6090 3782 6092 3834
rect 5846 3780 5852 3782
rect 5908 3780 5932 3782
rect 5988 3780 6012 3782
rect 6068 3780 6092 3782
rect 6148 3780 6154 3782
rect 5846 3760 6154 3780
rect 7478 3292 7786 3312
rect 7478 3290 7484 3292
rect 7540 3290 7564 3292
rect 7620 3290 7644 3292
rect 7700 3290 7724 3292
rect 7780 3290 7786 3292
rect 7540 3238 7542 3290
rect 7722 3238 7724 3290
rect 7478 3236 7484 3238
rect 7540 3236 7564 3238
rect 7620 3236 7644 3238
rect 7700 3236 7724 3238
rect 7780 3236 7786 3238
rect 7478 3216 7786 3236
rect 9048 3058 9076 3878
rect 9110 3836 9418 3856
rect 9110 3834 9116 3836
rect 9172 3834 9196 3836
rect 9252 3834 9276 3836
rect 9332 3834 9356 3836
rect 9412 3834 9418 3836
rect 9172 3782 9174 3834
rect 9354 3782 9356 3834
rect 9110 3780 9116 3782
rect 9172 3780 9196 3782
rect 9252 3780 9276 3782
rect 9332 3780 9356 3782
rect 9412 3780 9418 3782
rect 9110 3760 9418 3780
rect 9784 3534 9812 4422
rect 9876 4282 9904 4558
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 10060 4185 10088 4422
rect 10046 4176 10102 4185
rect 10046 4111 10102 4120
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10152 3738 10180 4082
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10048 3392 10100 3398
rect 10046 3360 10048 3369
rect 10100 3360 10102 3369
rect 10046 3295 10102 3304
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 5846 2748 6154 2768
rect 5846 2746 5852 2748
rect 5908 2746 5932 2748
rect 5988 2746 6012 2748
rect 6068 2746 6092 2748
rect 6148 2746 6154 2748
rect 5908 2694 5910 2746
rect 6090 2694 6092 2746
rect 5846 2692 5852 2694
rect 5908 2692 5932 2694
rect 5988 2692 6012 2694
rect 6068 2692 6092 2694
rect 6148 2692 6154 2694
rect 5846 2672 6154 2692
rect 9110 2748 9418 2768
rect 9110 2746 9116 2748
rect 9172 2746 9196 2748
rect 9252 2746 9276 2748
rect 9332 2746 9356 2748
rect 9412 2746 9418 2748
rect 9172 2694 9174 2746
rect 9354 2694 9356 2746
rect 9110 2692 9116 2694
rect 9172 2692 9196 2694
rect 9252 2692 9276 2694
rect 9332 2692 9356 2694
rect 9412 2692 9418 2694
rect 9110 2672 9418 2692
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 3988 1465 4016 2382
rect 4080 1873 4108 2382
rect 4214 2204 4522 2224
rect 4214 2202 4220 2204
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4516 2202 4522 2204
rect 4276 2150 4278 2202
rect 4458 2150 4460 2202
rect 4214 2148 4220 2150
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4516 2148 4522 2150
rect 4214 2128 4522 2148
rect 4066 1864 4122 1873
rect 4066 1799 4122 1808
rect 3974 1456 4030 1465
rect 3974 1391 4030 1400
rect 5276 1086 5304 2382
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 7478 2204 7786 2224
rect 7478 2202 7484 2204
rect 7540 2202 7564 2204
rect 7620 2202 7644 2204
rect 7700 2202 7724 2204
rect 7780 2202 7786 2204
rect 7540 2150 7542 2202
rect 7722 2150 7724 2202
rect 7478 2148 7484 2150
rect 7540 2148 7564 2150
rect 7620 2148 7644 2150
rect 7700 2148 7724 2150
rect 7780 2148 7786 2150
rect 7478 2128 7786 2148
rect 5264 1080 5316 1086
rect 5264 1022 5316 1028
rect 2870 640 2926 649
rect 2870 575 2926 584
rect 1398 232 1454 241
rect 1398 167 1454 176
rect 5998 0 6054 800
rect 9324 377 9352 2246
rect 9508 1873 9536 2790
rect 9692 2446 9720 3062
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10060 2553 10088 2790
rect 10046 2544 10102 2553
rect 10046 2479 10102 2488
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9494 1864 9550 1873
rect 9494 1799 9550 1808
rect 9600 1057 9628 2246
rect 9586 1048 9642 1057
rect 9586 983 9642 992
rect 9310 368 9366 377
rect 9310 303 9366 312
<< via2 >>
rect 2962 79600 3018 79656
rect 1398 79192 1454 79248
rect 2588 77818 2644 77820
rect 2668 77818 2724 77820
rect 2748 77818 2804 77820
rect 2828 77818 2884 77820
rect 2588 77766 2634 77818
rect 2634 77766 2644 77818
rect 2668 77766 2698 77818
rect 2698 77766 2710 77818
rect 2710 77766 2724 77818
rect 2748 77766 2762 77818
rect 2762 77766 2774 77818
rect 2774 77766 2804 77818
rect 2828 77766 2838 77818
rect 2838 77766 2884 77818
rect 2588 77764 2644 77766
rect 2668 77764 2724 77766
rect 2748 77764 2804 77766
rect 2828 77764 2884 77766
rect 9954 79464 10010 79520
rect 3698 78784 3754 78840
rect 3422 77968 3478 78024
rect 1398 74976 1454 75032
rect 110 50380 166 50416
rect 110 50360 112 50380
rect 112 50360 164 50380
rect 164 50360 166 50380
rect 110 46572 166 46574
rect 110 46520 112 46572
rect 112 46520 164 46572
rect 164 46520 166 46572
rect 110 46518 166 46520
rect 1582 74568 1638 74624
rect 1122 72700 1124 72720
rect 1124 72700 1176 72720
rect 1176 72700 1178 72720
rect 1122 72664 1178 72700
rect 1398 72800 1454 72856
rect 1582 72392 1638 72448
rect 1582 71032 1638 71088
rect 1582 70624 1638 70680
rect 1582 70216 1638 70272
rect 1306 67632 1362 67688
rect 1398 67224 1454 67280
rect 1398 66816 1454 66872
rect 1582 68040 1638 68096
rect 478 53352 534 53408
rect 294 44376 350 44432
rect 938 60560 994 60616
rect 754 32816 810 32872
rect 1674 67668 1676 67688
rect 1676 67668 1728 67688
rect 1728 67668 1730 67688
rect 1674 67632 1730 67668
rect 1582 66156 1638 66192
rect 1582 66136 1584 66156
rect 1584 66136 1636 66156
rect 1636 66136 1638 66156
rect 1582 66000 1638 66056
rect 1490 64912 1546 64968
rect 1398 62056 1454 62112
rect 1674 63452 1676 63472
rect 1676 63452 1728 63472
rect 1728 63452 1730 63472
rect 1674 63416 1730 63452
rect 1582 63008 1638 63064
rect 1122 58928 1178 58984
rect 1122 58792 1178 58848
rect 1674 62192 1730 62248
rect 1582 61376 1638 61432
rect 1766 61240 1822 61296
rect 1398 57432 1454 57488
rect 1122 56344 1178 56400
rect 1306 55140 1362 55176
rect 1306 55120 1308 55140
rect 1308 55120 1360 55140
rect 1360 55120 1362 55140
rect 1582 59064 1638 59120
rect 1582 57024 1638 57080
rect 1674 56616 1730 56672
rect 1582 55392 1638 55448
rect 1766 55392 1822 55448
rect 1766 54304 1822 54360
rect 1490 54032 1546 54088
rect 1398 52672 1454 52728
rect 1306 51584 1362 51640
rect 1306 51176 1362 51232
rect 1214 50904 1270 50960
rect 1122 50632 1178 50688
rect 1122 49836 1178 49872
rect 1122 49816 1124 49836
rect 1124 49816 1176 49836
rect 1176 49816 1178 49836
rect 1122 48320 1178 48376
rect 1030 41384 1086 41440
rect 938 38528 994 38584
rect 938 36896 994 36952
rect 1122 39208 1178 39264
rect 1122 38664 1178 38720
rect 1398 50904 1454 50960
rect 1582 52264 1638 52320
rect 1582 52148 1638 52184
rect 1582 52128 1584 52148
rect 1584 52128 1636 52148
rect 1636 52128 1638 52148
rect 1766 51312 1822 51368
rect 1766 51176 1822 51232
rect 1674 51040 1730 51096
rect 1674 50360 1730 50416
rect 1490 50224 1546 50280
rect 1398 48456 1454 48512
rect 1582 48048 1638 48104
rect 1582 47640 1638 47696
rect 1398 47368 1454 47424
rect 1398 46552 1454 46608
rect 1398 45600 1454 45656
rect 1766 48184 1822 48240
rect 1674 46824 1730 46880
rect 1490 45328 1546 45384
rect 1398 44240 1454 44296
rect 1582 45076 1638 45112
rect 1582 45056 1584 45076
rect 1584 45056 1636 45076
rect 1636 45056 1638 45076
rect 1582 44648 1638 44704
rect 1306 42744 1362 42800
rect 1582 44104 1638 44160
rect 1490 43016 1546 43072
rect 1306 41556 1308 41576
rect 1308 41556 1360 41576
rect 1360 41556 1362 41576
rect 1306 41520 1362 41556
rect 1306 41384 1362 41440
rect 1398 39344 1454 39400
rect 1306 38800 1362 38856
rect 1306 38528 1362 38584
rect 2042 69808 2098 69864
rect 1950 60968 2006 61024
rect 2226 73208 2282 73264
rect 2226 71576 2282 71632
rect 2226 68992 2282 69048
rect 2226 67360 2282 67416
rect 2962 77016 3018 77072
rect 2588 76730 2644 76732
rect 2668 76730 2724 76732
rect 2748 76730 2804 76732
rect 2828 76730 2884 76732
rect 2588 76678 2634 76730
rect 2634 76678 2644 76730
rect 2668 76678 2698 76730
rect 2698 76678 2710 76730
rect 2710 76678 2724 76730
rect 2748 76678 2762 76730
rect 2762 76678 2774 76730
rect 2774 76678 2804 76730
rect 2828 76678 2838 76730
rect 2838 76678 2884 76730
rect 2588 76676 2644 76678
rect 2668 76676 2724 76678
rect 2748 76676 2804 76678
rect 2828 76676 2884 76678
rect 2502 75792 2558 75848
rect 2588 75642 2644 75644
rect 2668 75642 2724 75644
rect 2748 75642 2804 75644
rect 2828 75642 2884 75644
rect 2588 75590 2634 75642
rect 2634 75590 2644 75642
rect 2668 75590 2698 75642
rect 2698 75590 2710 75642
rect 2710 75590 2724 75642
rect 2748 75590 2762 75642
rect 2762 75590 2774 75642
rect 2774 75590 2804 75642
rect 2828 75590 2838 75642
rect 2838 75590 2884 75642
rect 2588 75588 2644 75590
rect 2668 75588 2724 75590
rect 2748 75588 2804 75590
rect 2828 75588 2884 75590
rect 2502 74976 2558 75032
rect 2588 74554 2644 74556
rect 2668 74554 2724 74556
rect 2748 74554 2804 74556
rect 2828 74554 2884 74556
rect 2588 74502 2634 74554
rect 2634 74502 2644 74554
rect 2668 74502 2698 74554
rect 2698 74502 2710 74554
rect 2710 74502 2724 74554
rect 2748 74502 2762 74554
rect 2762 74502 2774 74554
rect 2774 74502 2804 74554
rect 2828 74502 2838 74554
rect 2838 74502 2884 74554
rect 2588 74500 2644 74502
rect 2668 74500 2724 74502
rect 2748 74500 2804 74502
rect 2828 74500 2884 74502
rect 2962 74024 3018 74080
rect 2870 73616 2926 73672
rect 2588 73466 2644 73468
rect 2668 73466 2724 73468
rect 2748 73466 2804 73468
rect 2828 73466 2884 73468
rect 2588 73414 2634 73466
rect 2634 73414 2644 73466
rect 2668 73414 2698 73466
rect 2698 73414 2710 73466
rect 2710 73414 2724 73466
rect 2748 73414 2762 73466
rect 2762 73414 2774 73466
rect 2774 73414 2804 73466
rect 2828 73414 2838 73466
rect 2838 73414 2884 73466
rect 2588 73412 2644 73414
rect 2668 73412 2724 73414
rect 2748 73412 2804 73414
rect 2828 73412 2884 73414
rect 2686 72684 2742 72720
rect 2686 72664 2688 72684
rect 2688 72664 2740 72684
rect 2740 72664 2742 72684
rect 2588 72378 2644 72380
rect 2668 72378 2724 72380
rect 2748 72378 2804 72380
rect 2828 72378 2884 72380
rect 2588 72326 2634 72378
rect 2634 72326 2644 72378
rect 2668 72326 2698 72378
rect 2698 72326 2710 72378
rect 2710 72326 2724 72378
rect 2748 72326 2762 72378
rect 2762 72326 2774 72378
rect 2774 72326 2804 72378
rect 2828 72326 2838 72378
rect 2838 72326 2884 72378
rect 2588 72324 2644 72326
rect 2668 72324 2724 72326
rect 2748 72324 2804 72326
rect 2828 72324 2884 72326
rect 2870 72020 2872 72040
rect 2872 72020 2924 72040
rect 2924 72020 2926 72040
rect 2870 71984 2926 72020
rect 2588 71290 2644 71292
rect 2668 71290 2724 71292
rect 2748 71290 2804 71292
rect 2828 71290 2884 71292
rect 2588 71238 2634 71290
rect 2634 71238 2644 71290
rect 2668 71238 2698 71290
rect 2698 71238 2710 71290
rect 2710 71238 2724 71290
rect 2748 71238 2762 71290
rect 2762 71238 2774 71290
rect 2774 71238 2804 71290
rect 2828 71238 2838 71290
rect 2838 71238 2884 71290
rect 2588 71236 2644 71238
rect 2668 71236 2724 71238
rect 2748 71236 2804 71238
rect 2828 71236 2884 71238
rect 2588 70202 2644 70204
rect 2668 70202 2724 70204
rect 2748 70202 2804 70204
rect 2828 70202 2884 70204
rect 2588 70150 2634 70202
rect 2634 70150 2644 70202
rect 2668 70150 2698 70202
rect 2698 70150 2710 70202
rect 2710 70150 2724 70202
rect 2748 70150 2762 70202
rect 2762 70150 2774 70202
rect 2774 70150 2804 70202
rect 2828 70150 2838 70202
rect 2838 70150 2884 70202
rect 2588 70148 2644 70150
rect 2668 70148 2724 70150
rect 2748 70148 2804 70150
rect 2828 70148 2884 70150
rect 3330 76472 3386 76528
rect 9586 78648 9642 78704
rect 4066 78376 4122 78432
rect 3974 77560 4030 77616
rect 9494 77968 9550 78024
rect 5852 77818 5908 77820
rect 5932 77818 5988 77820
rect 6012 77818 6068 77820
rect 6092 77818 6148 77820
rect 5852 77766 5898 77818
rect 5898 77766 5908 77818
rect 5932 77766 5962 77818
rect 5962 77766 5974 77818
rect 5974 77766 5988 77818
rect 6012 77766 6026 77818
rect 6026 77766 6038 77818
rect 6038 77766 6068 77818
rect 6092 77766 6102 77818
rect 6102 77766 6148 77818
rect 5852 77764 5908 77766
rect 5932 77764 5988 77766
rect 6012 77764 6068 77766
rect 6092 77764 6148 77766
rect 9116 77818 9172 77820
rect 9196 77818 9252 77820
rect 9276 77818 9332 77820
rect 9356 77818 9412 77820
rect 9116 77766 9162 77818
rect 9162 77766 9172 77818
rect 9196 77766 9226 77818
rect 9226 77766 9238 77818
rect 9238 77766 9252 77818
rect 9276 77766 9290 77818
rect 9290 77766 9302 77818
rect 9302 77766 9332 77818
rect 9356 77766 9366 77818
rect 9366 77766 9412 77818
rect 9116 77764 9172 77766
rect 9196 77764 9252 77766
rect 9276 77764 9332 77766
rect 9356 77764 9412 77766
rect 2870 69400 2926 69456
rect 2686 69264 2742 69320
rect 2588 69114 2644 69116
rect 2668 69114 2724 69116
rect 2748 69114 2804 69116
rect 2828 69114 2884 69116
rect 2588 69062 2634 69114
rect 2634 69062 2644 69114
rect 2668 69062 2698 69114
rect 2698 69062 2710 69114
rect 2710 69062 2724 69114
rect 2748 69062 2762 69114
rect 2762 69062 2774 69114
rect 2774 69062 2804 69114
rect 2828 69062 2838 69114
rect 2838 69062 2884 69114
rect 2588 69060 2644 69062
rect 2668 69060 2724 69062
rect 2748 69060 2804 69062
rect 2828 69060 2884 69062
rect 2226 64096 2282 64152
rect 2318 62636 2320 62656
rect 2320 62636 2372 62656
rect 2372 62636 2374 62656
rect 2318 62600 2374 62636
rect 2962 68584 3018 68640
rect 2588 68026 2644 68028
rect 2668 68026 2724 68028
rect 2748 68026 2804 68028
rect 2828 68026 2884 68028
rect 2588 67974 2634 68026
rect 2634 67974 2644 68026
rect 2668 67974 2698 68026
rect 2698 67974 2710 68026
rect 2710 67974 2724 68026
rect 2748 67974 2762 68026
rect 2762 67974 2774 68026
rect 2774 67974 2804 68026
rect 2828 67974 2838 68026
rect 2838 67974 2884 68026
rect 2588 67972 2644 67974
rect 2668 67972 2724 67974
rect 2748 67972 2804 67974
rect 2828 67972 2884 67974
rect 2588 66938 2644 66940
rect 2668 66938 2724 66940
rect 2748 66938 2804 66940
rect 2828 66938 2884 66940
rect 2588 66886 2634 66938
rect 2634 66886 2644 66938
rect 2668 66886 2698 66938
rect 2698 66886 2710 66938
rect 2710 66886 2724 66938
rect 2748 66886 2762 66938
rect 2762 66886 2774 66938
rect 2774 66886 2804 66938
rect 2828 66886 2838 66938
rect 2838 66886 2884 66938
rect 2588 66884 2644 66886
rect 2668 66884 2724 66886
rect 2748 66884 2804 66886
rect 2828 66884 2884 66886
rect 2318 60696 2374 60752
rect 2318 60016 2374 60072
rect 2318 59880 2374 59936
rect 2588 65850 2644 65852
rect 2668 65850 2724 65852
rect 2748 65850 2804 65852
rect 2828 65850 2884 65852
rect 2588 65798 2634 65850
rect 2634 65798 2644 65850
rect 2668 65798 2698 65850
rect 2698 65798 2710 65850
rect 2710 65798 2724 65850
rect 2748 65798 2762 65850
rect 2762 65798 2774 65850
rect 2774 65798 2804 65850
rect 2828 65798 2838 65850
rect 2838 65798 2884 65850
rect 2588 65796 2644 65798
rect 2668 65796 2724 65798
rect 2748 65796 2804 65798
rect 2828 65796 2884 65798
rect 3054 66408 3110 66464
rect 2962 65592 3018 65648
rect 2588 64762 2644 64764
rect 2668 64762 2724 64764
rect 2748 64762 2804 64764
rect 2828 64762 2884 64764
rect 2588 64710 2634 64762
rect 2634 64710 2644 64762
rect 2668 64710 2698 64762
rect 2698 64710 2710 64762
rect 2710 64710 2724 64762
rect 2748 64710 2762 64762
rect 2762 64710 2774 64762
rect 2774 64710 2804 64762
rect 2828 64710 2838 64762
rect 2838 64710 2884 64762
rect 2588 64708 2644 64710
rect 2668 64708 2724 64710
rect 2748 64708 2804 64710
rect 2828 64708 2884 64710
rect 3054 64504 3110 64560
rect 3054 64268 3056 64288
rect 3056 64268 3108 64288
rect 3108 64268 3110 64288
rect 3054 64232 3110 64268
rect 2588 63674 2644 63676
rect 2668 63674 2724 63676
rect 2748 63674 2804 63676
rect 2828 63674 2884 63676
rect 2588 63622 2634 63674
rect 2634 63622 2644 63674
rect 2668 63622 2698 63674
rect 2698 63622 2710 63674
rect 2710 63622 2724 63674
rect 2748 63622 2762 63674
rect 2762 63622 2774 63674
rect 2774 63622 2804 63674
rect 2828 63622 2838 63674
rect 2838 63622 2884 63674
rect 2588 63620 2644 63622
rect 2668 63620 2724 63622
rect 2748 63620 2804 63622
rect 2828 63620 2884 63622
rect 2870 62872 2926 62928
rect 2588 62586 2644 62588
rect 2668 62586 2724 62588
rect 2748 62586 2804 62588
rect 2828 62586 2884 62588
rect 2588 62534 2634 62586
rect 2634 62534 2644 62586
rect 2668 62534 2698 62586
rect 2698 62534 2710 62586
rect 2710 62534 2724 62586
rect 2748 62534 2762 62586
rect 2762 62534 2774 62586
rect 2774 62534 2804 62586
rect 2828 62534 2838 62586
rect 2838 62534 2884 62586
rect 2588 62532 2644 62534
rect 2668 62532 2724 62534
rect 2748 62532 2804 62534
rect 2828 62532 2884 62534
rect 3054 63824 3110 63880
rect 2686 61804 2742 61840
rect 2686 61784 2688 61804
rect 2688 61784 2740 61804
rect 2740 61784 2742 61804
rect 2588 61498 2644 61500
rect 2668 61498 2724 61500
rect 2748 61498 2804 61500
rect 2828 61498 2884 61500
rect 2588 61446 2634 61498
rect 2634 61446 2644 61498
rect 2668 61446 2698 61498
rect 2698 61446 2710 61498
rect 2710 61446 2724 61498
rect 2748 61446 2762 61498
rect 2762 61446 2774 61498
rect 2774 61446 2804 61498
rect 2828 61446 2838 61498
rect 2838 61446 2884 61498
rect 2588 61444 2644 61446
rect 2668 61444 2724 61446
rect 2748 61444 2804 61446
rect 2828 61444 2884 61446
rect 2502 60968 2558 61024
rect 2778 60832 2834 60888
rect 2962 60696 3018 60752
rect 2962 60580 3018 60616
rect 2962 60560 2964 60580
rect 2964 60560 3016 60580
rect 3016 60560 3018 60580
rect 2588 60410 2644 60412
rect 2668 60410 2724 60412
rect 2748 60410 2804 60412
rect 2828 60410 2884 60412
rect 2588 60358 2634 60410
rect 2634 60358 2644 60410
rect 2668 60358 2698 60410
rect 2698 60358 2710 60410
rect 2710 60358 2724 60410
rect 2748 60358 2762 60410
rect 2762 60358 2774 60410
rect 2774 60358 2804 60410
rect 2828 60358 2838 60410
rect 2838 60358 2884 60410
rect 2588 60356 2644 60358
rect 2668 60356 2724 60358
rect 2748 60356 2804 60358
rect 2828 60356 2884 60358
rect 2134 59472 2190 59528
rect 1950 57432 2006 57488
rect 2226 58792 2282 58848
rect 2042 53624 2098 53680
rect 1766 42336 1822 42392
rect 1950 42880 2006 42936
rect 1950 42744 2006 42800
rect 1858 41792 1914 41848
rect 1674 41384 1730 41440
rect 1582 38528 1638 38584
rect 1582 38392 1638 38448
rect 1306 38256 1362 38312
rect 1490 38256 1546 38312
rect 1122 31320 1178 31376
rect 1122 30268 1124 30288
rect 1124 30268 1176 30288
rect 1176 30268 1178 30288
rect 1122 30232 1178 30268
rect 1214 27920 1270 27976
rect 1214 22752 1270 22808
rect 1214 21936 1270 21992
rect 1582 36080 1638 36136
rect 1582 35128 1638 35184
rect 1398 33496 1454 33552
rect 1582 34740 1638 34776
rect 1582 34720 1584 34740
rect 1584 34720 1636 34740
rect 1636 34720 1638 34740
rect 1490 33224 1546 33280
rect 1490 32816 1546 32872
rect 1398 31864 1454 31920
rect 1674 32136 1730 32192
rect 1490 31456 1546 31512
rect 1398 27512 1454 27568
rect 1398 25336 1454 25392
rect 1398 24928 1454 24984
rect 1398 23160 1454 23216
rect 1398 22344 1454 22400
rect 1398 21528 1454 21584
rect 1398 21120 1454 21176
rect 2410 57568 2466 57624
rect 2318 55664 2374 55720
rect 2318 55256 2374 55312
rect 2318 53080 2374 53136
rect 2134 52672 2190 52728
rect 2134 51176 2190 51232
rect 2134 50768 2190 50824
rect 2778 59608 2834 59664
rect 2594 59472 2650 59528
rect 2588 59322 2644 59324
rect 2668 59322 2724 59324
rect 2748 59322 2804 59324
rect 2828 59322 2884 59324
rect 2588 59270 2634 59322
rect 2634 59270 2644 59322
rect 2668 59270 2698 59322
rect 2698 59270 2710 59322
rect 2710 59270 2724 59322
rect 2748 59270 2762 59322
rect 2762 59270 2774 59322
rect 2774 59270 2804 59322
rect 2828 59270 2838 59322
rect 2838 59270 2884 59322
rect 2588 59268 2644 59270
rect 2668 59268 2724 59270
rect 2748 59268 2804 59270
rect 2828 59268 2884 59270
rect 2686 58540 2742 58576
rect 2686 58520 2688 58540
rect 2688 58520 2740 58540
rect 2740 58520 2742 58540
rect 2588 58234 2644 58236
rect 2668 58234 2724 58236
rect 2748 58234 2804 58236
rect 2828 58234 2884 58236
rect 2588 58182 2634 58234
rect 2634 58182 2644 58234
rect 2668 58182 2698 58234
rect 2698 58182 2710 58234
rect 2710 58182 2724 58234
rect 2748 58182 2762 58234
rect 2762 58182 2774 58234
rect 2774 58182 2804 58234
rect 2828 58182 2838 58234
rect 2838 58182 2884 58234
rect 2588 58180 2644 58182
rect 2668 58180 2724 58182
rect 2748 58180 2804 58182
rect 2828 58180 2884 58182
rect 2594 57840 2650 57896
rect 2686 57296 2742 57352
rect 2588 57146 2644 57148
rect 2668 57146 2724 57148
rect 2748 57146 2804 57148
rect 2828 57146 2884 57148
rect 2588 57094 2634 57146
rect 2634 57094 2644 57146
rect 2668 57094 2698 57146
rect 2698 57094 2710 57146
rect 2710 57094 2724 57146
rect 2748 57094 2762 57146
rect 2762 57094 2774 57146
rect 2774 57094 2804 57146
rect 2828 57094 2838 57146
rect 2838 57094 2884 57146
rect 2588 57092 2644 57094
rect 2668 57092 2724 57094
rect 2748 57092 2804 57094
rect 2828 57092 2884 57094
rect 2686 56228 2742 56264
rect 2686 56208 2688 56228
rect 2688 56208 2740 56228
rect 2740 56208 2742 56228
rect 2588 56058 2644 56060
rect 2668 56058 2724 56060
rect 2748 56058 2804 56060
rect 2828 56058 2884 56060
rect 2588 56006 2634 56058
rect 2634 56006 2644 56058
rect 2668 56006 2698 56058
rect 2698 56006 2710 56058
rect 2710 56006 2724 56058
rect 2748 56006 2762 56058
rect 2762 56006 2774 56058
rect 2774 56006 2804 56058
rect 2828 56006 2838 56058
rect 2838 56006 2884 56058
rect 2588 56004 2644 56006
rect 2668 56004 2724 56006
rect 2748 56004 2804 56006
rect 2828 56004 2884 56006
rect 2870 55700 2872 55720
rect 2872 55700 2924 55720
rect 2924 55700 2926 55720
rect 2870 55664 2926 55700
rect 3054 60288 3110 60344
rect 3054 55256 3110 55312
rect 3238 63416 3294 63472
rect 3238 60832 3294 60888
rect 3238 60716 3294 60752
rect 3238 60696 3240 60716
rect 3240 60696 3292 60716
rect 3292 60696 3294 60716
rect 2588 54970 2644 54972
rect 2668 54970 2724 54972
rect 2748 54970 2804 54972
rect 2828 54970 2884 54972
rect 2588 54918 2634 54970
rect 2634 54918 2644 54970
rect 2668 54918 2698 54970
rect 2698 54918 2710 54970
rect 2710 54918 2724 54970
rect 2748 54918 2762 54970
rect 2762 54918 2774 54970
rect 2774 54918 2804 54970
rect 2828 54918 2838 54970
rect 2838 54918 2884 54970
rect 2588 54916 2644 54918
rect 2668 54916 2724 54918
rect 2748 54916 2804 54918
rect 2828 54916 2884 54918
rect 2778 54476 2780 54496
rect 2780 54476 2832 54496
rect 2832 54476 2834 54496
rect 2778 54440 2834 54476
rect 2588 53882 2644 53884
rect 2668 53882 2724 53884
rect 2748 53882 2804 53884
rect 2828 53882 2884 53884
rect 2588 53830 2634 53882
rect 2634 53830 2644 53882
rect 2668 53830 2698 53882
rect 2698 53830 2710 53882
rect 2710 53830 2724 53882
rect 2748 53830 2762 53882
rect 2762 53830 2774 53882
rect 2774 53830 2804 53882
rect 2828 53830 2838 53882
rect 2838 53830 2884 53882
rect 2588 53828 2644 53830
rect 2668 53828 2724 53830
rect 2748 53828 2804 53830
rect 2828 53828 2884 53830
rect 2594 52944 2650 53000
rect 2588 52794 2644 52796
rect 2668 52794 2724 52796
rect 2748 52794 2804 52796
rect 2828 52794 2884 52796
rect 2588 52742 2634 52794
rect 2634 52742 2644 52794
rect 2668 52742 2698 52794
rect 2698 52742 2710 52794
rect 2710 52742 2724 52794
rect 2748 52742 2762 52794
rect 2762 52742 2774 52794
rect 2774 52742 2804 52794
rect 2828 52742 2838 52794
rect 2838 52742 2884 52794
rect 2588 52740 2644 52742
rect 2668 52740 2724 52742
rect 2748 52740 2804 52742
rect 2828 52740 2884 52742
rect 2870 51856 2926 51912
rect 2588 51706 2644 51708
rect 2668 51706 2724 51708
rect 2748 51706 2804 51708
rect 2828 51706 2884 51708
rect 2588 51654 2634 51706
rect 2634 51654 2644 51706
rect 2668 51654 2698 51706
rect 2698 51654 2710 51706
rect 2710 51654 2724 51706
rect 2748 51654 2762 51706
rect 2762 51654 2774 51706
rect 2774 51654 2804 51706
rect 2828 51654 2838 51706
rect 2838 51654 2884 51706
rect 2588 51652 2644 51654
rect 2668 51652 2724 51654
rect 2748 51652 2804 51654
rect 2828 51652 2884 51654
rect 2588 50618 2644 50620
rect 2668 50618 2724 50620
rect 2748 50618 2804 50620
rect 2828 50618 2884 50620
rect 2588 50566 2634 50618
rect 2634 50566 2644 50618
rect 2668 50566 2698 50618
rect 2698 50566 2710 50618
rect 2710 50566 2724 50618
rect 2748 50566 2762 50618
rect 2762 50566 2774 50618
rect 2774 50566 2804 50618
rect 2828 50566 2838 50618
rect 2838 50566 2884 50618
rect 2588 50564 2644 50566
rect 2668 50564 2724 50566
rect 2748 50564 2804 50566
rect 2828 50564 2884 50566
rect 2962 50088 3018 50144
rect 2778 49680 2834 49736
rect 2588 49530 2644 49532
rect 2668 49530 2724 49532
rect 2748 49530 2804 49532
rect 2828 49530 2884 49532
rect 2588 49478 2634 49530
rect 2634 49478 2644 49530
rect 2668 49478 2698 49530
rect 2698 49478 2710 49530
rect 2710 49478 2724 49530
rect 2748 49478 2762 49530
rect 2762 49478 2774 49530
rect 2774 49478 2804 49530
rect 2828 49478 2838 49530
rect 2838 49478 2884 49530
rect 2588 49476 2644 49478
rect 2668 49476 2724 49478
rect 2748 49476 2804 49478
rect 2828 49476 2884 49478
rect 2502 49272 2558 49328
rect 2318 48864 2374 48920
rect 2594 49136 2650 49192
rect 2502 49000 2558 49056
rect 2778 49272 2834 49328
rect 2870 49136 2926 49192
rect 2410 48184 2466 48240
rect 2410 47912 2466 47968
rect 2962 48628 2964 48648
rect 2964 48628 3016 48648
rect 3016 48628 3018 48648
rect 2962 48592 3018 48628
rect 2588 48442 2644 48444
rect 2668 48442 2724 48444
rect 2748 48442 2804 48444
rect 2828 48442 2884 48444
rect 2588 48390 2634 48442
rect 2634 48390 2644 48442
rect 2668 48390 2698 48442
rect 2698 48390 2710 48442
rect 2710 48390 2724 48442
rect 2748 48390 2762 48442
rect 2762 48390 2774 48442
rect 2774 48390 2804 48442
rect 2828 48390 2838 48442
rect 2838 48390 2884 48442
rect 2588 48388 2644 48390
rect 2668 48388 2724 48390
rect 2748 48388 2804 48390
rect 2828 48388 2884 48390
rect 2778 48220 2780 48240
rect 2780 48220 2832 48240
rect 2832 48220 2834 48240
rect 2778 48184 2834 48220
rect 2686 47776 2742 47832
rect 2588 47354 2644 47356
rect 2668 47354 2724 47356
rect 2748 47354 2804 47356
rect 2828 47354 2884 47356
rect 2588 47302 2634 47354
rect 2634 47302 2644 47354
rect 2668 47302 2698 47354
rect 2698 47302 2710 47354
rect 2710 47302 2724 47354
rect 2748 47302 2762 47354
rect 2762 47302 2774 47354
rect 2774 47302 2804 47354
rect 2828 47302 2838 47354
rect 2838 47302 2884 47354
rect 2588 47300 2644 47302
rect 2668 47300 2724 47302
rect 2748 47300 2804 47302
rect 2828 47300 2884 47302
rect 2588 46266 2644 46268
rect 2668 46266 2724 46268
rect 2748 46266 2804 46268
rect 2828 46266 2884 46268
rect 2588 46214 2634 46266
rect 2634 46214 2644 46266
rect 2668 46214 2698 46266
rect 2698 46214 2710 46266
rect 2710 46214 2724 46266
rect 2748 46214 2762 46266
rect 2762 46214 2774 46266
rect 2774 46214 2804 46266
rect 2828 46214 2838 46266
rect 2838 46214 2884 46266
rect 2588 46212 2644 46214
rect 2668 46212 2724 46214
rect 2748 46212 2804 46214
rect 2828 46212 2884 46214
rect 2686 46008 2742 46064
rect 2870 45872 2926 45928
rect 2870 45600 2926 45656
rect 2588 45178 2644 45180
rect 2668 45178 2724 45180
rect 2748 45178 2804 45180
rect 2828 45178 2884 45180
rect 2588 45126 2634 45178
rect 2634 45126 2644 45178
rect 2668 45126 2698 45178
rect 2698 45126 2710 45178
rect 2710 45126 2724 45178
rect 2748 45126 2762 45178
rect 2762 45126 2774 45178
rect 2774 45126 2804 45178
rect 2828 45126 2838 45178
rect 2838 45126 2884 45178
rect 2588 45124 2644 45126
rect 2668 45124 2724 45126
rect 2748 45124 2804 45126
rect 2828 45124 2884 45126
rect 3238 51584 3294 51640
rect 3146 50904 3202 50960
rect 3146 49000 3202 49056
rect 3146 47640 3202 47696
rect 2588 44090 2644 44092
rect 2668 44090 2724 44092
rect 2748 44090 2804 44092
rect 2828 44090 2884 44092
rect 2588 44038 2634 44090
rect 2634 44038 2644 44090
rect 2668 44038 2698 44090
rect 2698 44038 2710 44090
rect 2710 44038 2724 44090
rect 2748 44038 2762 44090
rect 2762 44038 2774 44090
rect 2774 44038 2804 44090
rect 2828 44038 2838 44090
rect 2838 44038 2884 44090
rect 2588 44036 2644 44038
rect 2668 44036 2724 44038
rect 2748 44036 2804 44038
rect 2828 44036 2884 44038
rect 2226 38936 2282 38992
rect 2686 43832 2742 43888
rect 3698 75384 3754 75440
rect 4220 77274 4276 77276
rect 4300 77274 4356 77276
rect 4380 77274 4436 77276
rect 4460 77274 4516 77276
rect 4220 77222 4266 77274
rect 4266 77222 4276 77274
rect 4300 77222 4330 77274
rect 4330 77222 4342 77274
rect 4342 77222 4356 77274
rect 4380 77222 4394 77274
rect 4394 77222 4406 77274
rect 4406 77222 4436 77274
rect 4460 77222 4470 77274
rect 4470 77222 4516 77274
rect 4220 77220 4276 77222
rect 4300 77220 4356 77222
rect 4380 77220 4436 77222
rect 4460 77220 4516 77222
rect 7484 77274 7540 77276
rect 7564 77274 7620 77276
rect 7644 77274 7700 77276
rect 7724 77274 7780 77276
rect 7484 77222 7530 77274
rect 7530 77222 7540 77274
rect 7564 77222 7594 77274
rect 7594 77222 7606 77274
rect 7606 77222 7620 77274
rect 7644 77222 7658 77274
rect 7658 77222 7670 77274
rect 7670 77222 7700 77274
rect 7724 77222 7734 77274
rect 7734 77222 7780 77274
rect 7484 77220 7540 77222
rect 7564 77220 7620 77222
rect 7644 77220 7700 77222
rect 7724 77220 7780 77222
rect 5852 76730 5908 76732
rect 5932 76730 5988 76732
rect 6012 76730 6068 76732
rect 6092 76730 6148 76732
rect 5852 76678 5898 76730
rect 5898 76678 5908 76730
rect 5932 76678 5962 76730
rect 5962 76678 5974 76730
rect 5974 76678 5988 76730
rect 6012 76678 6026 76730
rect 6026 76678 6038 76730
rect 6038 76678 6068 76730
rect 6092 76678 6102 76730
rect 6102 76678 6148 76730
rect 5852 76676 5908 76678
rect 5932 76676 5988 76678
rect 6012 76676 6068 76678
rect 6092 76676 6148 76678
rect 3974 76200 4030 76256
rect 4220 76186 4276 76188
rect 4300 76186 4356 76188
rect 4380 76186 4436 76188
rect 4460 76186 4516 76188
rect 4220 76134 4266 76186
rect 4266 76134 4276 76186
rect 4300 76134 4330 76186
rect 4330 76134 4342 76186
rect 4342 76134 4356 76186
rect 4380 76134 4394 76186
rect 4394 76134 4406 76186
rect 4406 76134 4436 76186
rect 4460 76134 4470 76186
rect 4470 76134 4516 76186
rect 4220 76132 4276 76134
rect 4300 76132 4356 76134
rect 4380 76132 4436 76134
rect 4460 76132 4516 76134
rect 7484 76186 7540 76188
rect 7564 76186 7620 76188
rect 7644 76186 7700 76188
rect 7724 76186 7780 76188
rect 7484 76134 7530 76186
rect 7530 76134 7540 76186
rect 7564 76134 7594 76186
rect 7594 76134 7606 76186
rect 7606 76134 7620 76186
rect 7644 76134 7658 76186
rect 7658 76134 7670 76186
rect 7670 76134 7700 76186
rect 7724 76134 7734 76186
rect 7734 76134 7780 76186
rect 7484 76132 7540 76134
rect 7564 76132 7620 76134
rect 7644 76132 7700 76134
rect 7724 76132 7780 76134
rect 4220 75098 4276 75100
rect 4300 75098 4356 75100
rect 4380 75098 4436 75100
rect 4460 75098 4516 75100
rect 4220 75046 4266 75098
rect 4266 75046 4276 75098
rect 4300 75046 4330 75098
rect 4330 75046 4342 75098
rect 4342 75046 4356 75098
rect 4380 75046 4394 75098
rect 4394 75046 4406 75098
rect 4406 75046 4436 75098
rect 4460 75046 4470 75098
rect 4470 75046 4516 75098
rect 4220 75044 4276 75046
rect 4300 75044 4356 75046
rect 4380 75044 4436 75046
rect 4460 75044 4516 75046
rect 4220 74010 4276 74012
rect 4300 74010 4356 74012
rect 4380 74010 4436 74012
rect 4460 74010 4516 74012
rect 4220 73958 4266 74010
rect 4266 73958 4276 74010
rect 4300 73958 4330 74010
rect 4330 73958 4342 74010
rect 4342 73958 4356 74010
rect 4380 73958 4394 74010
rect 4394 73958 4406 74010
rect 4406 73958 4436 74010
rect 4460 73958 4470 74010
rect 4470 73958 4516 74010
rect 4220 73956 4276 73958
rect 4300 73956 4356 73958
rect 4380 73956 4436 73958
rect 4460 73956 4516 73958
rect 4220 72922 4276 72924
rect 4300 72922 4356 72924
rect 4380 72922 4436 72924
rect 4460 72922 4516 72924
rect 4220 72870 4266 72922
rect 4266 72870 4276 72922
rect 4300 72870 4330 72922
rect 4330 72870 4342 72922
rect 4342 72870 4356 72922
rect 4380 72870 4394 72922
rect 4394 72870 4406 72922
rect 4406 72870 4436 72922
rect 4460 72870 4470 72922
rect 4470 72870 4516 72922
rect 4220 72868 4276 72870
rect 4300 72868 4356 72870
rect 4380 72868 4436 72870
rect 4460 72868 4516 72870
rect 3422 60968 3478 61024
rect 3514 58404 3570 58440
rect 3514 58384 3516 58404
rect 3516 58384 3568 58404
rect 3568 58384 3570 58404
rect 3698 61784 3754 61840
rect 3698 61668 3754 61704
rect 3698 61648 3700 61668
rect 3700 61648 3752 61668
rect 3752 61648 3754 61668
rect 3790 61376 3846 61432
rect 3514 55800 3570 55856
rect 3514 54984 3570 55040
rect 3606 51312 3662 51368
rect 3514 49544 3570 49600
rect 3330 48728 3386 48784
rect 3330 48048 3386 48104
rect 3514 47796 3570 47832
rect 3514 47776 3516 47796
rect 3516 47776 3568 47796
rect 3568 47776 3570 47796
rect 3330 47232 3386 47288
rect 3054 43424 3110 43480
rect 2588 43002 2644 43004
rect 2668 43002 2724 43004
rect 2748 43002 2804 43004
rect 2828 43002 2884 43004
rect 2588 42950 2634 43002
rect 2634 42950 2644 43002
rect 2668 42950 2698 43002
rect 2698 42950 2710 43002
rect 2710 42950 2724 43002
rect 2748 42950 2762 43002
rect 2762 42950 2774 43002
rect 2774 42950 2804 43002
rect 2828 42950 2838 43002
rect 2838 42950 2884 43002
rect 2588 42948 2644 42950
rect 2668 42948 2724 42950
rect 2748 42948 2804 42950
rect 2828 42948 2884 42950
rect 2778 42744 2834 42800
rect 3146 43152 3202 43208
rect 2588 41914 2644 41916
rect 2668 41914 2724 41916
rect 2748 41914 2804 41916
rect 2828 41914 2884 41916
rect 2588 41862 2634 41914
rect 2634 41862 2644 41914
rect 2668 41862 2698 41914
rect 2698 41862 2710 41914
rect 2710 41862 2724 41914
rect 2748 41862 2762 41914
rect 2762 41862 2774 41914
rect 2774 41862 2804 41914
rect 2828 41862 2838 41914
rect 2838 41862 2884 41914
rect 2588 41860 2644 41862
rect 2668 41860 2724 41862
rect 2748 41860 2804 41862
rect 2828 41860 2884 41862
rect 2962 41112 3018 41168
rect 2870 40976 2926 41032
rect 2588 40826 2644 40828
rect 2668 40826 2724 40828
rect 2748 40826 2804 40828
rect 2828 40826 2884 40828
rect 2588 40774 2634 40826
rect 2634 40774 2644 40826
rect 2668 40774 2698 40826
rect 2698 40774 2710 40826
rect 2710 40774 2724 40826
rect 2748 40774 2762 40826
rect 2762 40774 2774 40826
rect 2774 40774 2804 40826
rect 2828 40774 2838 40826
rect 2838 40774 2884 40826
rect 2588 40772 2644 40774
rect 2668 40772 2724 40774
rect 2748 40772 2804 40774
rect 2828 40772 2884 40774
rect 2594 40432 2650 40488
rect 2588 39738 2644 39740
rect 2668 39738 2724 39740
rect 2748 39738 2804 39740
rect 2828 39738 2884 39740
rect 2588 39686 2634 39738
rect 2634 39686 2644 39738
rect 2668 39686 2698 39738
rect 2698 39686 2710 39738
rect 2710 39686 2724 39738
rect 2748 39686 2762 39738
rect 2762 39686 2774 39738
rect 2774 39686 2804 39738
rect 2828 39686 2838 39738
rect 2838 39686 2884 39738
rect 2588 39684 2644 39686
rect 2668 39684 2724 39686
rect 2748 39684 2804 39686
rect 2828 39684 2884 39686
rect 3422 43596 3424 43616
rect 3424 43596 3476 43616
rect 3476 43596 3478 43616
rect 3422 43560 3478 43596
rect 3790 49952 3846 50008
rect 4220 71834 4276 71836
rect 4300 71834 4356 71836
rect 4380 71834 4436 71836
rect 4460 71834 4516 71836
rect 4220 71782 4266 71834
rect 4266 71782 4276 71834
rect 4300 71782 4330 71834
rect 4330 71782 4342 71834
rect 4342 71782 4356 71834
rect 4380 71782 4394 71834
rect 4394 71782 4406 71834
rect 4406 71782 4436 71834
rect 4460 71782 4470 71834
rect 4470 71782 4516 71834
rect 4220 71780 4276 71782
rect 4300 71780 4356 71782
rect 4380 71780 4436 71782
rect 4460 71780 4516 71782
rect 4220 70746 4276 70748
rect 4300 70746 4356 70748
rect 4380 70746 4436 70748
rect 4460 70746 4516 70748
rect 4220 70694 4266 70746
rect 4266 70694 4276 70746
rect 4300 70694 4330 70746
rect 4330 70694 4342 70746
rect 4342 70694 4356 70746
rect 4380 70694 4394 70746
rect 4394 70694 4406 70746
rect 4406 70694 4436 70746
rect 4460 70694 4470 70746
rect 4470 70694 4516 70746
rect 4220 70692 4276 70694
rect 4300 70692 4356 70694
rect 4380 70692 4436 70694
rect 4460 70692 4516 70694
rect 4220 69658 4276 69660
rect 4300 69658 4356 69660
rect 4380 69658 4436 69660
rect 4460 69658 4516 69660
rect 4220 69606 4266 69658
rect 4266 69606 4276 69658
rect 4300 69606 4330 69658
rect 4330 69606 4342 69658
rect 4342 69606 4356 69658
rect 4380 69606 4394 69658
rect 4394 69606 4406 69658
rect 4406 69606 4436 69658
rect 4460 69606 4470 69658
rect 4470 69606 4516 69658
rect 4220 69604 4276 69606
rect 4300 69604 4356 69606
rect 4380 69604 4436 69606
rect 4460 69604 4516 69606
rect 3974 65048 4030 65104
rect 4220 68570 4276 68572
rect 4300 68570 4356 68572
rect 4380 68570 4436 68572
rect 4460 68570 4516 68572
rect 4220 68518 4266 68570
rect 4266 68518 4276 68570
rect 4300 68518 4330 68570
rect 4330 68518 4342 68570
rect 4342 68518 4356 68570
rect 4380 68518 4394 68570
rect 4394 68518 4406 68570
rect 4406 68518 4436 68570
rect 4460 68518 4470 68570
rect 4470 68518 4516 68570
rect 4220 68516 4276 68518
rect 4300 68516 4356 68518
rect 4380 68516 4436 68518
rect 4460 68516 4516 68518
rect 4220 67482 4276 67484
rect 4300 67482 4356 67484
rect 4380 67482 4436 67484
rect 4460 67482 4516 67484
rect 4220 67430 4266 67482
rect 4266 67430 4276 67482
rect 4300 67430 4330 67482
rect 4330 67430 4342 67482
rect 4342 67430 4356 67482
rect 4380 67430 4394 67482
rect 4394 67430 4406 67482
rect 4406 67430 4436 67482
rect 4460 67430 4470 67482
rect 4470 67430 4516 67482
rect 4220 67428 4276 67430
rect 4300 67428 4356 67430
rect 4380 67428 4436 67430
rect 4460 67428 4516 67430
rect 4220 66394 4276 66396
rect 4300 66394 4356 66396
rect 4380 66394 4436 66396
rect 4460 66394 4516 66396
rect 4220 66342 4266 66394
rect 4266 66342 4276 66394
rect 4300 66342 4330 66394
rect 4330 66342 4342 66394
rect 4342 66342 4356 66394
rect 4380 66342 4394 66394
rect 4394 66342 4406 66394
rect 4406 66342 4436 66394
rect 4460 66342 4470 66394
rect 4470 66342 4516 66394
rect 4220 66340 4276 66342
rect 4300 66340 4356 66342
rect 4380 66340 4436 66342
rect 4460 66340 4516 66342
rect 4220 65306 4276 65308
rect 4300 65306 4356 65308
rect 4380 65306 4436 65308
rect 4460 65306 4516 65308
rect 4220 65254 4266 65306
rect 4266 65254 4276 65306
rect 4300 65254 4330 65306
rect 4330 65254 4342 65306
rect 4342 65254 4356 65306
rect 4380 65254 4394 65306
rect 4394 65254 4406 65306
rect 4406 65254 4436 65306
rect 4460 65254 4470 65306
rect 4470 65254 4516 65306
rect 4220 65252 4276 65254
rect 4300 65252 4356 65254
rect 4380 65252 4436 65254
rect 4460 65252 4516 65254
rect 3974 61376 4030 61432
rect 4220 64218 4276 64220
rect 4300 64218 4356 64220
rect 4380 64218 4436 64220
rect 4460 64218 4516 64220
rect 4220 64166 4266 64218
rect 4266 64166 4276 64218
rect 4300 64166 4330 64218
rect 4330 64166 4342 64218
rect 4342 64166 4356 64218
rect 4380 64166 4394 64218
rect 4394 64166 4406 64218
rect 4406 64166 4436 64218
rect 4460 64166 4470 64218
rect 4470 64166 4516 64218
rect 4220 64164 4276 64166
rect 4300 64164 4356 64166
rect 4380 64164 4436 64166
rect 4460 64164 4516 64166
rect 4220 63130 4276 63132
rect 4300 63130 4356 63132
rect 4380 63130 4436 63132
rect 4460 63130 4516 63132
rect 4220 63078 4266 63130
rect 4266 63078 4276 63130
rect 4300 63078 4330 63130
rect 4330 63078 4342 63130
rect 4342 63078 4356 63130
rect 4380 63078 4394 63130
rect 4394 63078 4406 63130
rect 4406 63078 4436 63130
rect 4460 63078 4470 63130
rect 4470 63078 4516 63130
rect 4220 63076 4276 63078
rect 4300 63076 4356 63078
rect 4380 63076 4436 63078
rect 4460 63076 4516 63078
rect 4220 62042 4276 62044
rect 4300 62042 4356 62044
rect 4380 62042 4436 62044
rect 4460 62042 4516 62044
rect 4220 61990 4266 62042
rect 4266 61990 4276 62042
rect 4300 61990 4330 62042
rect 4330 61990 4342 62042
rect 4342 61990 4356 62042
rect 4380 61990 4394 62042
rect 4394 61990 4406 62042
rect 4406 61990 4436 62042
rect 4460 61990 4470 62042
rect 4470 61990 4516 62042
rect 4220 61988 4276 61990
rect 4300 61988 4356 61990
rect 4380 61988 4436 61990
rect 4460 61988 4516 61990
rect 4220 60954 4276 60956
rect 4300 60954 4356 60956
rect 4380 60954 4436 60956
rect 4460 60954 4516 60956
rect 4220 60902 4266 60954
rect 4266 60902 4276 60954
rect 4300 60902 4330 60954
rect 4330 60902 4342 60954
rect 4342 60902 4356 60954
rect 4380 60902 4394 60954
rect 4394 60902 4406 60954
rect 4406 60902 4436 60954
rect 4460 60902 4470 60954
rect 4470 60902 4516 60954
rect 4220 60900 4276 60902
rect 4300 60900 4356 60902
rect 4380 60900 4436 60902
rect 4460 60900 4516 60902
rect 4066 60560 4122 60616
rect 4066 60424 4122 60480
rect 3974 58656 4030 58712
rect 4220 59866 4276 59868
rect 4300 59866 4356 59868
rect 4380 59866 4436 59868
rect 4460 59866 4516 59868
rect 4220 59814 4266 59866
rect 4266 59814 4276 59866
rect 4300 59814 4330 59866
rect 4330 59814 4342 59866
rect 4342 59814 4356 59866
rect 4380 59814 4394 59866
rect 4394 59814 4406 59866
rect 4406 59814 4436 59866
rect 4460 59814 4470 59866
rect 4470 59814 4516 59866
rect 4220 59812 4276 59814
rect 4300 59812 4356 59814
rect 4380 59812 4436 59814
rect 4460 59812 4516 59814
rect 4220 58778 4276 58780
rect 4300 58778 4356 58780
rect 4380 58778 4436 58780
rect 4460 58778 4516 58780
rect 4220 58726 4266 58778
rect 4266 58726 4276 58778
rect 4300 58726 4330 58778
rect 4330 58726 4342 58778
rect 4342 58726 4356 58778
rect 4380 58726 4394 58778
rect 4394 58726 4406 58778
rect 4406 58726 4436 58778
rect 4460 58726 4470 58778
rect 4470 58726 4516 58778
rect 4220 58724 4276 58726
rect 4300 58724 4356 58726
rect 4380 58724 4436 58726
rect 4460 58724 4516 58726
rect 4220 57690 4276 57692
rect 4300 57690 4356 57692
rect 4380 57690 4436 57692
rect 4460 57690 4516 57692
rect 4220 57638 4266 57690
rect 4266 57638 4276 57690
rect 4300 57638 4330 57690
rect 4330 57638 4342 57690
rect 4342 57638 4356 57690
rect 4380 57638 4394 57690
rect 4394 57638 4406 57690
rect 4406 57638 4436 57690
rect 4460 57638 4470 57690
rect 4470 57638 4516 57690
rect 4220 57636 4276 57638
rect 4300 57636 4356 57638
rect 4380 57636 4436 57638
rect 4460 57636 4516 57638
rect 4220 56602 4276 56604
rect 4300 56602 4356 56604
rect 4380 56602 4436 56604
rect 4460 56602 4516 56604
rect 4220 56550 4266 56602
rect 4266 56550 4276 56602
rect 4300 56550 4330 56602
rect 4330 56550 4342 56602
rect 4342 56550 4356 56602
rect 4380 56550 4394 56602
rect 4394 56550 4406 56602
rect 4406 56550 4436 56602
rect 4460 56550 4470 56602
rect 4470 56550 4516 56602
rect 4220 56548 4276 56550
rect 4300 56548 4356 56550
rect 4380 56548 4436 56550
rect 4460 56548 4516 56550
rect 4158 55700 4160 55720
rect 4160 55700 4212 55720
rect 4212 55700 4214 55720
rect 4158 55664 4214 55700
rect 4220 55514 4276 55516
rect 4300 55514 4356 55516
rect 4380 55514 4436 55516
rect 4460 55514 4516 55516
rect 4220 55462 4266 55514
rect 4266 55462 4276 55514
rect 4300 55462 4330 55514
rect 4330 55462 4342 55514
rect 4342 55462 4356 55514
rect 4380 55462 4394 55514
rect 4394 55462 4406 55514
rect 4406 55462 4436 55514
rect 4460 55462 4470 55514
rect 4470 55462 4516 55514
rect 4220 55460 4276 55462
rect 4300 55460 4356 55462
rect 4380 55460 4436 55462
rect 4460 55460 4516 55462
rect 4342 55156 4344 55176
rect 4344 55156 4396 55176
rect 4396 55156 4398 55176
rect 4342 55120 4398 55156
rect 4220 54426 4276 54428
rect 4300 54426 4356 54428
rect 4380 54426 4436 54428
rect 4460 54426 4516 54428
rect 4220 54374 4266 54426
rect 4266 54374 4276 54426
rect 4300 54374 4330 54426
rect 4330 54374 4342 54426
rect 4342 54374 4356 54426
rect 4380 54374 4394 54426
rect 4394 54374 4406 54426
rect 4406 54374 4436 54426
rect 4460 54374 4470 54426
rect 4470 54374 4516 54426
rect 4220 54372 4276 54374
rect 4300 54372 4356 54374
rect 4380 54372 4436 54374
rect 4460 54372 4516 54374
rect 4220 53338 4276 53340
rect 4300 53338 4356 53340
rect 4380 53338 4436 53340
rect 4460 53338 4516 53340
rect 4220 53286 4266 53338
rect 4266 53286 4276 53338
rect 4300 53286 4330 53338
rect 4330 53286 4342 53338
rect 4342 53286 4356 53338
rect 4380 53286 4394 53338
rect 4394 53286 4406 53338
rect 4406 53286 4436 53338
rect 4460 53286 4470 53338
rect 4470 53286 4516 53338
rect 4220 53284 4276 53286
rect 4300 53284 4356 53286
rect 4380 53284 4436 53286
rect 4460 53284 4516 53286
rect 4158 52692 4214 52728
rect 4158 52672 4160 52692
rect 4160 52672 4212 52692
rect 4212 52672 4214 52692
rect 4220 52250 4276 52252
rect 4300 52250 4356 52252
rect 4380 52250 4436 52252
rect 4460 52250 4516 52252
rect 4220 52198 4266 52250
rect 4266 52198 4276 52250
rect 4300 52198 4330 52250
rect 4330 52198 4342 52250
rect 4342 52198 4356 52250
rect 4380 52198 4394 52250
rect 4394 52198 4406 52250
rect 4406 52198 4436 52250
rect 4460 52198 4470 52250
rect 4470 52198 4516 52250
rect 4220 52196 4276 52198
rect 4300 52196 4356 52198
rect 4380 52196 4436 52198
rect 4460 52196 4516 52198
rect 4618 51448 4674 51504
rect 4220 51162 4276 51164
rect 4300 51162 4356 51164
rect 4380 51162 4436 51164
rect 4460 51162 4516 51164
rect 4220 51110 4266 51162
rect 4266 51110 4276 51162
rect 4300 51110 4330 51162
rect 4330 51110 4342 51162
rect 4342 51110 4356 51162
rect 4380 51110 4394 51162
rect 4394 51110 4406 51162
rect 4406 51110 4436 51162
rect 4460 51110 4470 51162
rect 4470 51110 4516 51162
rect 4802 52808 4858 52864
rect 4220 51108 4276 51110
rect 4300 51108 4356 51110
rect 4380 51108 4436 51110
rect 4460 51108 4516 51110
rect 4066 50904 4122 50960
rect 3790 48184 3846 48240
rect 3422 41656 3478 41712
rect 3514 41520 3570 41576
rect 3698 47096 3754 47152
rect 3698 46572 3754 46608
rect 3698 46552 3700 46572
rect 3700 46552 3752 46572
rect 3752 46552 3754 46572
rect 3882 47096 3938 47152
rect 3974 46688 4030 46744
rect 3882 46436 3938 46472
rect 3882 46416 3884 46436
rect 3884 46416 3936 46436
rect 3936 46416 3938 46436
rect 3606 41384 3662 41440
rect 3606 41248 3662 41304
rect 3514 41112 3570 41168
rect 3422 40976 3478 41032
rect 3422 40432 3478 40488
rect 3330 39908 3386 39944
rect 3330 39888 3332 39908
rect 3332 39888 3384 39908
rect 3384 39888 3386 39908
rect 2594 38800 2650 38856
rect 2778 38800 2834 38856
rect 2588 38650 2644 38652
rect 2668 38650 2724 38652
rect 2748 38650 2804 38652
rect 2828 38650 2884 38652
rect 2588 38598 2634 38650
rect 2634 38598 2644 38650
rect 2668 38598 2698 38650
rect 2698 38598 2710 38650
rect 2710 38598 2724 38650
rect 2748 38598 2762 38650
rect 2762 38598 2774 38650
rect 2774 38598 2804 38650
rect 2828 38598 2838 38650
rect 2838 38598 2884 38650
rect 2588 38596 2644 38598
rect 2668 38596 2724 38598
rect 2748 38596 2804 38598
rect 2828 38596 2884 38598
rect 3146 38664 3202 38720
rect 3146 38548 3202 38584
rect 3146 38528 3148 38548
rect 3148 38528 3200 38548
rect 3200 38528 3202 38548
rect 1858 37848 1914 37904
rect 1674 29144 1730 29200
rect 1858 30096 1914 30152
rect 2318 38120 2374 38176
rect 2318 36488 2374 36544
rect 2318 35556 2374 35592
rect 2318 35536 2320 35556
rect 2320 35536 2372 35556
rect 2372 35536 2374 35556
rect 2778 38392 2834 38448
rect 2588 37562 2644 37564
rect 2668 37562 2724 37564
rect 2748 37562 2804 37564
rect 2828 37562 2884 37564
rect 2588 37510 2634 37562
rect 2634 37510 2644 37562
rect 2668 37510 2698 37562
rect 2698 37510 2710 37562
rect 2710 37510 2724 37562
rect 2748 37510 2762 37562
rect 2762 37510 2774 37562
rect 2774 37510 2804 37562
rect 2828 37510 2838 37562
rect 2838 37510 2884 37562
rect 2588 37508 2644 37510
rect 2668 37508 2724 37510
rect 2748 37508 2804 37510
rect 2828 37508 2884 37510
rect 2588 36474 2644 36476
rect 2668 36474 2724 36476
rect 2748 36474 2804 36476
rect 2828 36474 2884 36476
rect 2588 36422 2634 36474
rect 2634 36422 2644 36474
rect 2668 36422 2698 36474
rect 2698 36422 2710 36474
rect 2710 36422 2724 36474
rect 2748 36422 2762 36474
rect 2762 36422 2774 36474
rect 2774 36422 2804 36474
rect 2828 36422 2838 36474
rect 2838 36422 2884 36474
rect 2588 36420 2644 36422
rect 2668 36420 2724 36422
rect 2748 36420 2804 36422
rect 2828 36420 2884 36422
rect 3330 38256 3386 38312
rect 3146 37848 3202 37904
rect 2962 36080 3018 36136
rect 2588 35386 2644 35388
rect 2668 35386 2724 35388
rect 2748 35386 2804 35388
rect 2828 35386 2884 35388
rect 2588 35334 2634 35386
rect 2634 35334 2644 35386
rect 2668 35334 2698 35386
rect 2698 35334 2710 35386
rect 2710 35334 2724 35386
rect 2748 35334 2762 35386
rect 2762 35334 2774 35386
rect 2774 35334 2804 35386
rect 2828 35334 2838 35386
rect 2838 35334 2884 35386
rect 2588 35332 2644 35334
rect 2668 35332 2724 35334
rect 2748 35332 2804 35334
rect 2828 35332 2884 35334
rect 2134 32680 2190 32736
rect 2318 32544 2374 32600
rect 2042 30096 2098 30152
rect 1858 26832 1914 26888
rect 1766 23840 1822 23896
rect 1398 20576 1454 20632
rect 1398 20168 1454 20224
rect 1490 17584 1546 17640
rect 1398 17176 1454 17232
rect 1582 16768 1638 16824
rect 1490 15544 1546 15600
rect 2134 26696 2190 26752
rect 2042 22072 2098 22128
rect 1674 14728 1730 14784
rect 1582 12552 1638 12608
rect 1582 12280 1638 12336
rect 1306 11736 1362 11792
rect 1214 11192 1270 11248
rect 1306 10784 1362 10840
rect 1398 10376 1454 10432
rect 1306 9968 1362 10024
rect 1398 9560 1454 9616
rect 1398 9152 1454 9208
rect 1398 8608 1454 8664
rect 1398 8200 1454 8256
rect 1398 7828 1400 7848
rect 1400 7828 1452 7848
rect 1452 7828 1454 7848
rect 1398 7792 1454 7828
rect 1398 7404 1454 7440
rect 1398 7384 1400 7404
rect 1400 7384 1452 7404
rect 1452 7384 1454 7404
rect 1950 14320 2006 14376
rect 2778 34448 2834 34504
rect 2588 34298 2644 34300
rect 2668 34298 2724 34300
rect 2748 34298 2804 34300
rect 2828 34298 2884 34300
rect 2588 34246 2634 34298
rect 2634 34246 2644 34298
rect 2668 34246 2698 34298
rect 2698 34246 2710 34298
rect 2710 34246 2724 34298
rect 2748 34246 2762 34298
rect 2762 34246 2774 34298
rect 2774 34246 2804 34298
rect 2828 34246 2838 34298
rect 2838 34246 2884 34298
rect 2588 34244 2644 34246
rect 2668 34244 2724 34246
rect 2748 34244 2804 34246
rect 2828 34244 2884 34246
rect 3054 33904 3110 33960
rect 2588 33210 2644 33212
rect 2668 33210 2724 33212
rect 2748 33210 2804 33212
rect 2828 33210 2884 33212
rect 2588 33158 2634 33210
rect 2634 33158 2644 33210
rect 2668 33158 2698 33210
rect 2698 33158 2710 33210
rect 2710 33158 2724 33210
rect 2748 33158 2762 33210
rect 2762 33158 2774 33210
rect 2774 33158 2804 33210
rect 2828 33158 2838 33210
rect 2838 33158 2884 33210
rect 2588 33156 2644 33158
rect 2668 33156 2724 33158
rect 2748 33156 2804 33158
rect 2828 33156 2884 33158
rect 2778 32816 2834 32872
rect 2588 32122 2644 32124
rect 2668 32122 2724 32124
rect 2748 32122 2804 32124
rect 2828 32122 2884 32124
rect 2588 32070 2634 32122
rect 2634 32070 2644 32122
rect 2668 32070 2698 32122
rect 2698 32070 2710 32122
rect 2710 32070 2724 32122
rect 2748 32070 2762 32122
rect 2762 32070 2774 32122
rect 2774 32070 2804 32122
rect 2828 32070 2838 32122
rect 2838 32070 2884 32122
rect 2588 32068 2644 32070
rect 2668 32068 2724 32070
rect 2748 32068 2804 32070
rect 2828 32068 2884 32070
rect 2318 30232 2374 30288
rect 3054 32292 3110 32328
rect 3054 32272 3056 32292
rect 3056 32272 3108 32292
rect 3108 32272 3110 32292
rect 2588 31034 2644 31036
rect 2668 31034 2724 31036
rect 2748 31034 2804 31036
rect 2828 31034 2884 31036
rect 2588 30982 2634 31034
rect 2634 30982 2644 31034
rect 2668 30982 2698 31034
rect 2698 30982 2710 31034
rect 2710 30982 2724 31034
rect 2748 30982 2762 31034
rect 2762 30982 2774 31034
rect 2774 30982 2804 31034
rect 2828 30982 2838 31034
rect 2838 30982 2884 31034
rect 2588 30980 2644 30982
rect 2668 30980 2724 30982
rect 2748 30980 2804 30982
rect 2828 30980 2884 30982
rect 2778 30540 2780 30560
rect 2780 30540 2832 30560
rect 2832 30540 2834 30560
rect 2778 30504 2834 30540
rect 2588 29946 2644 29948
rect 2668 29946 2724 29948
rect 2748 29946 2804 29948
rect 2828 29946 2884 29948
rect 2588 29894 2634 29946
rect 2634 29894 2644 29946
rect 2668 29894 2698 29946
rect 2698 29894 2710 29946
rect 2710 29894 2724 29946
rect 2748 29894 2762 29946
rect 2762 29894 2774 29946
rect 2774 29894 2804 29946
rect 2828 29894 2838 29946
rect 2838 29894 2884 29946
rect 2588 29892 2644 29894
rect 2668 29892 2724 29894
rect 2748 29892 2804 29894
rect 2828 29892 2884 29894
rect 2778 29572 2834 29608
rect 2778 29552 2780 29572
rect 2780 29552 2832 29572
rect 2832 29552 2834 29572
rect 2962 29280 3018 29336
rect 2588 28858 2644 28860
rect 2668 28858 2724 28860
rect 2748 28858 2804 28860
rect 2828 28858 2884 28860
rect 2588 28806 2634 28858
rect 2634 28806 2644 28858
rect 2668 28806 2698 28858
rect 2698 28806 2710 28858
rect 2710 28806 2724 28858
rect 2748 28806 2762 28858
rect 2762 28806 2774 28858
rect 2774 28806 2804 28858
rect 2828 28806 2838 28858
rect 2838 28806 2884 28858
rect 2588 28804 2644 28806
rect 2668 28804 2724 28806
rect 2748 28804 2804 28806
rect 2828 28804 2884 28806
rect 3514 37732 3570 37768
rect 3514 37712 3516 37732
rect 3516 37712 3568 37732
rect 3568 37712 3570 37732
rect 3422 37304 3478 37360
rect 3422 36644 3478 36680
rect 3422 36624 3424 36644
rect 3424 36624 3476 36644
rect 3476 36624 3478 36644
rect 2318 22208 2374 22264
rect 2226 21936 2282 21992
rect 2226 18128 2282 18184
rect 2962 28600 3018 28656
rect 2588 27770 2644 27772
rect 2668 27770 2724 27772
rect 2748 27770 2804 27772
rect 2828 27770 2884 27772
rect 2588 27718 2634 27770
rect 2634 27718 2644 27770
rect 2668 27718 2698 27770
rect 2698 27718 2710 27770
rect 2710 27718 2724 27770
rect 2748 27718 2762 27770
rect 2762 27718 2774 27770
rect 2774 27718 2804 27770
rect 2828 27718 2838 27770
rect 2838 27718 2884 27770
rect 2588 27716 2644 27718
rect 2668 27716 2724 27718
rect 2748 27716 2804 27718
rect 2828 27716 2884 27718
rect 2778 27572 2834 27628
rect 2588 26682 2644 26684
rect 2668 26682 2724 26684
rect 2748 26682 2804 26684
rect 2828 26682 2884 26684
rect 2588 26630 2634 26682
rect 2634 26630 2644 26682
rect 2668 26630 2698 26682
rect 2698 26630 2710 26682
rect 2710 26630 2724 26682
rect 2748 26630 2762 26682
rect 2762 26630 2774 26682
rect 2774 26630 2804 26682
rect 2828 26630 2838 26682
rect 2838 26630 2884 26682
rect 2588 26628 2644 26630
rect 2668 26628 2724 26630
rect 2748 26628 2804 26630
rect 2828 26628 2884 26630
rect 2594 25744 2650 25800
rect 2588 25594 2644 25596
rect 2668 25594 2724 25596
rect 2748 25594 2804 25596
rect 2828 25594 2884 25596
rect 2588 25542 2634 25594
rect 2634 25542 2644 25594
rect 2668 25542 2698 25594
rect 2698 25542 2710 25594
rect 2710 25542 2724 25594
rect 2748 25542 2762 25594
rect 2762 25542 2774 25594
rect 2774 25542 2804 25594
rect 2828 25542 2838 25594
rect 2838 25542 2884 25594
rect 2588 25540 2644 25542
rect 2668 25540 2724 25542
rect 2748 25540 2804 25542
rect 2828 25540 2884 25542
rect 2778 24812 2834 24848
rect 2778 24792 2780 24812
rect 2780 24792 2832 24812
rect 2832 24792 2834 24812
rect 2588 24506 2644 24508
rect 2668 24506 2724 24508
rect 2748 24506 2804 24508
rect 2828 24506 2884 24508
rect 2588 24454 2634 24506
rect 2634 24454 2644 24506
rect 2668 24454 2698 24506
rect 2698 24454 2710 24506
rect 2710 24454 2724 24506
rect 2748 24454 2762 24506
rect 2762 24454 2774 24506
rect 2774 24454 2804 24506
rect 2828 24454 2838 24506
rect 2838 24454 2884 24506
rect 2588 24452 2644 24454
rect 2668 24452 2724 24454
rect 2748 24452 2804 24454
rect 2828 24452 2884 24454
rect 2962 24112 3018 24168
rect 2778 23604 2780 23624
rect 2780 23604 2832 23624
rect 2832 23604 2834 23624
rect 2778 23568 2834 23604
rect 2588 23418 2644 23420
rect 2668 23418 2724 23420
rect 2748 23418 2804 23420
rect 2828 23418 2884 23420
rect 2588 23366 2634 23418
rect 2634 23366 2644 23418
rect 2668 23366 2698 23418
rect 2698 23366 2710 23418
rect 2710 23366 2724 23418
rect 2748 23366 2762 23418
rect 2762 23366 2774 23418
rect 2774 23366 2804 23418
rect 2828 23366 2838 23418
rect 2838 23366 2884 23418
rect 2588 23364 2644 23366
rect 2668 23364 2724 23366
rect 2748 23364 2804 23366
rect 2828 23364 2884 23366
rect 2588 22330 2644 22332
rect 2668 22330 2724 22332
rect 2748 22330 2804 22332
rect 2828 22330 2884 22332
rect 2588 22278 2634 22330
rect 2634 22278 2644 22330
rect 2668 22278 2698 22330
rect 2698 22278 2710 22330
rect 2710 22278 2724 22330
rect 2748 22278 2762 22330
rect 2762 22278 2774 22330
rect 2774 22278 2804 22330
rect 2828 22278 2838 22330
rect 2838 22278 2884 22330
rect 2588 22276 2644 22278
rect 2668 22276 2724 22278
rect 2748 22276 2804 22278
rect 2828 22276 2884 22278
rect 2502 22072 2558 22128
rect 3054 22772 3110 22808
rect 3054 22752 3056 22772
rect 3056 22752 3108 22772
rect 3108 22752 3110 22772
rect 2588 21242 2644 21244
rect 2668 21242 2724 21244
rect 2748 21242 2804 21244
rect 2828 21242 2884 21244
rect 2588 21190 2634 21242
rect 2634 21190 2644 21242
rect 2668 21190 2698 21242
rect 2698 21190 2710 21242
rect 2710 21190 2724 21242
rect 2748 21190 2762 21242
rect 2762 21190 2774 21242
rect 2774 21190 2804 21242
rect 2828 21190 2838 21242
rect 2838 21190 2884 21242
rect 2588 21188 2644 21190
rect 2668 21188 2724 21190
rect 2748 21188 2804 21190
rect 2828 21188 2884 21190
rect 2588 20154 2644 20156
rect 2668 20154 2724 20156
rect 2748 20154 2804 20156
rect 2828 20154 2884 20156
rect 2588 20102 2634 20154
rect 2634 20102 2644 20154
rect 2668 20102 2698 20154
rect 2698 20102 2710 20154
rect 2710 20102 2724 20154
rect 2748 20102 2762 20154
rect 2762 20102 2774 20154
rect 2774 20102 2804 20154
rect 2828 20102 2838 20154
rect 2838 20102 2884 20154
rect 2588 20100 2644 20102
rect 2668 20100 2724 20102
rect 2748 20100 2804 20102
rect 2828 20100 2884 20102
rect 2870 19352 2926 19408
rect 2778 19216 2834 19272
rect 2588 19066 2644 19068
rect 2668 19066 2724 19068
rect 2748 19066 2804 19068
rect 2828 19066 2884 19068
rect 2588 19014 2634 19066
rect 2634 19014 2644 19066
rect 2668 19014 2698 19066
rect 2698 19014 2710 19066
rect 2710 19014 2724 19066
rect 2748 19014 2762 19066
rect 2762 19014 2774 19066
rect 2774 19014 2804 19066
rect 2828 19014 2838 19066
rect 2838 19014 2884 19066
rect 2588 19012 2644 19014
rect 2668 19012 2724 19014
rect 2748 19012 2804 19014
rect 2828 19012 2884 19014
rect 2870 18536 2926 18592
rect 2588 17978 2644 17980
rect 2668 17978 2724 17980
rect 2748 17978 2804 17980
rect 2828 17978 2884 17980
rect 2588 17926 2634 17978
rect 2634 17926 2644 17978
rect 2668 17926 2698 17978
rect 2698 17926 2710 17978
rect 2710 17926 2724 17978
rect 2748 17926 2762 17978
rect 2762 17926 2774 17978
rect 2774 17926 2804 17978
rect 2828 17926 2838 17978
rect 2838 17926 2884 17978
rect 2588 17924 2644 17926
rect 2668 17924 2724 17926
rect 2748 17924 2804 17926
rect 2828 17924 2884 17926
rect 2588 16890 2644 16892
rect 2668 16890 2724 16892
rect 2748 16890 2804 16892
rect 2828 16890 2884 16892
rect 2588 16838 2634 16890
rect 2634 16838 2644 16890
rect 2668 16838 2698 16890
rect 2698 16838 2710 16890
rect 2710 16838 2724 16890
rect 2748 16838 2762 16890
rect 2762 16838 2774 16890
rect 2774 16838 2804 16890
rect 2828 16838 2838 16890
rect 2838 16838 2884 16890
rect 2588 16836 2644 16838
rect 2668 16836 2724 16838
rect 2748 16836 2804 16838
rect 2828 16836 2884 16838
rect 2778 15952 2834 16008
rect 2588 15802 2644 15804
rect 2668 15802 2724 15804
rect 2748 15802 2804 15804
rect 2828 15802 2884 15804
rect 2588 15750 2634 15802
rect 2634 15750 2644 15802
rect 2668 15750 2698 15802
rect 2698 15750 2710 15802
rect 2710 15750 2724 15802
rect 2748 15750 2762 15802
rect 2762 15750 2774 15802
rect 2774 15750 2804 15802
rect 2828 15750 2838 15802
rect 2838 15750 2884 15802
rect 2588 15748 2644 15750
rect 2668 15748 2724 15750
rect 2748 15748 2804 15750
rect 2828 15748 2884 15750
rect 2042 13096 2098 13152
rect 1582 6704 1638 6760
rect 1306 5616 1362 5672
rect 1398 5208 1454 5264
rect 1398 4020 1400 4040
rect 1400 4020 1452 4040
rect 1452 4020 1454 4040
rect 1398 3984 1454 4020
rect 2870 14864 2926 14920
rect 2588 14714 2644 14716
rect 2668 14714 2724 14716
rect 2748 14714 2804 14716
rect 2828 14714 2884 14716
rect 2588 14662 2634 14714
rect 2634 14662 2644 14714
rect 2668 14662 2698 14714
rect 2698 14662 2710 14714
rect 2710 14662 2724 14714
rect 2748 14662 2762 14714
rect 2762 14662 2774 14714
rect 2774 14662 2804 14714
rect 2828 14662 2838 14714
rect 2838 14662 2884 14714
rect 2588 14660 2644 14662
rect 2668 14660 2724 14662
rect 2748 14660 2804 14662
rect 2828 14660 2884 14662
rect 3146 15036 3148 15056
rect 3148 15036 3200 15056
rect 3200 15036 3202 15056
rect 3146 15000 3202 15036
rect 2588 13626 2644 13628
rect 2668 13626 2724 13628
rect 2748 13626 2804 13628
rect 2828 13626 2884 13628
rect 2588 13574 2634 13626
rect 2634 13574 2644 13626
rect 2668 13574 2698 13626
rect 2698 13574 2710 13626
rect 2710 13574 2724 13626
rect 2748 13574 2762 13626
rect 2762 13574 2774 13626
rect 2774 13574 2804 13626
rect 2828 13574 2838 13626
rect 2838 13574 2884 13626
rect 2588 13572 2644 13574
rect 2668 13572 2724 13574
rect 2748 13572 2804 13574
rect 2828 13572 2884 13574
rect 1858 6160 1914 6216
rect 2226 6976 2282 7032
rect 2226 6568 2282 6624
rect 2588 12538 2644 12540
rect 2668 12538 2724 12540
rect 2748 12538 2804 12540
rect 2828 12538 2884 12540
rect 2588 12486 2634 12538
rect 2634 12486 2644 12538
rect 2668 12486 2698 12538
rect 2698 12486 2710 12538
rect 2710 12486 2724 12538
rect 2748 12486 2762 12538
rect 2762 12486 2774 12538
rect 2774 12486 2804 12538
rect 2828 12486 2838 12538
rect 2838 12486 2884 12538
rect 2588 12484 2644 12486
rect 2668 12484 2724 12486
rect 2748 12484 2804 12486
rect 2828 12484 2884 12486
rect 2588 11450 2644 11452
rect 2668 11450 2724 11452
rect 2748 11450 2804 11452
rect 2828 11450 2884 11452
rect 2588 11398 2634 11450
rect 2634 11398 2644 11450
rect 2668 11398 2698 11450
rect 2698 11398 2710 11450
rect 2710 11398 2724 11450
rect 2748 11398 2762 11450
rect 2762 11398 2774 11450
rect 2774 11398 2804 11450
rect 2828 11398 2838 11450
rect 2838 11398 2884 11450
rect 2588 11396 2644 11398
rect 2668 11396 2724 11398
rect 2748 11396 2804 11398
rect 2828 11396 2884 11398
rect 2588 10362 2644 10364
rect 2668 10362 2724 10364
rect 2748 10362 2804 10364
rect 2828 10362 2884 10364
rect 2588 10310 2634 10362
rect 2634 10310 2644 10362
rect 2668 10310 2698 10362
rect 2698 10310 2710 10362
rect 2710 10310 2724 10362
rect 2748 10310 2762 10362
rect 2762 10310 2774 10362
rect 2774 10310 2804 10362
rect 2828 10310 2838 10362
rect 2838 10310 2884 10362
rect 2588 10308 2644 10310
rect 2668 10308 2724 10310
rect 2748 10308 2804 10310
rect 2828 10308 2884 10310
rect 3422 36488 3478 36544
rect 3422 32000 3478 32056
rect 3330 30776 3386 30832
rect 3330 28328 3386 28384
rect 3790 45600 3846 45656
rect 3974 45464 4030 45520
rect 3882 43832 3938 43888
rect 3790 43288 3846 43344
rect 3790 42880 3846 42936
rect 3790 42744 3846 42800
rect 3790 42084 3846 42120
rect 3790 42064 3792 42084
rect 3792 42064 3844 42084
rect 3844 42064 3846 42084
rect 3790 41928 3846 41984
rect 3790 41384 3846 41440
rect 3974 43152 4030 43208
rect 3974 42472 4030 42528
rect 3882 41248 3938 41304
rect 4618 50768 4674 50824
rect 4220 50074 4276 50076
rect 4300 50074 4356 50076
rect 4380 50074 4436 50076
rect 4460 50074 4516 50076
rect 4220 50022 4266 50074
rect 4266 50022 4276 50074
rect 4300 50022 4330 50074
rect 4330 50022 4342 50074
rect 4342 50022 4356 50074
rect 4380 50022 4394 50074
rect 4394 50022 4406 50074
rect 4406 50022 4436 50074
rect 4460 50022 4470 50074
rect 4470 50022 4516 50074
rect 4220 50020 4276 50022
rect 4300 50020 4356 50022
rect 4380 50020 4436 50022
rect 4460 50020 4516 50022
rect 4526 49308 4528 49328
rect 4528 49308 4580 49328
rect 4580 49308 4582 49328
rect 4526 49272 4582 49308
rect 4220 48986 4276 48988
rect 4300 48986 4356 48988
rect 4380 48986 4436 48988
rect 4460 48986 4516 48988
rect 4220 48934 4266 48986
rect 4266 48934 4276 48986
rect 4300 48934 4330 48986
rect 4330 48934 4342 48986
rect 4342 48934 4356 48986
rect 4380 48934 4394 48986
rect 4394 48934 4406 48986
rect 4406 48934 4436 48986
rect 4460 48934 4470 48986
rect 4470 48934 4516 48986
rect 4220 48932 4276 48934
rect 4300 48932 4356 48934
rect 4380 48932 4436 48934
rect 4460 48932 4516 48934
rect 4526 48456 4582 48512
rect 4526 48068 4582 48104
rect 4526 48048 4528 48068
rect 4528 48048 4580 48068
rect 4580 48048 4582 48068
rect 4220 47898 4276 47900
rect 4300 47898 4356 47900
rect 4380 47898 4436 47900
rect 4460 47898 4516 47900
rect 4220 47846 4266 47898
rect 4266 47846 4276 47898
rect 4300 47846 4330 47898
rect 4330 47846 4342 47898
rect 4342 47846 4356 47898
rect 4380 47846 4394 47898
rect 4394 47846 4406 47898
rect 4406 47846 4436 47898
rect 4460 47846 4470 47898
rect 4470 47846 4516 47898
rect 4220 47844 4276 47846
rect 4300 47844 4356 47846
rect 4380 47844 4436 47846
rect 4460 47844 4516 47846
rect 4618 47504 4674 47560
rect 4526 46996 4528 47016
rect 4528 46996 4580 47016
rect 4580 46996 4582 47016
rect 4526 46960 4582 46996
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4266 46810
rect 4266 46758 4276 46810
rect 4300 46758 4330 46810
rect 4330 46758 4342 46810
rect 4342 46758 4356 46810
rect 4380 46758 4394 46810
rect 4394 46758 4406 46810
rect 4406 46758 4436 46810
rect 4460 46758 4470 46810
rect 4470 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4802 50632 4858 50688
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4266 45722
rect 4266 45670 4276 45722
rect 4300 45670 4330 45722
rect 4330 45670 4342 45722
rect 4342 45670 4356 45722
rect 4380 45670 4394 45722
rect 4394 45670 4406 45722
rect 4406 45670 4436 45722
rect 4460 45670 4470 45722
rect 4470 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4266 44634
rect 4266 44582 4276 44634
rect 4300 44582 4330 44634
rect 4330 44582 4342 44634
rect 4342 44582 4356 44634
rect 4380 44582 4394 44634
rect 4394 44582 4406 44634
rect 4406 44582 4436 44634
rect 4460 44582 4470 44634
rect 4470 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4266 43546
rect 4266 43494 4276 43546
rect 4300 43494 4330 43546
rect 4330 43494 4342 43546
rect 4342 43494 4356 43546
rect 4380 43494 4394 43546
rect 4394 43494 4406 43546
rect 4406 43494 4436 43546
rect 4460 43494 4470 43546
rect 4470 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4158 43288 4214 43344
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4266 42458
rect 4266 42406 4276 42458
rect 4300 42406 4330 42458
rect 4330 42406 4342 42458
rect 4342 42406 4356 42458
rect 4380 42406 4394 42458
rect 4394 42406 4406 42458
rect 4406 42406 4436 42458
rect 4460 42406 4470 42458
rect 4470 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4266 41370
rect 4266 41318 4276 41370
rect 4300 41318 4330 41370
rect 4330 41318 4342 41370
rect 4342 41318 4356 41370
rect 4380 41318 4394 41370
rect 4394 41318 4406 41370
rect 4406 41318 4436 41370
rect 4460 41318 4470 41370
rect 4470 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 3974 39752 4030 39808
rect 3882 39344 3938 39400
rect 3790 39072 3846 39128
rect 3882 38392 3938 38448
rect 3790 37712 3846 37768
rect 3790 35264 3846 35320
rect 3698 35128 3754 35184
rect 3790 33768 3846 33824
rect 3606 27104 3662 27160
rect 3974 32000 4030 32056
rect 3974 31728 4030 31784
rect 3606 26424 3662 26480
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4266 40282
rect 4266 40230 4276 40282
rect 4300 40230 4330 40282
rect 4330 40230 4342 40282
rect 4342 40230 4356 40282
rect 4380 40230 4394 40282
rect 4394 40230 4406 40282
rect 4406 40230 4436 40282
rect 4460 40230 4470 40282
rect 4470 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4526 40024 4582 40080
rect 4250 39344 4306 39400
rect 4710 39888 4766 39944
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4266 39194
rect 4266 39142 4276 39194
rect 4300 39142 4330 39194
rect 4330 39142 4342 39194
rect 4342 39142 4356 39194
rect 4380 39142 4394 39194
rect 4394 39142 4406 39194
rect 4406 39142 4436 39194
rect 4460 39142 4470 39194
rect 4470 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4342 38936 4398 38992
rect 4342 38256 4398 38312
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4266 38106
rect 4266 38054 4276 38106
rect 4300 38054 4330 38106
rect 4330 38054 4342 38106
rect 4342 38054 4356 38106
rect 4380 38054 4394 38106
rect 4394 38054 4406 38106
rect 4406 38054 4436 38106
rect 4460 38054 4470 38106
rect 4470 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4266 37018
rect 4266 36966 4276 37018
rect 4300 36966 4330 37018
rect 4330 36966 4342 37018
rect 4342 36966 4356 37018
rect 4380 36966 4394 37018
rect 4394 36966 4406 37018
rect 4406 36966 4436 37018
rect 4460 36966 4470 37018
rect 4470 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4526 36796 4528 36816
rect 4528 36796 4580 36816
rect 4580 36796 4582 36816
rect 4526 36760 4582 36796
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4266 35930
rect 4266 35878 4276 35930
rect 4300 35878 4330 35930
rect 4330 35878 4342 35930
rect 4342 35878 4356 35930
rect 4380 35878 4394 35930
rect 4394 35878 4406 35930
rect 4406 35878 4436 35930
rect 4460 35878 4470 35930
rect 4470 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4618 35672 4674 35728
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4266 34842
rect 4266 34790 4276 34842
rect 4300 34790 4330 34842
rect 4330 34790 4342 34842
rect 4342 34790 4356 34842
rect 4380 34790 4394 34842
rect 4394 34790 4406 34842
rect 4406 34790 4436 34842
rect 4460 34790 4470 34842
rect 4470 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4158 33904 4214 33960
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4266 33754
rect 4266 33702 4276 33754
rect 4300 33702 4330 33754
rect 4330 33702 4342 33754
rect 4342 33702 4356 33754
rect 4380 33702 4394 33754
rect 4394 33702 4406 33754
rect 4406 33702 4436 33754
rect 4460 33702 4470 33754
rect 4470 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4266 32666
rect 4266 32614 4276 32666
rect 4300 32614 4330 32666
rect 4330 32614 4342 32666
rect 4342 32614 4356 32666
rect 4380 32614 4394 32666
rect 4394 32614 4406 32666
rect 4406 32614 4436 32666
rect 4460 32614 4470 32666
rect 4470 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4250 32408 4306 32464
rect 5078 58928 5134 58984
rect 4986 50904 5042 50960
rect 5078 50632 5134 50688
rect 4894 42064 4950 42120
rect 4802 35944 4858 36000
rect 4986 41792 5042 41848
rect 5852 75642 5908 75644
rect 5932 75642 5988 75644
rect 6012 75642 6068 75644
rect 6092 75642 6148 75644
rect 5852 75590 5898 75642
rect 5898 75590 5908 75642
rect 5932 75590 5962 75642
rect 5962 75590 5974 75642
rect 5974 75590 5988 75642
rect 6012 75590 6026 75642
rect 6026 75590 6038 75642
rect 6038 75590 6068 75642
rect 6092 75590 6102 75642
rect 6102 75590 6148 75642
rect 5852 75588 5908 75590
rect 5932 75588 5988 75590
rect 6012 75588 6068 75590
rect 6092 75588 6148 75590
rect 7484 75098 7540 75100
rect 7564 75098 7620 75100
rect 7644 75098 7700 75100
rect 7724 75098 7780 75100
rect 7484 75046 7530 75098
rect 7530 75046 7540 75098
rect 7564 75046 7594 75098
rect 7594 75046 7606 75098
rect 7606 75046 7620 75098
rect 7644 75046 7658 75098
rect 7658 75046 7670 75098
rect 7670 75046 7700 75098
rect 7724 75046 7734 75098
rect 7734 75046 7780 75098
rect 7484 75044 7540 75046
rect 7564 75044 7620 75046
rect 7644 75044 7700 75046
rect 7724 75044 7780 75046
rect 5852 74554 5908 74556
rect 5932 74554 5988 74556
rect 6012 74554 6068 74556
rect 6092 74554 6148 74556
rect 5852 74502 5898 74554
rect 5898 74502 5908 74554
rect 5932 74502 5962 74554
rect 5962 74502 5974 74554
rect 5974 74502 5988 74554
rect 6012 74502 6026 74554
rect 6026 74502 6038 74554
rect 6038 74502 6068 74554
rect 6092 74502 6102 74554
rect 6102 74502 6148 74554
rect 5852 74500 5908 74502
rect 5932 74500 5988 74502
rect 6012 74500 6068 74502
rect 6092 74500 6148 74502
rect 7484 74010 7540 74012
rect 7564 74010 7620 74012
rect 7644 74010 7700 74012
rect 7724 74010 7780 74012
rect 7484 73958 7530 74010
rect 7530 73958 7540 74010
rect 7564 73958 7594 74010
rect 7594 73958 7606 74010
rect 7606 73958 7620 74010
rect 7644 73958 7658 74010
rect 7658 73958 7670 74010
rect 7670 73958 7700 74010
rect 7724 73958 7734 74010
rect 7734 73958 7780 74010
rect 7484 73956 7540 73958
rect 7564 73956 7620 73958
rect 7644 73956 7700 73958
rect 7724 73956 7780 73958
rect 5852 73466 5908 73468
rect 5932 73466 5988 73468
rect 6012 73466 6068 73468
rect 6092 73466 6148 73468
rect 5852 73414 5898 73466
rect 5898 73414 5908 73466
rect 5932 73414 5962 73466
rect 5962 73414 5974 73466
rect 5974 73414 5988 73466
rect 6012 73414 6026 73466
rect 6026 73414 6038 73466
rect 6038 73414 6068 73466
rect 6092 73414 6102 73466
rect 6102 73414 6148 73466
rect 5852 73412 5908 73414
rect 5932 73412 5988 73414
rect 6012 73412 6068 73414
rect 6092 73412 6148 73414
rect 7484 72922 7540 72924
rect 7564 72922 7620 72924
rect 7644 72922 7700 72924
rect 7724 72922 7780 72924
rect 7484 72870 7530 72922
rect 7530 72870 7540 72922
rect 7564 72870 7594 72922
rect 7594 72870 7606 72922
rect 7606 72870 7620 72922
rect 7644 72870 7658 72922
rect 7658 72870 7670 72922
rect 7670 72870 7700 72922
rect 7724 72870 7734 72922
rect 7734 72870 7780 72922
rect 7484 72868 7540 72870
rect 7564 72868 7620 72870
rect 7644 72868 7700 72870
rect 7724 72868 7780 72870
rect 5446 66136 5502 66192
rect 5354 52672 5410 52728
rect 5354 52128 5410 52184
rect 5354 51032 5410 51088
rect 5354 50768 5410 50824
rect 5262 41248 5318 41304
rect 4986 40568 5042 40624
rect 4526 31728 4582 31784
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4266 31578
rect 4266 31526 4276 31578
rect 4300 31526 4330 31578
rect 4330 31526 4342 31578
rect 4342 31526 4356 31578
rect 4380 31526 4394 31578
rect 4394 31526 4406 31578
rect 4406 31526 4436 31578
rect 4460 31526 4470 31578
rect 4470 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4526 31320 4582 31376
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4266 30490
rect 4266 30438 4276 30490
rect 4300 30438 4330 30490
rect 4330 30438 4342 30490
rect 4342 30438 4356 30490
rect 4380 30438 4394 30490
rect 4394 30438 4406 30490
rect 4406 30438 4436 30490
rect 4460 30438 4470 30490
rect 4470 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4266 29402
rect 4266 29350 4276 29402
rect 4300 29350 4330 29402
rect 4330 29350 4342 29402
rect 4342 29350 4356 29402
rect 4380 29350 4394 29402
rect 4394 29350 4406 29402
rect 4406 29350 4436 29402
rect 4460 29350 4470 29402
rect 4470 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 3974 28192 4030 28248
rect 3514 26188 3516 26208
rect 3516 26188 3568 26208
rect 3568 26188 3570 26208
rect 3514 26152 3570 26188
rect 3330 24656 3386 24712
rect 3238 12960 3294 13016
rect 3238 12180 3240 12200
rect 3240 12180 3292 12200
rect 3292 12180 3294 12200
rect 3238 12144 3294 12180
rect 3422 24520 3478 24576
rect 3606 25200 3662 25256
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4266 28314
rect 4266 28262 4276 28314
rect 4300 28262 4330 28314
rect 4330 28262 4342 28314
rect 4342 28262 4356 28314
rect 4380 28262 4394 28314
rect 4394 28262 4406 28314
rect 4406 28262 4436 28314
rect 4460 28262 4470 28314
rect 4470 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4250 28056 4306 28112
rect 4250 27512 4306 27568
rect 4434 27376 4490 27432
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4266 27226
rect 4266 27174 4276 27226
rect 4300 27174 4330 27226
rect 4330 27174 4342 27226
rect 4342 27174 4356 27226
rect 4380 27174 4394 27226
rect 4394 27174 4406 27226
rect 4406 27174 4436 27226
rect 4460 27174 4470 27226
rect 4470 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4266 26138
rect 4266 26086 4276 26138
rect 4300 26086 4330 26138
rect 4330 26086 4342 26138
rect 4342 26086 4356 26138
rect 4380 26086 4394 26138
rect 4394 26086 4406 26138
rect 4406 26086 4436 26138
rect 4460 26086 4470 26138
rect 4470 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4526 25880 4582 25936
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4266 25050
rect 4266 24998 4276 25050
rect 4300 24998 4330 25050
rect 4330 24998 4342 25050
rect 4342 24998 4356 25050
rect 4380 24998 4394 25050
rect 4394 24998 4406 25050
rect 4406 24998 4436 25050
rect 4460 24998 4470 25050
rect 4470 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4986 31184 5042 31240
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4266 23962
rect 4266 23910 4276 23962
rect 4300 23910 4330 23962
rect 4330 23910 4342 23962
rect 4342 23910 4356 23962
rect 4380 23910 4394 23962
rect 4394 23910 4406 23962
rect 4406 23910 4436 23962
rect 4460 23910 4470 23962
rect 4470 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 3790 22616 3846 22672
rect 3790 22344 3846 22400
rect 3698 22208 3754 22264
rect 2870 9444 2926 9480
rect 2870 9424 2872 9444
rect 2872 9424 2924 9444
rect 2924 9424 2926 9444
rect 2588 9274 2644 9276
rect 2668 9274 2724 9276
rect 2748 9274 2804 9276
rect 2828 9274 2884 9276
rect 2588 9222 2634 9274
rect 2634 9222 2644 9274
rect 2668 9222 2698 9274
rect 2698 9222 2710 9274
rect 2710 9222 2724 9274
rect 2748 9222 2762 9274
rect 2762 9222 2774 9274
rect 2774 9222 2804 9274
rect 2828 9222 2838 9274
rect 2838 9222 2884 9274
rect 2588 9220 2644 9222
rect 2668 9220 2724 9222
rect 2748 9220 2804 9222
rect 2828 9220 2884 9222
rect 2962 9172 3018 9208
rect 2962 9152 2964 9172
rect 2964 9152 3016 9172
rect 3016 9152 3018 9172
rect 2588 8186 2644 8188
rect 2668 8186 2724 8188
rect 2748 8186 2804 8188
rect 2828 8186 2884 8188
rect 2588 8134 2634 8186
rect 2634 8134 2644 8186
rect 2668 8134 2698 8186
rect 2698 8134 2710 8186
rect 2710 8134 2724 8186
rect 2748 8134 2762 8186
rect 2762 8134 2774 8186
rect 2774 8134 2804 8186
rect 2828 8134 2838 8186
rect 2838 8134 2884 8186
rect 2588 8132 2644 8134
rect 2668 8132 2724 8134
rect 2748 8132 2804 8134
rect 2828 8132 2884 8134
rect 2588 7098 2644 7100
rect 2668 7098 2724 7100
rect 2748 7098 2804 7100
rect 2828 7098 2884 7100
rect 2588 7046 2634 7098
rect 2634 7046 2644 7098
rect 2668 7046 2698 7098
rect 2698 7046 2710 7098
rect 2710 7046 2724 7098
rect 2748 7046 2762 7098
rect 2762 7046 2774 7098
rect 2774 7046 2804 7098
rect 2828 7046 2838 7098
rect 2838 7046 2884 7098
rect 2588 7044 2644 7046
rect 2668 7044 2724 7046
rect 2748 7044 2804 7046
rect 2828 7044 2884 7046
rect 2588 6010 2644 6012
rect 2668 6010 2724 6012
rect 2748 6010 2804 6012
rect 2828 6010 2884 6012
rect 2588 5958 2634 6010
rect 2634 5958 2644 6010
rect 2668 5958 2698 6010
rect 2698 5958 2710 6010
rect 2710 5958 2724 6010
rect 2748 5958 2762 6010
rect 2762 5958 2774 6010
rect 2774 5958 2804 6010
rect 2828 5958 2838 6010
rect 2838 5958 2884 6010
rect 2588 5956 2644 5958
rect 2668 5956 2724 5958
rect 2748 5956 2804 5958
rect 2828 5956 2884 5958
rect 2588 4922 2644 4924
rect 2668 4922 2724 4924
rect 2748 4922 2804 4924
rect 2828 4922 2884 4924
rect 2588 4870 2634 4922
rect 2634 4870 2644 4922
rect 2668 4870 2698 4922
rect 2698 4870 2710 4922
rect 2710 4870 2724 4922
rect 2748 4870 2762 4922
rect 2762 4870 2774 4922
rect 2774 4870 2804 4922
rect 2828 4870 2838 4922
rect 2838 4870 2884 4922
rect 2588 4868 2644 4870
rect 2668 4868 2724 4870
rect 2748 4868 2804 4870
rect 2828 4868 2884 4870
rect 2962 4392 3018 4448
rect 2318 3168 2374 3224
rect 2588 3834 2644 3836
rect 2668 3834 2724 3836
rect 2748 3834 2804 3836
rect 2828 3834 2884 3836
rect 2588 3782 2634 3834
rect 2634 3782 2644 3834
rect 2668 3782 2698 3834
rect 2698 3782 2710 3834
rect 2710 3782 2724 3834
rect 2748 3782 2762 3834
rect 2762 3782 2774 3834
rect 2774 3782 2804 3834
rect 2828 3782 2838 3834
rect 2838 3782 2884 3834
rect 2588 3780 2644 3782
rect 2668 3780 2724 3782
rect 2748 3780 2804 3782
rect 2828 3780 2884 3782
rect 2962 3576 3018 3632
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4266 22874
rect 4266 22822 4276 22874
rect 4300 22822 4330 22874
rect 4330 22822 4342 22874
rect 4342 22822 4356 22874
rect 4380 22822 4394 22874
rect 4394 22822 4406 22874
rect 4406 22822 4436 22874
rect 4460 22822 4470 22874
rect 4470 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4266 21786
rect 4266 21734 4276 21786
rect 4300 21734 4330 21786
rect 4330 21734 4342 21786
rect 4342 21734 4356 21786
rect 4380 21734 4394 21786
rect 4394 21734 4406 21786
rect 4406 21734 4436 21786
rect 4460 21734 4470 21786
rect 4470 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4266 20698
rect 4266 20646 4276 20698
rect 4300 20646 4330 20698
rect 4330 20646 4342 20698
rect 4342 20646 4356 20698
rect 4380 20646 4394 20698
rect 4394 20646 4406 20698
rect 4406 20646 4436 20698
rect 4460 20646 4470 20698
rect 4470 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 3974 19796 3976 19816
rect 3976 19796 4028 19816
rect 4028 19796 4030 19816
rect 3974 19760 4030 19796
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4266 19610
rect 4266 19558 4276 19610
rect 4300 19558 4330 19610
rect 4330 19558 4342 19610
rect 4342 19558 4356 19610
rect 4380 19558 4394 19610
rect 4394 19558 4406 19610
rect 4406 19558 4436 19610
rect 4460 19558 4470 19610
rect 4470 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4266 18522
rect 4266 18470 4276 18522
rect 4300 18470 4330 18522
rect 4330 18470 4342 18522
rect 4342 18470 4356 18522
rect 4380 18470 4394 18522
rect 4394 18470 4406 18522
rect 4406 18470 4436 18522
rect 4460 18470 4470 18522
rect 4470 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4266 17434
rect 4266 17382 4276 17434
rect 4300 17382 4330 17434
rect 4330 17382 4342 17434
rect 4342 17382 4356 17434
rect 4380 17382 4394 17434
rect 4394 17382 4406 17434
rect 4406 17382 4436 17434
rect 4460 17382 4470 17434
rect 4470 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 3974 16360 4030 16416
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4266 16346
rect 4266 16294 4276 16346
rect 4300 16294 4330 16346
rect 4330 16294 4342 16346
rect 4342 16294 4356 16346
rect 4380 16294 4394 16346
rect 4394 16294 4406 16346
rect 4406 16294 4436 16346
rect 4460 16294 4470 16346
rect 4470 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 3974 15136 4030 15192
rect 3974 14184 4030 14240
rect 3974 13776 4030 13832
rect 3882 13368 3938 13424
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4266 15258
rect 4266 15206 4276 15258
rect 4300 15206 4330 15258
rect 4330 15206 4342 15258
rect 4342 15206 4356 15258
rect 4380 15206 4394 15258
rect 4394 15206 4406 15258
rect 4406 15206 4436 15258
rect 4460 15206 4470 15258
rect 4470 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4266 14170
rect 4266 14118 4276 14170
rect 4300 14118 4330 14170
rect 4330 14118 4342 14170
rect 4342 14118 4356 14170
rect 4380 14118 4394 14170
rect 4394 14118 4406 14170
rect 4406 14118 4436 14170
rect 4460 14118 4470 14170
rect 4470 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4266 13082
rect 4266 13030 4276 13082
rect 4300 13030 4330 13082
rect 4330 13030 4342 13082
rect 4342 13030 4356 13082
rect 4380 13030 4394 13082
rect 4394 13030 4406 13082
rect 4406 13030 4436 13082
rect 4460 13030 4470 13082
rect 4470 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 3698 8472 3754 8528
rect 3330 4664 3386 4720
rect 2588 2746 2644 2748
rect 2668 2746 2724 2748
rect 2748 2746 2804 2748
rect 2828 2746 2884 2748
rect 2588 2694 2634 2746
rect 2634 2694 2644 2746
rect 2668 2694 2698 2746
rect 2698 2694 2710 2746
rect 2710 2694 2724 2746
rect 2748 2694 2762 2746
rect 2762 2694 2774 2746
rect 2774 2694 2804 2746
rect 2828 2694 2838 2746
rect 2838 2694 2884 2746
rect 2588 2692 2644 2694
rect 2668 2692 2724 2694
rect 2748 2692 2804 2694
rect 2828 2692 2884 2694
rect 2778 2216 2834 2272
rect 2778 1028 2780 1048
rect 2780 1028 2832 1048
rect 2832 1028 2834 1048
rect 2778 992 2834 1028
rect 3698 5208 3754 5264
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4266 11994
rect 4266 11942 4276 11994
rect 4300 11942 4330 11994
rect 4330 11942 4342 11994
rect 4342 11942 4356 11994
rect 4380 11942 4394 11994
rect 4394 11942 4406 11994
rect 4406 11942 4436 11994
rect 4460 11942 4470 11994
rect 4470 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 3974 9016 4030 9072
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4266 10906
rect 4266 10854 4276 10906
rect 4300 10854 4330 10906
rect 4330 10854 4342 10906
rect 4342 10854 4356 10906
rect 4380 10854 4394 10906
rect 4394 10854 4406 10906
rect 4406 10854 4436 10906
rect 4460 10854 4470 10906
rect 4470 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 5262 40840 5318 40896
rect 5170 32136 5226 32192
rect 5170 27920 5226 27976
rect 5852 72378 5908 72380
rect 5932 72378 5988 72380
rect 6012 72378 6068 72380
rect 6092 72378 6148 72380
rect 5852 72326 5898 72378
rect 5898 72326 5908 72378
rect 5932 72326 5962 72378
rect 5962 72326 5974 72378
rect 5974 72326 5988 72378
rect 6012 72326 6026 72378
rect 6026 72326 6038 72378
rect 6038 72326 6068 72378
rect 6092 72326 6102 72378
rect 6102 72326 6148 72378
rect 5852 72324 5908 72326
rect 5932 72324 5988 72326
rect 6012 72324 6068 72326
rect 6092 72324 6148 72326
rect 7484 71834 7540 71836
rect 7564 71834 7620 71836
rect 7644 71834 7700 71836
rect 7724 71834 7780 71836
rect 7484 71782 7530 71834
rect 7530 71782 7540 71834
rect 7564 71782 7594 71834
rect 7594 71782 7606 71834
rect 7606 71782 7620 71834
rect 7644 71782 7658 71834
rect 7658 71782 7670 71834
rect 7670 71782 7700 71834
rect 7724 71782 7734 71834
rect 7734 71782 7780 71834
rect 7484 71780 7540 71782
rect 7564 71780 7620 71782
rect 7644 71780 7700 71782
rect 7724 71780 7780 71782
rect 5852 71290 5908 71292
rect 5932 71290 5988 71292
rect 6012 71290 6068 71292
rect 6092 71290 6148 71292
rect 5852 71238 5898 71290
rect 5898 71238 5908 71290
rect 5932 71238 5962 71290
rect 5962 71238 5974 71290
rect 5974 71238 5988 71290
rect 6012 71238 6026 71290
rect 6026 71238 6038 71290
rect 6038 71238 6068 71290
rect 6092 71238 6102 71290
rect 6102 71238 6148 71290
rect 5852 71236 5908 71238
rect 5932 71236 5988 71238
rect 6012 71236 6068 71238
rect 6092 71236 6148 71238
rect 7484 70746 7540 70748
rect 7564 70746 7620 70748
rect 7644 70746 7700 70748
rect 7724 70746 7780 70748
rect 7484 70694 7530 70746
rect 7530 70694 7540 70746
rect 7564 70694 7594 70746
rect 7594 70694 7606 70746
rect 7606 70694 7620 70746
rect 7644 70694 7658 70746
rect 7658 70694 7670 70746
rect 7670 70694 7700 70746
rect 7724 70694 7734 70746
rect 7734 70694 7780 70746
rect 7484 70692 7540 70694
rect 7564 70692 7620 70694
rect 7644 70692 7700 70694
rect 7724 70692 7780 70694
rect 5852 70202 5908 70204
rect 5932 70202 5988 70204
rect 6012 70202 6068 70204
rect 6092 70202 6148 70204
rect 5852 70150 5898 70202
rect 5898 70150 5908 70202
rect 5932 70150 5962 70202
rect 5962 70150 5974 70202
rect 5974 70150 5988 70202
rect 6012 70150 6026 70202
rect 6026 70150 6038 70202
rect 6038 70150 6068 70202
rect 6092 70150 6102 70202
rect 6102 70150 6148 70202
rect 5852 70148 5908 70150
rect 5932 70148 5988 70150
rect 6012 70148 6068 70150
rect 6092 70148 6148 70150
rect 7484 69658 7540 69660
rect 7564 69658 7620 69660
rect 7644 69658 7700 69660
rect 7724 69658 7780 69660
rect 7484 69606 7530 69658
rect 7530 69606 7540 69658
rect 7564 69606 7594 69658
rect 7594 69606 7606 69658
rect 7606 69606 7620 69658
rect 7644 69606 7658 69658
rect 7658 69606 7670 69658
rect 7670 69606 7700 69658
rect 7724 69606 7734 69658
rect 7734 69606 7780 69658
rect 7484 69604 7540 69606
rect 7564 69604 7620 69606
rect 7644 69604 7700 69606
rect 7724 69604 7780 69606
rect 5852 69114 5908 69116
rect 5932 69114 5988 69116
rect 6012 69114 6068 69116
rect 6092 69114 6148 69116
rect 5852 69062 5898 69114
rect 5898 69062 5908 69114
rect 5932 69062 5962 69114
rect 5962 69062 5974 69114
rect 5974 69062 5988 69114
rect 6012 69062 6026 69114
rect 6026 69062 6038 69114
rect 6038 69062 6068 69114
rect 6092 69062 6102 69114
rect 6102 69062 6148 69114
rect 5852 69060 5908 69062
rect 5932 69060 5988 69062
rect 6012 69060 6068 69062
rect 6092 69060 6148 69062
rect 7484 68570 7540 68572
rect 7564 68570 7620 68572
rect 7644 68570 7700 68572
rect 7724 68570 7780 68572
rect 7484 68518 7530 68570
rect 7530 68518 7540 68570
rect 7564 68518 7594 68570
rect 7594 68518 7606 68570
rect 7606 68518 7620 68570
rect 7644 68518 7658 68570
rect 7658 68518 7670 68570
rect 7670 68518 7700 68570
rect 7724 68518 7734 68570
rect 7734 68518 7780 68570
rect 7484 68516 7540 68518
rect 7564 68516 7620 68518
rect 7644 68516 7700 68518
rect 7724 68516 7780 68518
rect 5852 68026 5908 68028
rect 5932 68026 5988 68028
rect 6012 68026 6068 68028
rect 6092 68026 6148 68028
rect 5852 67974 5898 68026
rect 5898 67974 5908 68026
rect 5932 67974 5962 68026
rect 5962 67974 5974 68026
rect 5974 67974 5988 68026
rect 6012 67974 6026 68026
rect 6026 67974 6038 68026
rect 6038 67974 6068 68026
rect 6092 67974 6102 68026
rect 6102 67974 6148 68026
rect 5852 67972 5908 67974
rect 5932 67972 5988 67974
rect 6012 67972 6068 67974
rect 6092 67972 6148 67974
rect 7484 67482 7540 67484
rect 7564 67482 7620 67484
rect 7644 67482 7700 67484
rect 7724 67482 7780 67484
rect 7484 67430 7530 67482
rect 7530 67430 7540 67482
rect 7564 67430 7594 67482
rect 7594 67430 7606 67482
rect 7606 67430 7620 67482
rect 7644 67430 7658 67482
rect 7658 67430 7670 67482
rect 7670 67430 7700 67482
rect 7724 67430 7734 67482
rect 7734 67430 7780 67482
rect 7484 67428 7540 67430
rect 7564 67428 7620 67430
rect 7644 67428 7700 67430
rect 7724 67428 7780 67430
rect 5852 66938 5908 66940
rect 5932 66938 5988 66940
rect 6012 66938 6068 66940
rect 6092 66938 6148 66940
rect 5852 66886 5898 66938
rect 5898 66886 5908 66938
rect 5932 66886 5962 66938
rect 5962 66886 5974 66938
rect 5974 66886 5988 66938
rect 6012 66886 6026 66938
rect 6026 66886 6038 66938
rect 6038 66886 6068 66938
rect 6092 66886 6102 66938
rect 6102 66886 6148 66938
rect 5852 66884 5908 66886
rect 5932 66884 5988 66886
rect 6012 66884 6068 66886
rect 6092 66884 6148 66886
rect 7484 66394 7540 66396
rect 7564 66394 7620 66396
rect 7644 66394 7700 66396
rect 7724 66394 7780 66396
rect 7484 66342 7530 66394
rect 7530 66342 7540 66394
rect 7564 66342 7594 66394
rect 7594 66342 7606 66394
rect 7606 66342 7620 66394
rect 7644 66342 7658 66394
rect 7658 66342 7670 66394
rect 7670 66342 7700 66394
rect 7724 66342 7734 66394
rect 7734 66342 7780 66394
rect 7484 66340 7540 66342
rect 7564 66340 7620 66342
rect 7644 66340 7700 66342
rect 7724 66340 7780 66342
rect 5852 65850 5908 65852
rect 5932 65850 5988 65852
rect 6012 65850 6068 65852
rect 6092 65850 6148 65852
rect 5852 65798 5898 65850
rect 5898 65798 5908 65850
rect 5932 65798 5962 65850
rect 5962 65798 5974 65850
rect 5974 65798 5988 65850
rect 6012 65798 6026 65850
rect 6026 65798 6038 65850
rect 6038 65798 6068 65850
rect 6092 65798 6102 65850
rect 6102 65798 6148 65850
rect 5852 65796 5908 65798
rect 5932 65796 5988 65798
rect 6012 65796 6068 65798
rect 6092 65796 6148 65798
rect 9402 77152 9458 77208
rect 9116 76730 9172 76732
rect 9196 76730 9252 76732
rect 9276 76730 9332 76732
rect 9356 76730 9412 76732
rect 9116 76678 9162 76730
rect 9162 76678 9172 76730
rect 9196 76678 9226 76730
rect 9226 76678 9238 76730
rect 9238 76678 9252 76730
rect 9276 76678 9290 76730
rect 9290 76678 9302 76730
rect 9302 76678 9332 76730
rect 9356 76678 9366 76730
rect 9366 76678 9412 76730
rect 9116 76676 9172 76678
rect 9196 76676 9252 76678
rect 9276 76676 9332 76678
rect 9356 76676 9412 76678
rect 9116 75642 9172 75644
rect 9196 75642 9252 75644
rect 9276 75642 9332 75644
rect 9356 75642 9412 75644
rect 9116 75590 9162 75642
rect 9162 75590 9172 75642
rect 9196 75590 9226 75642
rect 9226 75590 9238 75642
rect 9238 75590 9252 75642
rect 9276 75590 9290 75642
rect 9290 75590 9302 75642
rect 9302 75590 9332 75642
rect 9356 75590 9366 75642
rect 9366 75590 9412 75642
rect 9116 75588 9172 75590
rect 9196 75588 9252 75590
rect 9276 75588 9332 75590
rect 9356 75588 9412 75590
rect 9116 74554 9172 74556
rect 9196 74554 9252 74556
rect 9276 74554 9332 74556
rect 9356 74554 9412 74556
rect 9116 74502 9162 74554
rect 9162 74502 9172 74554
rect 9196 74502 9226 74554
rect 9226 74502 9238 74554
rect 9238 74502 9252 74554
rect 9276 74502 9290 74554
rect 9290 74502 9302 74554
rect 9302 74502 9332 74554
rect 9356 74502 9366 74554
rect 9366 74502 9412 74554
rect 9116 74500 9172 74502
rect 9196 74500 9252 74502
rect 9276 74500 9332 74502
rect 9356 74500 9412 74502
rect 9116 73466 9172 73468
rect 9196 73466 9252 73468
rect 9276 73466 9332 73468
rect 9356 73466 9412 73468
rect 9116 73414 9162 73466
rect 9162 73414 9172 73466
rect 9196 73414 9226 73466
rect 9226 73414 9238 73466
rect 9238 73414 9252 73466
rect 9276 73414 9290 73466
rect 9290 73414 9302 73466
rect 9302 73414 9332 73466
rect 9356 73414 9366 73466
rect 9366 73414 9412 73466
rect 9116 73412 9172 73414
rect 9196 73412 9252 73414
rect 9276 73412 9332 73414
rect 9356 73412 9412 73414
rect 9116 72378 9172 72380
rect 9196 72378 9252 72380
rect 9276 72378 9332 72380
rect 9356 72378 9412 72380
rect 9116 72326 9162 72378
rect 9162 72326 9172 72378
rect 9196 72326 9226 72378
rect 9226 72326 9238 72378
rect 9238 72326 9252 72378
rect 9276 72326 9290 72378
rect 9290 72326 9302 72378
rect 9302 72326 9332 72378
rect 9356 72326 9366 72378
rect 9366 72326 9412 72378
rect 9116 72324 9172 72326
rect 9196 72324 9252 72326
rect 9276 72324 9332 72326
rect 9356 72324 9412 72326
rect 9116 71290 9172 71292
rect 9196 71290 9252 71292
rect 9276 71290 9332 71292
rect 9356 71290 9412 71292
rect 9116 71238 9162 71290
rect 9162 71238 9172 71290
rect 9196 71238 9226 71290
rect 9226 71238 9238 71290
rect 9238 71238 9252 71290
rect 9276 71238 9290 71290
rect 9290 71238 9302 71290
rect 9302 71238 9332 71290
rect 9356 71238 9366 71290
rect 9366 71238 9412 71290
rect 9116 71236 9172 71238
rect 9196 71236 9252 71238
rect 9276 71236 9332 71238
rect 9356 71236 9412 71238
rect 9116 70202 9172 70204
rect 9196 70202 9252 70204
rect 9276 70202 9332 70204
rect 9356 70202 9412 70204
rect 9116 70150 9162 70202
rect 9162 70150 9172 70202
rect 9196 70150 9226 70202
rect 9226 70150 9238 70202
rect 9238 70150 9252 70202
rect 9276 70150 9290 70202
rect 9290 70150 9302 70202
rect 9302 70150 9332 70202
rect 9356 70150 9366 70202
rect 9366 70150 9412 70202
rect 9116 70148 9172 70150
rect 9196 70148 9252 70150
rect 9276 70148 9332 70150
rect 9356 70148 9412 70150
rect 9116 69114 9172 69116
rect 9196 69114 9252 69116
rect 9276 69114 9332 69116
rect 9356 69114 9412 69116
rect 9116 69062 9162 69114
rect 9162 69062 9172 69114
rect 9196 69062 9226 69114
rect 9226 69062 9238 69114
rect 9238 69062 9252 69114
rect 9276 69062 9290 69114
rect 9290 69062 9302 69114
rect 9302 69062 9332 69114
rect 9356 69062 9366 69114
rect 9366 69062 9412 69114
rect 9116 69060 9172 69062
rect 9196 69060 9252 69062
rect 9276 69060 9332 69062
rect 9356 69060 9412 69062
rect 9116 68026 9172 68028
rect 9196 68026 9252 68028
rect 9276 68026 9332 68028
rect 9356 68026 9412 68028
rect 9116 67974 9162 68026
rect 9162 67974 9172 68026
rect 9196 67974 9226 68026
rect 9226 67974 9238 68026
rect 9238 67974 9252 68026
rect 9276 67974 9290 68026
rect 9290 67974 9302 68026
rect 9302 67974 9332 68026
rect 9356 67974 9366 68026
rect 9366 67974 9412 68026
rect 9116 67972 9172 67974
rect 9196 67972 9252 67974
rect 9276 67972 9332 67974
rect 9356 67972 9412 67974
rect 9116 66938 9172 66940
rect 9196 66938 9252 66940
rect 9276 66938 9332 66940
rect 9356 66938 9412 66940
rect 9116 66886 9162 66938
rect 9162 66886 9172 66938
rect 9196 66886 9226 66938
rect 9226 66886 9238 66938
rect 9238 66886 9252 66938
rect 9276 66886 9290 66938
rect 9290 66886 9302 66938
rect 9302 66886 9332 66938
rect 9356 66886 9366 66938
rect 9366 66886 9412 66938
rect 9116 66884 9172 66886
rect 9196 66884 9252 66886
rect 9276 66884 9332 66886
rect 9356 66884 9412 66886
rect 7484 65306 7540 65308
rect 7564 65306 7620 65308
rect 7644 65306 7700 65308
rect 7724 65306 7780 65308
rect 7484 65254 7530 65306
rect 7530 65254 7540 65306
rect 7564 65254 7594 65306
rect 7594 65254 7606 65306
rect 7606 65254 7620 65306
rect 7644 65254 7658 65306
rect 7658 65254 7670 65306
rect 7670 65254 7700 65306
rect 7724 65254 7734 65306
rect 7734 65254 7780 65306
rect 7484 65252 7540 65254
rect 7564 65252 7620 65254
rect 7644 65252 7700 65254
rect 7724 65252 7780 65254
rect 9116 65850 9172 65852
rect 9196 65850 9252 65852
rect 9276 65850 9332 65852
rect 9356 65850 9412 65852
rect 9116 65798 9162 65850
rect 9162 65798 9172 65850
rect 9196 65798 9226 65850
rect 9226 65798 9238 65850
rect 9238 65798 9252 65850
rect 9276 65798 9290 65850
rect 9290 65798 9302 65850
rect 9302 65798 9332 65850
rect 9356 65798 9366 65850
rect 9366 65798 9412 65850
rect 9116 65796 9172 65798
rect 9196 65796 9252 65798
rect 9276 65796 9332 65798
rect 9356 65796 9412 65798
rect 5852 64762 5908 64764
rect 5932 64762 5988 64764
rect 6012 64762 6068 64764
rect 6092 64762 6148 64764
rect 5852 64710 5898 64762
rect 5898 64710 5908 64762
rect 5932 64710 5962 64762
rect 5962 64710 5974 64762
rect 5974 64710 5988 64762
rect 6012 64710 6026 64762
rect 6026 64710 6038 64762
rect 6038 64710 6068 64762
rect 6092 64710 6102 64762
rect 6102 64710 6148 64762
rect 5852 64708 5908 64710
rect 5932 64708 5988 64710
rect 6012 64708 6068 64710
rect 6092 64708 6148 64710
rect 9116 64762 9172 64764
rect 9196 64762 9252 64764
rect 9276 64762 9332 64764
rect 9356 64762 9412 64764
rect 9116 64710 9162 64762
rect 9162 64710 9172 64762
rect 9196 64710 9226 64762
rect 9226 64710 9238 64762
rect 9238 64710 9252 64762
rect 9276 64710 9290 64762
rect 9290 64710 9302 64762
rect 9302 64710 9332 64762
rect 9356 64710 9366 64762
rect 9366 64710 9412 64762
rect 9116 64708 9172 64710
rect 9196 64708 9252 64710
rect 9276 64708 9332 64710
rect 9356 64708 9412 64710
rect 7484 64218 7540 64220
rect 7564 64218 7620 64220
rect 7644 64218 7700 64220
rect 7724 64218 7780 64220
rect 7484 64166 7530 64218
rect 7530 64166 7540 64218
rect 7564 64166 7594 64218
rect 7594 64166 7606 64218
rect 7606 64166 7620 64218
rect 7644 64166 7658 64218
rect 7658 64166 7670 64218
rect 7670 64166 7700 64218
rect 7724 64166 7734 64218
rect 7734 64166 7780 64218
rect 7484 64164 7540 64166
rect 7564 64164 7620 64166
rect 7644 64164 7700 64166
rect 7724 64164 7780 64166
rect 5852 63674 5908 63676
rect 5932 63674 5988 63676
rect 6012 63674 6068 63676
rect 6092 63674 6148 63676
rect 5852 63622 5898 63674
rect 5898 63622 5908 63674
rect 5932 63622 5962 63674
rect 5962 63622 5974 63674
rect 5974 63622 5988 63674
rect 6012 63622 6026 63674
rect 6026 63622 6038 63674
rect 6038 63622 6068 63674
rect 6092 63622 6102 63674
rect 6102 63622 6148 63674
rect 5852 63620 5908 63622
rect 5932 63620 5988 63622
rect 6012 63620 6068 63622
rect 6092 63620 6148 63622
rect 7484 63130 7540 63132
rect 7564 63130 7620 63132
rect 7644 63130 7700 63132
rect 7724 63130 7780 63132
rect 7484 63078 7530 63130
rect 7530 63078 7540 63130
rect 7564 63078 7594 63130
rect 7594 63078 7606 63130
rect 7606 63078 7620 63130
rect 7644 63078 7658 63130
rect 7658 63078 7670 63130
rect 7670 63078 7700 63130
rect 7724 63078 7734 63130
rect 7734 63078 7780 63130
rect 7484 63076 7540 63078
rect 7564 63076 7620 63078
rect 7644 63076 7700 63078
rect 7724 63076 7780 63078
rect 5852 62586 5908 62588
rect 5932 62586 5988 62588
rect 6012 62586 6068 62588
rect 6092 62586 6148 62588
rect 5852 62534 5898 62586
rect 5898 62534 5908 62586
rect 5932 62534 5962 62586
rect 5962 62534 5974 62586
rect 5974 62534 5988 62586
rect 6012 62534 6026 62586
rect 6026 62534 6038 62586
rect 6038 62534 6068 62586
rect 6092 62534 6102 62586
rect 6102 62534 6148 62586
rect 5852 62532 5908 62534
rect 5932 62532 5988 62534
rect 6012 62532 6068 62534
rect 6092 62532 6148 62534
rect 5852 61498 5908 61500
rect 5932 61498 5988 61500
rect 6012 61498 6068 61500
rect 6092 61498 6148 61500
rect 5852 61446 5898 61498
rect 5898 61446 5908 61498
rect 5932 61446 5962 61498
rect 5962 61446 5974 61498
rect 5974 61446 5988 61498
rect 6012 61446 6026 61498
rect 6026 61446 6038 61498
rect 6038 61446 6068 61498
rect 6092 61446 6102 61498
rect 6102 61446 6148 61498
rect 5852 61444 5908 61446
rect 5932 61444 5988 61446
rect 6012 61444 6068 61446
rect 6092 61444 6148 61446
rect 5852 60410 5908 60412
rect 5932 60410 5988 60412
rect 6012 60410 6068 60412
rect 6092 60410 6148 60412
rect 5852 60358 5898 60410
rect 5898 60358 5908 60410
rect 5932 60358 5962 60410
rect 5962 60358 5974 60410
rect 5974 60358 5988 60410
rect 6012 60358 6026 60410
rect 6026 60358 6038 60410
rect 6038 60358 6068 60410
rect 6092 60358 6102 60410
rect 6102 60358 6148 60410
rect 5852 60356 5908 60358
rect 5932 60356 5988 60358
rect 6012 60356 6068 60358
rect 6092 60356 6148 60358
rect 9116 63674 9172 63676
rect 9196 63674 9252 63676
rect 9276 63674 9332 63676
rect 9356 63674 9412 63676
rect 9116 63622 9162 63674
rect 9162 63622 9172 63674
rect 9196 63622 9226 63674
rect 9226 63622 9238 63674
rect 9238 63622 9252 63674
rect 9276 63622 9290 63674
rect 9290 63622 9302 63674
rect 9302 63622 9332 63674
rect 9356 63622 9366 63674
rect 9366 63622 9412 63674
rect 9116 63620 9172 63622
rect 9196 63620 9252 63622
rect 9276 63620 9332 63622
rect 9356 63620 9412 63622
rect 7484 62042 7540 62044
rect 7564 62042 7620 62044
rect 7644 62042 7700 62044
rect 7724 62042 7780 62044
rect 7484 61990 7530 62042
rect 7530 61990 7540 62042
rect 7564 61990 7594 62042
rect 7594 61990 7606 62042
rect 7606 61990 7620 62042
rect 7644 61990 7658 62042
rect 7658 61990 7670 62042
rect 7670 61990 7700 62042
rect 7724 61990 7734 62042
rect 7734 61990 7780 62042
rect 7484 61988 7540 61990
rect 7564 61988 7620 61990
rect 7644 61988 7700 61990
rect 7724 61988 7780 61990
rect 7484 60954 7540 60956
rect 7564 60954 7620 60956
rect 7644 60954 7700 60956
rect 7724 60954 7780 60956
rect 7484 60902 7530 60954
rect 7530 60902 7540 60954
rect 7564 60902 7594 60954
rect 7594 60902 7606 60954
rect 7606 60902 7620 60954
rect 7644 60902 7658 60954
rect 7658 60902 7670 60954
rect 7670 60902 7700 60954
rect 7724 60902 7734 60954
rect 7734 60902 7780 60954
rect 7484 60900 7540 60902
rect 7564 60900 7620 60902
rect 7644 60900 7700 60902
rect 7724 60900 7780 60902
rect 6182 60016 6238 60072
rect 7484 59866 7540 59868
rect 7564 59866 7620 59868
rect 7644 59866 7700 59868
rect 7724 59866 7780 59868
rect 7484 59814 7530 59866
rect 7530 59814 7540 59866
rect 7564 59814 7594 59866
rect 7594 59814 7606 59866
rect 7606 59814 7620 59866
rect 7644 59814 7658 59866
rect 7658 59814 7670 59866
rect 7670 59814 7700 59866
rect 7724 59814 7734 59866
rect 7734 59814 7780 59866
rect 7484 59812 7540 59814
rect 7564 59812 7620 59814
rect 7644 59812 7700 59814
rect 7724 59812 7780 59814
rect 5852 59322 5908 59324
rect 5932 59322 5988 59324
rect 6012 59322 6068 59324
rect 6092 59322 6148 59324
rect 5852 59270 5898 59322
rect 5898 59270 5908 59322
rect 5932 59270 5962 59322
rect 5962 59270 5974 59322
rect 5974 59270 5988 59322
rect 6012 59270 6026 59322
rect 6026 59270 6038 59322
rect 6038 59270 6068 59322
rect 6092 59270 6102 59322
rect 6102 59270 6148 59322
rect 5852 59268 5908 59270
rect 5932 59268 5988 59270
rect 6012 59268 6068 59270
rect 6092 59268 6148 59270
rect 7484 58778 7540 58780
rect 7564 58778 7620 58780
rect 7644 58778 7700 58780
rect 7724 58778 7780 58780
rect 7484 58726 7530 58778
rect 7530 58726 7540 58778
rect 7564 58726 7594 58778
rect 7594 58726 7606 58778
rect 7606 58726 7620 58778
rect 7644 58726 7658 58778
rect 7658 58726 7670 58778
rect 7670 58726 7700 58778
rect 7724 58726 7734 58778
rect 7734 58726 7780 58778
rect 7484 58724 7540 58726
rect 7564 58724 7620 58726
rect 7644 58724 7700 58726
rect 7724 58724 7780 58726
rect 5852 58234 5908 58236
rect 5932 58234 5988 58236
rect 6012 58234 6068 58236
rect 6092 58234 6148 58236
rect 5852 58182 5898 58234
rect 5898 58182 5908 58234
rect 5932 58182 5962 58234
rect 5962 58182 5974 58234
rect 5974 58182 5988 58234
rect 6012 58182 6026 58234
rect 6026 58182 6038 58234
rect 6038 58182 6068 58234
rect 6092 58182 6102 58234
rect 6102 58182 6148 58234
rect 5852 58180 5908 58182
rect 5932 58180 5988 58182
rect 6012 58180 6068 58182
rect 6092 58180 6148 58182
rect 7484 57690 7540 57692
rect 7564 57690 7620 57692
rect 7644 57690 7700 57692
rect 7724 57690 7780 57692
rect 7484 57638 7530 57690
rect 7530 57638 7540 57690
rect 7564 57638 7594 57690
rect 7594 57638 7606 57690
rect 7606 57638 7620 57690
rect 7644 57638 7658 57690
rect 7658 57638 7670 57690
rect 7670 57638 7700 57690
rect 7724 57638 7734 57690
rect 7734 57638 7780 57690
rect 7484 57636 7540 57638
rect 7564 57636 7620 57638
rect 7644 57636 7700 57638
rect 7724 57636 7780 57638
rect 5852 57146 5908 57148
rect 5932 57146 5988 57148
rect 6012 57146 6068 57148
rect 6092 57146 6148 57148
rect 5852 57094 5898 57146
rect 5898 57094 5908 57146
rect 5932 57094 5962 57146
rect 5962 57094 5974 57146
rect 5974 57094 5988 57146
rect 6012 57094 6026 57146
rect 6026 57094 6038 57146
rect 6038 57094 6068 57146
rect 6092 57094 6102 57146
rect 6102 57094 6148 57146
rect 5852 57092 5908 57094
rect 5932 57092 5988 57094
rect 6012 57092 6068 57094
rect 6092 57092 6148 57094
rect 5852 56058 5908 56060
rect 5932 56058 5988 56060
rect 6012 56058 6068 56060
rect 6092 56058 6148 56060
rect 5852 56006 5898 56058
rect 5898 56006 5908 56058
rect 5932 56006 5962 56058
rect 5962 56006 5974 56058
rect 5974 56006 5988 56058
rect 6012 56006 6026 56058
rect 6026 56006 6038 56058
rect 6038 56006 6068 56058
rect 6092 56006 6102 56058
rect 6102 56006 6148 56058
rect 5852 56004 5908 56006
rect 5932 56004 5988 56006
rect 6012 56004 6068 56006
rect 6092 56004 6148 56006
rect 5852 54970 5908 54972
rect 5932 54970 5988 54972
rect 6012 54970 6068 54972
rect 6092 54970 6148 54972
rect 5852 54918 5898 54970
rect 5898 54918 5908 54970
rect 5932 54918 5962 54970
rect 5962 54918 5974 54970
rect 5974 54918 5988 54970
rect 6012 54918 6026 54970
rect 6026 54918 6038 54970
rect 6038 54918 6068 54970
rect 6092 54918 6102 54970
rect 6102 54918 6148 54970
rect 5852 54916 5908 54918
rect 5932 54916 5988 54918
rect 6012 54916 6068 54918
rect 6092 54916 6148 54918
rect 5852 53882 5908 53884
rect 5932 53882 5988 53884
rect 6012 53882 6068 53884
rect 6092 53882 6148 53884
rect 5852 53830 5898 53882
rect 5898 53830 5908 53882
rect 5932 53830 5962 53882
rect 5962 53830 5974 53882
rect 5974 53830 5988 53882
rect 6012 53830 6026 53882
rect 6026 53830 6038 53882
rect 6038 53830 6068 53882
rect 6092 53830 6102 53882
rect 6102 53830 6148 53882
rect 5852 53828 5908 53830
rect 5932 53828 5988 53830
rect 6012 53828 6068 53830
rect 6092 53828 6148 53830
rect 5852 52794 5908 52796
rect 5932 52794 5988 52796
rect 6012 52794 6068 52796
rect 6092 52794 6148 52796
rect 5852 52742 5898 52794
rect 5898 52742 5908 52794
rect 5932 52742 5962 52794
rect 5962 52742 5974 52794
rect 5974 52742 5988 52794
rect 6012 52742 6026 52794
rect 6026 52742 6038 52794
rect 6038 52742 6068 52794
rect 6092 52742 6102 52794
rect 6102 52742 6148 52794
rect 5852 52740 5908 52742
rect 5932 52740 5988 52742
rect 6012 52740 6068 52742
rect 6092 52740 6148 52742
rect 5852 51706 5908 51708
rect 5932 51706 5988 51708
rect 6012 51706 6068 51708
rect 6092 51706 6148 51708
rect 5852 51654 5898 51706
rect 5898 51654 5908 51706
rect 5932 51654 5962 51706
rect 5962 51654 5974 51706
rect 5974 51654 5988 51706
rect 6012 51654 6026 51706
rect 6026 51654 6038 51706
rect 6038 51654 6068 51706
rect 6092 51654 6102 51706
rect 6102 51654 6148 51706
rect 5852 51652 5908 51654
rect 5932 51652 5988 51654
rect 6012 51652 6068 51654
rect 6092 51652 6148 51654
rect 5852 50618 5908 50620
rect 5932 50618 5988 50620
rect 6012 50618 6068 50620
rect 6092 50618 6148 50620
rect 5852 50566 5898 50618
rect 5898 50566 5908 50618
rect 5932 50566 5962 50618
rect 5962 50566 5974 50618
rect 5974 50566 5988 50618
rect 6012 50566 6026 50618
rect 6026 50566 6038 50618
rect 6038 50566 6068 50618
rect 6092 50566 6102 50618
rect 6102 50566 6148 50618
rect 5852 50564 5908 50566
rect 5932 50564 5988 50566
rect 6012 50564 6068 50566
rect 6092 50564 6148 50566
rect 5852 49530 5908 49532
rect 5932 49530 5988 49532
rect 6012 49530 6068 49532
rect 6092 49530 6148 49532
rect 5852 49478 5898 49530
rect 5898 49478 5908 49530
rect 5932 49478 5962 49530
rect 5962 49478 5974 49530
rect 5974 49478 5988 49530
rect 6012 49478 6026 49530
rect 6026 49478 6038 49530
rect 6038 49478 6068 49530
rect 6092 49478 6102 49530
rect 6102 49478 6148 49530
rect 5852 49476 5908 49478
rect 5932 49476 5988 49478
rect 6012 49476 6068 49478
rect 6092 49476 6148 49478
rect 5852 48442 5908 48444
rect 5932 48442 5988 48444
rect 6012 48442 6068 48444
rect 6092 48442 6148 48444
rect 5852 48390 5898 48442
rect 5898 48390 5908 48442
rect 5932 48390 5962 48442
rect 5962 48390 5974 48442
rect 5974 48390 5988 48442
rect 6012 48390 6026 48442
rect 6026 48390 6038 48442
rect 6038 48390 6068 48442
rect 6092 48390 6102 48442
rect 6102 48390 6148 48442
rect 5852 48388 5908 48390
rect 5932 48388 5988 48390
rect 6012 48388 6068 48390
rect 6092 48388 6148 48390
rect 5852 47354 5908 47356
rect 5932 47354 5988 47356
rect 6012 47354 6068 47356
rect 6092 47354 6148 47356
rect 5852 47302 5898 47354
rect 5898 47302 5908 47354
rect 5932 47302 5962 47354
rect 5962 47302 5974 47354
rect 5974 47302 5988 47354
rect 6012 47302 6026 47354
rect 6026 47302 6038 47354
rect 6038 47302 6068 47354
rect 6092 47302 6102 47354
rect 6102 47302 6148 47354
rect 5852 47300 5908 47302
rect 5932 47300 5988 47302
rect 6012 47300 6068 47302
rect 6092 47300 6148 47302
rect 5538 45600 5594 45656
rect 5852 46266 5908 46268
rect 5932 46266 5988 46268
rect 6012 46266 6068 46268
rect 6092 46266 6148 46268
rect 5852 46214 5898 46266
rect 5898 46214 5908 46266
rect 5932 46214 5962 46266
rect 5962 46214 5974 46266
rect 5974 46214 5988 46266
rect 6012 46214 6026 46266
rect 6026 46214 6038 46266
rect 6038 46214 6068 46266
rect 6092 46214 6102 46266
rect 6102 46214 6148 46266
rect 5852 46212 5908 46214
rect 5932 46212 5988 46214
rect 6012 46212 6068 46214
rect 6092 46212 6148 46214
rect 5852 45178 5908 45180
rect 5932 45178 5988 45180
rect 6012 45178 6068 45180
rect 6092 45178 6148 45180
rect 5852 45126 5898 45178
rect 5898 45126 5908 45178
rect 5932 45126 5962 45178
rect 5962 45126 5974 45178
rect 5974 45126 5988 45178
rect 6012 45126 6026 45178
rect 6026 45126 6038 45178
rect 6038 45126 6068 45178
rect 6092 45126 6102 45178
rect 6102 45126 6148 45178
rect 5852 45124 5908 45126
rect 5932 45124 5988 45126
rect 6012 45124 6068 45126
rect 6092 45124 6148 45126
rect 5852 44090 5908 44092
rect 5932 44090 5988 44092
rect 6012 44090 6068 44092
rect 6092 44090 6148 44092
rect 5852 44038 5898 44090
rect 5898 44038 5908 44090
rect 5932 44038 5962 44090
rect 5962 44038 5974 44090
rect 5974 44038 5988 44090
rect 6012 44038 6026 44090
rect 6026 44038 6038 44090
rect 6038 44038 6068 44090
rect 6092 44038 6102 44090
rect 6102 44038 6148 44090
rect 5852 44036 5908 44038
rect 5932 44036 5988 44038
rect 6012 44036 6068 44038
rect 6092 44036 6148 44038
rect 5852 43002 5908 43004
rect 5932 43002 5988 43004
rect 6012 43002 6068 43004
rect 6092 43002 6148 43004
rect 5852 42950 5898 43002
rect 5898 42950 5908 43002
rect 5932 42950 5962 43002
rect 5962 42950 5974 43002
rect 5974 42950 5988 43002
rect 6012 42950 6026 43002
rect 6026 42950 6038 43002
rect 6038 42950 6068 43002
rect 6092 42950 6102 43002
rect 6102 42950 6148 43002
rect 5852 42948 5908 42950
rect 5932 42948 5988 42950
rect 6012 42948 6068 42950
rect 6092 42948 6148 42950
rect 5852 41914 5908 41916
rect 5932 41914 5988 41916
rect 6012 41914 6068 41916
rect 6092 41914 6148 41916
rect 5852 41862 5898 41914
rect 5898 41862 5908 41914
rect 5932 41862 5962 41914
rect 5962 41862 5974 41914
rect 5974 41862 5988 41914
rect 6012 41862 6026 41914
rect 6026 41862 6038 41914
rect 6038 41862 6068 41914
rect 6092 41862 6102 41914
rect 6102 41862 6148 41914
rect 5852 41860 5908 41862
rect 5932 41860 5988 41862
rect 6012 41860 6068 41862
rect 6092 41860 6148 41862
rect 5852 40826 5908 40828
rect 5932 40826 5988 40828
rect 6012 40826 6068 40828
rect 6092 40826 6148 40828
rect 5852 40774 5898 40826
rect 5898 40774 5908 40826
rect 5932 40774 5962 40826
rect 5962 40774 5974 40826
rect 5974 40774 5988 40826
rect 6012 40774 6026 40826
rect 6026 40774 6038 40826
rect 6038 40774 6068 40826
rect 6092 40774 6102 40826
rect 6102 40774 6148 40826
rect 5852 40772 5908 40774
rect 5932 40772 5988 40774
rect 6012 40772 6068 40774
rect 6092 40772 6148 40774
rect 5852 39738 5908 39740
rect 5932 39738 5988 39740
rect 6012 39738 6068 39740
rect 6092 39738 6148 39740
rect 5852 39686 5898 39738
rect 5898 39686 5908 39738
rect 5932 39686 5962 39738
rect 5962 39686 5974 39738
rect 5974 39686 5988 39738
rect 6012 39686 6026 39738
rect 6026 39686 6038 39738
rect 6038 39686 6068 39738
rect 6092 39686 6102 39738
rect 6102 39686 6148 39738
rect 5852 39684 5908 39686
rect 5932 39684 5988 39686
rect 6012 39684 6068 39686
rect 6092 39684 6148 39686
rect 5852 38650 5908 38652
rect 5932 38650 5988 38652
rect 6012 38650 6068 38652
rect 6092 38650 6148 38652
rect 5852 38598 5898 38650
rect 5898 38598 5908 38650
rect 5932 38598 5962 38650
rect 5962 38598 5974 38650
rect 5974 38598 5988 38650
rect 6012 38598 6026 38650
rect 6026 38598 6038 38650
rect 6038 38598 6068 38650
rect 6092 38598 6102 38650
rect 6102 38598 6148 38650
rect 5852 38596 5908 38598
rect 5932 38596 5988 38598
rect 6012 38596 6068 38598
rect 6092 38596 6148 38598
rect 5852 37562 5908 37564
rect 5932 37562 5988 37564
rect 6012 37562 6068 37564
rect 6092 37562 6148 37564
rect 5852 37510 5898 37562
rect 5898 37510 5908 37562
rect 5932 37510 5962 37562
rect 5962 37510 5974 37562
rect 5974 37510 5988 37562
rect 6012 37510 6026 37562
rect 6026 37510 6038 37562
rect 6038 37510 6068 37562
rect 6092 37510 6102 37562
rect 6102 37510 6148 37562
rect 5852 37508 5908 37510
rect 5932 37508 5988 37510
rect 6012 37508 6068 37510
rect 6092 37508 6148 37510
rect 5852 36474 5908 36476
rect 5932 36474 5988 36476
rect 6012 36474 6068 36476
rect 6092 36474 6148 36476
rect 5852 36422 5898 36474
rect 5898 36422 5908 36474
rect 5932 36422 5962 36474
rect 5962 36422 5974 36474
rect 5974 36422 5988 36474
rect 6012 36422 6026 36474
rect 6026 36422 6038 36474
rect 6038 36422 6068 36474
rect 6092 36422 6102 36474
rect 6102 36422 6148 36474
rect 5852 36420 5908 36422
rect 5932 36420 5988 36422
rect 6012 36420 6068 36422
rect 6092 36420 6148 36422
rect 5852 35386 5908 35388
rect 5932 35386 5988 35388
rect 6012 35386 6068 35388
rect 6092 35386 6148 35388
rect 5852 35334 5898 35386
rect 5898 35334 5908 35386
rect 5932 35334 5962 35386
rect 5962 35334 5974 35386
rect 5974 35334 5988 35386
rect 6012 35334 6026 35386
rect 6026 35334 6038 35386
rect 6038 35334 6068 35386
rect 6092 35334 6102 35386
rect 6102 35334 6148 35386
rect 5852 35332 5908 35334
rect 5932 35332 5988 35334
rect 6012 35332 6068 35334
rect 6092 35332 6148 35334
rect 5852 34298 5908 34300
rect 5932 34298 5988 34300
rect 6012 34298 6068 34300
rect 6092 34298 6148 34300
rect 5852 34246 5898 34298
rect 5898 34246 5908 34298
rect 5932 34246 5962 34298
rect 5962 34246 5974 34298
rect 5974 34246 5988 34298
rect 6012 34246 6026 34298
rect 6026 34246 6038 34298
rect 6038 34246 6068 34298
rect 6092 34246 6102 34298
rect 6102 34246 6148 34298
rect 5852 34244 5908 34246
rect 5932 34244 5988 34246
rect 6012 34244 6068 34246
rect 6092 34244 6148 34246
rect 5852 33210 5908 33212
rect 5932 33210 5988 33212
rect 6012 33210 6068 33212
rect 6092 33210 6148 33212
rect 5852 33158 5898 33210
rect 5898 33158 5908 33210
rect 5932 33158 5962 33210
rect 5962 33158 5974 33210
rect 5974 33158 5988 33210
rect 6012 33158 6026 33210
rect 6026 33158 6038 33210
rect 6038 33158 6068 33210
rect 6092 33158 6102 33210
rect 6102 33158 6148 33210
rect 5852 33156 5908 33158
rect 5932 33156 5988 33158
rect 6012 33156 6068 33158
rect 6092 33156 6148 33158
rect 5630 32136 5686 32192
rect 5538 31592 5594 31648
rect 5538 31048 5594 31104
rect 5446 28192 5502 28248
rect 5852 32122 5908 32124
rect 5932 32122 5988 32124
rect 6012 32122 6068 32124
rect 6092 32122 6148 32124
rect 5852 32070 5898 32122
rect 5898 32070 5908 32122
rect 5932 32070 5962 32122
rect 5962 32070 5974 32122
rect 5974 32070 5988 32122
rect 6012 32070 6026 32122
rect 6026 32070 6038 32122
rect 6038 32070 6068 32122
rect 6092 32070 6102 32122
rect 6102 32070 6148 32122
rect 5852 32068 5908 32070
rect 5932 32068 5988 32070
rect 6012 32068 6068 32070
rect 6092 32068 6148 32070
rect 5852 31034 5908 31036
rect 5932 31034 5988 31036
rect 6012 31034 6068 31036
rect 6092 31034 6148 31036
rect 5852 30982 5898 31034
rect 5898 30982 5908 31034
rect 5932 30982 5962 31034
rect 5962 30982 5974 31034
rect 5974 30982 5988 31034
rect 6012 30982 6026 31034
rect 6026 30982 6038 31034
rect 6038 30982 6068 31034
rect 6092 30982 6102 31034
rect 6102 30982 6148 31034
rect 5852 30980 5908 30982
rect 5932 30980 5988 30982
rect 6012 30980 6068 30982
rect 6092 30980 6148 30982
rect 5852 29946 5908 29948
rect 5932 29946 5988 29948
rect 6012 29946 6068 29948
rect 6092 29946 6148 29948
rect 5852 29894 5898 29946
rect 5898 29894 5908 29946
rect 5932 29894 5962 29946
rect 5962 29894 5974 29946
rect 5974 29894 5988 29946
rect 6012 29894 6026 29946
rect 6026 29894 6038 29946
rect 6038 29894 6068 29946
rect 6092 29894 6102 29946
rect 6102 29894 6148 29946
rect 5852 29892 5908 29894
rect 5932 29892 5988 29894
rect 6012 29892 6068 29894
rect 6092 29892 6148 29894
rect 5852 28858 5908 28860
rect 5932 28858 5988 28860
rect 6012 28858 6068 28860
rect 6092 28858 6148 28860
rect 5852 28806 5898 28858
rect 5898 28806 5908 28858
rect 5932 28806 5962 28858
rect 5962 28806 5974 28858
rect 5974 28806 5988 28858
rect 6012 28806 6026 28858
rect 6026 28806 6038 28858
rect 6038 28806 6068 28858
rect 6092 28806 6102 28858
rect 6102 28806 6148 28858
rect 5852 28804 5908 28806
rect 5932 28804 5988 28806
rect 6012 28804 6068 28806
rect 6092 28804 6148 28806
rect 5852 27770 5908 27772
rect 5932 27770 5988 27772
rect 6012 27770 6068 27772
rect 6092 27770 6148 27772
rect 5852 27718 5898 27770
rect 5898 27718 5908 27770
rect 5932 27718 5962 27770
rect 5962 27718 5974 27770
rect 5974 27718 5988 27770
rect 6012 27718 6026 27770
rect 6026 27718 6038 27770
rect 6038 27718 6068 27770
rect 6092 27718 6102 27770
rect 6102 27718 6148 27770
rect 5852 27716 5908 27718
rect 5932 27716 5988 27718
rect 6012 27716 6068 27718
rect 6092 27716 6148 27718
rect 5852 26682 5908 26684
rect 5932 26682 5988 26684
rect 6012 26682 6068 26684
rect 6092 26682 6148 26684
rect 5852 26630 5898 26682
rect 5898 26630 5908 26682
rect 5932 26630 5962 26682
rect 5962 26630 5974 26682
rect 5974 26630 5988 26682
rect 6012 26630 6026 26682
rect 6026 26630 6038 26682
rect 6038 26630 6068 26682
rect 6092 26630 6102 26682
rect 6102 26630 6148 26682
rect 5852 26628 5908 26630
rect 5932 26628 5988 26630
rect 6012 26628 6068 26630
rect 6092 26628 6148 26630
rect 9116 62586 9172 62588
rect 9196 62586 9252 62588
rect 9276 62586 9332 62588
rect 9356 62586 9412 62588
rect 9116 62534 9162 62586
rect 9162 62534 9172 62586
rect 9196 62534 9226 62586
rect 9226 62534 9238 62586
rect 9238 62534 9252 62586
rect 9276 62534 9290 62586
rect 9290 62534 9302 62586
rect 9302 62534 9332 62586
rect 9356 62534 9366 62586
rect 9366 62534 9412 62586
rect 9116 62532 9172 62534
rect 9196 62532 9252 62534
rect 9276 62532 9332 62534
rect 9356 62532 9412 62534
rect 9116 61498 9172 61500
rect 9196 61498 9252 61500
rect 9276 61498 9332 61500
rect 9356 61498 9412 61500
rect 9116 61446 9162 61498
rect 9162 61446 9172 61498
rect 9196 61446 9226 61498
rect 9226 61446 9238 61498
rect 9238 61446 9252 61498
rect 9276 61446 9290 61498
rect 9290 61446 9302 61498
rect 9302 61446 9332 61498
rect 9356 61446 9366 61498
rect 9366 61446 9412 61498
rect 9116 61444 9172 61446
rect 9196 61444 9252 61446
rect 9276 61444 9332 61446
rect 9356 61444 9412 61446
rect 9116 60410 9172 60412
rect 9196 60410 9252 60412
rect 9276 60410 9332 60412
rect 9356 60410 9412 60412
rect 9116 60358 9162 60410
rect 9162 60358 9172 60410
rect 9196 60358 9226 60410
rect 9226 60358 9238 60410
rect 9238 60358 9252 60410
rect 9276 60358 9290 60410
rect 9290 60358 9302 60410
rect 9302 60358 9332 60410
rect 9356 60358 9366 60410
rect 9366 60358 9412 60410
rect 9116 60356 9172 60358
rect 9196 60356 9252 60358
rect 9276 60356 9332 60358
rect 9356 60356 9412 60358
rect 9116 59322 9172 59324
rect 9196 59322 9252 59324
rect 9276 59322 9332 59324
rect 9356 59322 9412 59324
rect 9116 59270 9162 59322
rect 9162 59270 9172 59322
rect 9196 59270 9226 59322
rect 9226 59270 9238 59322
rect 9238 59270 9252 59322
rect 9276 59270 9290 59322
rect 9290 59270 9302 59322
rect 9302 59270 9332 59322
rect 9356 59270 9366 59322
rect 9366 59270 9412 59322
rect 9116 59268 9172 59270
rect 9196 59268 9252 59270
rect 9276 59268 9332 59270
rect 9356 59268 9412 59270
rect 9116 58234 9172 58236
rect 9196 58234 9252 58236
rect 9276 58234 9332 58236
rect 9356 58234 9412 58236
rect 9116 58182 9162 58234
rect 9162 58182 9172 58234
rect 9196 58182 9226 58234
rect 9226 58182 9238 58234
rect 9238 58182 9252 58234
rect 9276 58182 9290 58234
rect 9290 58182 9302 58234
rect 9302 58182 9332 58234
rect 9356 58182 9366 58234
rect 9366 58182 9412 58234
rect 9116 58180 9172 58182
rect 9196 58180 9252 58182
rect 9276 58180 9332 58182
rect 9356 58180 9412 58182
rect 9494 57976 9550 58032
rect 9494 57160 9550 57216
rect 9116 57146 9172 57148
rect 9196 57146 9252 57148
rect 9276 57146 9332 57148
rect 9356 57146 9412 57148
rect 9116 57094 9162 57146
rect 9162 57094 9172 57146
rect 9196 57094 9226 57146
rect 9226 57094 9238 57146
rect 9238 57094 9252 57146
rect 9276 57094 9290 57146
rect 9290 57094 9302 57146
rect 9302 57094 9332 57146
rect 9356 57094 9366 57146
rect 9366 57094 9412 57146
rect 9116 57092 9172 57094
rect 9196 57092 9252 57094
rect 9276 57092 9332 57094
rect 9356 57092 9412 57094
rect 7484 56602 7540 56604
rect 7564 56602 7620 56604
rect 7644 56602 7700 56604
rect 7724 56602 7780 56604
rect 7484 56550 7530 56602
rect 7530 56550 7540 56602
rect 7564 56550 7594 56602
rect 7594 56550 7606 56602
rect 7606 56550 7620 56602
rect 7644 56550 7658 56602
rect 7658 56550 7670 56602
rect 7670 56550 7700 56602
rect 7724 56550 7734 56602
rect 7734 56550 7780 56602
rect 7484 56548 7540 56550
rect 7564 56548 7620 56550
rect 7644 56548 7700 56550
rect 7724 56548 7780 56550
rect 7484 55514 7540 55516
rect 7564 55514 7620 55516
rect 7644 55514 7700 55516
rect 7724 55514 7780 55516
rect 7484 55462 7530 55514
rect 7530 55462 7540 55514
rect 7564 55462 7594 55514
rect 7594 55462 7606 55514
rect 7606 55462 7620 55514
rect 7644 55462 7658 55514
rect 7658 55462 7670 55514
rect 7670 55462 7700 55514
rect 7724 55462 7734 55514
rect 7734 55462 7780 55514
rect 7484 55460 7540 55462
rect 7564 55460 7620 55462
rect 7644 55460 7700 55462
rect 7724 55460 7780 55462
rect 7484 54426 7540 54428
rect 7564 54426 7620 54428
rect 7644 54426 7700 54428
rect 7724 54426 7780 54428
rect 7484 54374 7530 54426
rect 7530 54374 7540 54426
rect 7564 54374 7594 54426
rect 7594 54374 7606 54426
rect 7606 54374 7620 54426
rect 7644 54374 7658 54426
rect 7658 54374 7670 54426
rect 7670 54374 7700 54426
rect 7724 54374 7734 54426
rect 7734 54374 7780 54426
rect 7484 54372 7540 54374
rect 7564 54372 7620 54374
rect 7644 54372 7700 54374
rect 7724 54372 7780 54374
rect 7484 53338 7540 53340
rect 7564 53338 7620 53340
rect 7644 53338 7700 53340
rect 7724 53338 7780 53340
rect 7484 53286 7530 53338
rect 7530 53286 7540 53338
rect 7564 53286 7594 53338
rect 7594 53286 7606 53338
rect 7606 53286 7620 53338
rect 7644 53286 7658 53338
rect 7658 53286 7670 53338
rect 7670 53286 7700 53338
rect 7724 53286 7734 53338
rect 7734 53286 7780 53338
rect 7484 53284 7540 53286
rect 7564 53284 7620 53286
rect 7644 53284 7700 53286
rect 7724 53284 7780 53286
rect 6550 49816 6606 49872
rect 6734 41248 6790 41304
rect 7484 52250 7540 52252
rect 7564 52250 7620 52252
rect 7644 52250 7700 52252
rect 7724 52250 7780 52252
rect 7484 52198 7530 52250
rect 7530 52198 7540 52250
rect 7564 52198 7594 52250
rect 7594 52198 7606 52250
rect 7606 52198 7620 52250
rect 7644 52198 7658 52250
rect 7658 52198 7670 52250
rect 7670 52198 7700 52250
rect 7724 52198 7734 52250
rect 7734 52198 7780 52250
rect 7484 52196 7540 52198
rect 7564 52196 7620 52198
rect 7644 52196 7700 52198
rect 7724 52196 7780 52198
rect 7484 51162 7540 51164
rect 7564 51162 7620 51164
rect 7644 51162 7700 51164
rect 7724 51162 7780 51164
rect 7484 51110 7530 51162
rect 7530 51110 7540 51162
rect 7564 51110 7594 51162
rect 7594 51110 7606 51162
rect 7606 51110 7620 51162
rect 7644 51110 7658 51162
rect 7658 51110 7670 51162
rect 7670 51110 7700 51162
rect 7724 51110 7734 51162
rect 7734 51110 7780 51162
rect 7484 51108 7540 51110
rect 7564 51108 7620 51110
rect 7644 51108 7700 51110
rect 7724 51108 7780 51110
rect 9310 56344 9366 56400
rect 9116 56058 9172 56060
rect 9196 56058 9252 56060
rect 9276 56058 9332 56060
rect 9356 56058 9412 56060
rect 9116 56006 9162 56058
rect 9162 56006 9172 56058
rect 9196 56006 9226 56058
rect 9226 56006 9238 56058
rect 9238 56006 9252 56058
rect 9276 56006 9290 56058
rect 9290 56006 9302 56058
rect 9302 56006 9332 56058
rect 9356 56006 9366 56058
rect 9366 56006 9412 56058
rect 9116 56004 9172 56006
rect 9196 56004 9252 56006
rect 9276 56004 9332 56006
rect 9356 56004 9412 56006
rect 9116 54970 9172 54972
rect 9196 54970 9252 54972
rect 9276 54970 9332 54972
rect 9356 54970 9412 54972
rect 9116 54918 9162 54970
rect 9162 54918 9172 54970
rect 9196 54918 9226 54970
rect 9226 54918 9238 54970
rect 9238 54918 9252 54970
rect 9276 54918 9290 54970
rect 9290 54918 9302 54970
rect 9302 54918 9332 54970
rect 9356 54918 9366 54970
rect 9366 54918 9412 54970
rect 9116 54916 9172 54918
rect 9196 54916 9252 54918
rect 9276 54916 9332 54918
rect 9356 54916 9412 54918
rect 9586 54848 9642 54904
rect 9116 53882 9172 53884
rect 9196 53882 9252 53884
rect 9276 53882 9332 53884
rect 9356 53882 9412 53884
rect 9116 53830 9162 53882
rect 9162 53830 9172 53882
rect 9196 53830 9226 53882
rect 9226 53830 9238 53882
rect 9238 53830 9252 53882
rect 9276 53830 9290 53882
rect 9290 53830 9302 53882
rect 9302 53830 9332 53882
rect 9356 53830 9366 53882
rect 9366 53830 9412 53882
rect 9116 53828 9172 53830
rect 9196 53828 9252 53830
rect 9276 53828 9332 53830
rect 9356 53828 9412 53830
rect 9116 52794 9172 52796
rect 9196 52794 9252 52796
rect 9276 52794 9332 52796
rect 9356 52794 9412 52796
rect 9116 52742 9162 52794
rect 9162 52742 9172 52794
rect 9196 52742 9226 52794
rect 9226 52742 9238 52794
rect 9238 52742 9252 52794
rect 9276 52742 9290 52794
rect 9290 52742 9302 52794
rect 9302 52742 9332 52794
rect 9356 52742 9366 52794
rect 9366 52742 9412 52794
rect 9116 52740 9172 52742
rect 9196 52740 9252 52742
rect 9276 52740 9332 52742
rect 9356 52740 9412 52742
rect 9116 51706 9172 51708
rect 9196 51706 9252 51708
rect 9276 51706 9332 51708
rect 9356 51706 9412 51708
rect 9116 51654 9162 51706
rect 9162 51654 9172 51706
rect 9196 51654 9226 51706
rect 9226 51654 9238 51706
rect 9238 51654 9252 51706
rect 9276 51654 9290 51706
rect 9290 51654 9302 51706
rect 9302 51654 9332 51706
rect 9356 51654 9366 51706
rect 9366 51654 9412 51706
rect 9116 51652 9172 51654
rect 9196 51652 9252 51654
rect 9276 51652 9332 51654
rect 9356 51652 9412 51654
rect 9116 50618 9172 50620
rect 9196 50618 9252 50620
rect 9276 50618 9332 50620
rect 9356 50618 9412 50620
rect 9116 50566 9162 50618
rect 9162 50566 9172 50618
rect 9196 50566 9226 50618
rect 9226 50566 9238 50618
rect 9238 50566 9252 50618
rect 9276 50566 9290 50618
rect 9290 50566 9302 50618
rect 9302 50566 9332 50618
rect 9356 50566 9366 50618
rect 9366 50566 9412 50618
rect 9116 50564 9172 50566
rect 9196 50564 9252 50566
rect 9276 50564 9332 50566
rect 9356 50564 9412 50566
rect 7484 50074 7540 50076
rect 7564 50074 7620 50076
rect 7644 50074 7700 50076
rect 7724 50074 7780 50076
rect 7484 50022 7530 50074
rect 7530 50022 7540 50074
rect 7564 50022 7594 50074
rect 7594 50022 7606 50074
rect 7606 50022 7620 50074
rect 7644 50022 7658 50074
rect 7658 50022 7670 50074
rect 7670 50022 7700 50074
rect 7724 50022 7734 50074
rect 7734 50022 7780 50074
rect 7484 50020 7540 50022
rect 7564 50020 7620 50022
rect 7644 50020 7700 50022
rect 7724 50020 7780 50022
rect 9116 49530 9172 49532
rect 9196 49530 9252 49532
rect 9276 49530 9332 49532
rect 9356 49530 9412 49532
rect 9116 49478 9162 49530
rect 9162 49478 9172 49530
rect 9196 49478 9226 49530
rect 9226 49478 9238 49530
rect 9238 49478 9252 49530
rect 9276 49478 9290 49530
rect 9290 49478 9302 49530
rect 9302 49478 9332 49530
rect 9356 49478 9366 49530
rect 9366 49478 9412 49530
rect 9116 49476 9172 49478
rect 9196 49476 9252 49478
rect 9276 49476 9332 49478
rect 9356 49476 9412 49478
rect 9586 49408 9642 49464
rect 7484 48986 7540 48988
rect 7564 48986 7620 48988
rect 7644 48986 7700 48988
rect 7724 48986 7780 48988
rect 7484 48934 7530 48986
rect 7530 48934 7540 48986
rect 7564 48934 7594 48986
rect 7594 48934 7606 48986
rect 7606 48934 7620 48986
rect 7644 48934 7658 48986
rect 7658 48934 7670 48986
rect 7670 48934 7700 48986
rect 7724 48934 7734 48986
rect 7734 48934 7780 48986
rect 7484 48932 7540 48934
rect 7564 48932 7620 48934
rect 7644 48932 7700 48934
rect 7724 48932 7780 48934
rect 9116 48442 9172 48444
rect 9196 48442 9252 48444
rect 9276 48442 9332 48444
rect 9356 48442 9412 48444
rect 9116 48390 9162 48442
rect 9162 48390 9172 48442
rect 9196 48390 9226 48442
rect 9226 48390 9238 48442
rect 9238 48390 9252 48442
rect 9276 48390 9290 48442
rect 9290 48390 9302 48442
rect 9302 48390 9332 48442
rect 9356 48390 9366 48442
rect 9366 48390 9412 48442
rect 9116 48388 9172 48390
rect 9196 48388 9252 48390
rect 9276 48388 9332 48390
rect 9356 48388 9412 48390
rect 7484 47898 7540 47900
rect 7564 47898 7620 47900
rect 7644 47898 7700 47900
rect 7724 47898 7780 47900
rect 7484 47846 7530 47898
rect 7530 47846 7540 47898
rect 7564 47846 7594 47898
rect 7594 47846 7606 47898
rect 7606 47846 7620 47898
rect 7644 47846 7658 47898
rect 7658 47846 7670 47898
rect 7670 47846 7700 47898
rect 7724 47846 7734 47898
rect 7734 47846 7780 47898
rect 7484 47844 7540 47846
rect 7564 47844 7620 47846
rect 7644 47844 7700 47846
rect 7724 47844 7780 47846
rect 9116 47354 9172 47356
rect 9196 47354 9252 47356
rect 9276 47354 9332 47356
rect 9356 47354 9412 47356
rect 9116 47302 9162 47354
rect 9162 47302 9172 47354
rect 9196 47302 9226 47354
rect 9226 47302 9238 47354
rect 9238 47302 9252 47354
rect 9276 47302 9290 47354
rect 9290 47302 9302 47354
rect 9302 47302 9332 47354
rect 9356 47302 9366 47354
rect 9366 47302 9412 47354
rect 9116 47300 9172 47302
rect 9196 47300 9252 47302
rect 9276 47300 9332 47302
rect 9356 47300 9412 47302
rect 7484 46810 7540 46812
rect 7564 46810 7620 46812
rect 7644 46810 7700 46812
rect 7724 46810 7780 46812
rect 7484 46758 7530 46810
rect 7530 46758 7540 46810
rect 7564 46758 7594 46810
rect 7594 46758 7606 46810
rect 7606 46758 7620 46810
rect 7644 46758 7658 46810
rect 7658 46758 7670 46810
rect 7670 46758 7700 46810
rect 7724 46758 7734 46810
rect 7734 46758 7780 46810
rect 7484 46756 7540 46758
rect 7564 46756 7620 46758
rect 7644 46756 7700 46758
rect 7724 46756 7780 46758
rect 9116 46266 9172 46268
rect 9196 46266 9252 46268
rect 9276 46266 9332 46268
rect 9356 46266 9412 46268
rect 9116 46214 9162 46266
rect 9162 46214 9172 46266
rect 9196 46214 9226 46266
rect 9226 46214 9238 46266
rect 9238 46214 9252 46266
rect 9276 46214 9290 46266
rect 9290 46214 9302 46266
rect 9302 46214 9332 46266
rect 9356 46214 9366 46266
rect 9366 46214 9412 46266
rect 9116 46212 9172 46214
rect 9196 46212 9252 46214
rect 9276 46212 9332 46214
rect 9356 46212 9412 46214
rect 7484 45722 7540 45724
rect 7564 45722 7620 45724
rect 7644 45722 7700 45724
rect 7724 45722 7780 45724
rect 7484 45670 7530 45722
rect 7530 45670 7540 45722
rect 7564 45670 7594 45722
rect 7594 45670 7606 45722
rect 7606 45670 7620 45722
rect 7644 45670 7658 45722
rect 7658 45670 7670 45722
rect 7670 45670 7700 45722
rect 7724 45670 7734 45722
rect 7734 45670 7780 45722
rect 7484 45668 7540 45670
rect 7564 45668 7620 45670
rect 7644 45668 7700 45670
rect 7724 45668 7780 45670
rect 9116 45178 9172 45180
rect 9196 45178 9252 45180
rect 9276 45178 9332 45180
rect 9356 45178 9412 45180
rect 9116 45126 9162 45178
rect 9162 45126 9172 45178
rect 9196 45126 9226 45178
rect 9226 45126 9238 45178
rect 9238 45126 9252 45178
rect 9276 45126 9290 45178
rect 9290 45126 9302 45178
rect 9302 45126 9332 45178
rect 9356 45126 9366 45178
rect 9366 45126 9412 45178
rect 9116 45124 9172 45126
rect 9196 45124 9252 45126
rect 9276 45124 9332 45126
rect 9356 45124 9412 45126
rect 7484 44634 7540 44636
rect 7564 44634 7620 44636
rect 7644 44634 7700 44636
rect 7724 44634 7780 44636
rect 7484 44582 7530 44634
rect 7530 44582 7540 44634
rect 7564 44582 7594 44634
rect 7594 44582 7606 44634
rect 7606 44582 7620 44634
rect 7644 44582 7658 44634
rect 7658 44582 7670 44634
rect 7670 44582 7700 44634
rect 7724 44582 7734 44634
rect 7734 44582 7780 44634
rect 7484 44580 7540 44582
rect 7564 44580 7620 44582
rect 7644 44580 7700 44582
rect 7724 44580 7780 44582
rect 7484 43546 7540 43548
rect 7564 43546 7620 43548
rect 7644 43546 7700 43548
rect 7724 43546 7780 43548
rect 7484 43494 7530 43546
rect 7530 43494 7540 43546
rect 7564 43494 7594 43546
rect 7594 43494 7606 43546
rect 7606 43494 7620 43546
rect 7644 43494 7658 43546
rect 7658 43494 7670 43546
rect 7670 43494 7700 43546
rect 7724 43494 7734 43546
rect 7734 43494 7780 43546
rect 7484 43492 7540 43494
rect 7564 43492 7620 43494
rect 7644 43492 7700 43494
rect 7724 43492 7780 43494
rect 7484 42458 7540 42460
rect 7564 42458 7620 42460
rect 7644 42458 7700 42460
rect 7724 42458 7780 42460
rect 7484 42406 7530 42458
rect 7530 42406 7540 42458
rect 7564 42406 7594 42458
rect 7594 42406 7606 42458
rect 7606 42406 7620 42458
rect 7644 42406 7658 42458
rect 7658 42406 7670 42458
rect 7670 42406 7700 42458
rect 7724 42406 7734 42458
rect 7734 42406 7780 42458
rect 7484 42404 7540 42406
rect 7564 42404 7620 42406
rect 7644 42404 7700 42406
rect 7724 42404 7780 42406
rect 9116 44090 9172 44092
rect 9196 44090 9252 44092
rect 9276 44090 9332 44092
rect 9356 44090 9412 44092
rect 9116 44038 9162 44090
rect 9162 44038 9172 44090
rect 9196 44038 9226 44090
rect 9226 44038 9238 44090
rect 9238 44038 9252 44090
rect 9276 44038 9290 44090
rect 9290 44038 9302 44090
rect 9302 44038 9332 44090
rect 9356 44038 9366 44090
rect 9366 44038 9412 44090
rect 9116 44036 9172 44038
rect 9196 44036 9252 44038
rect 9276 44036 9332 44038
rect 9356 44036 9412 44038
rect 10138 76372 10140 76392
rect 10140 76372 10192 76392
rect 10192 76372 10194 76392
rect 10138 76336 10194 76372
rect 10138 75656 10194 75712
rect 10138 74840 10194 74896
rect 10138 74024 10194 74080
rect 10138 73344 10194 73400
rect 10138 72528 10194 72584
rect 10138 71712 10194 71768
rect 10138 71032 10194 71088
rect 10138 70216 10194 70272
rect 10138 69400 10194 69456
rect 10138 68756 10140 68776
rect 10140 68756 10192 68776
rect 10192 68756 10194 68776
rect 10138 68720 10194 68756
rect 10138 67904 10194 67960
rect 10138 67088 10194 67144
rect 10138 66408 10194 66464
rect 10138 65592 10194 65648
rect 10138 64776 10194 64832
rect 10138 64096 10194 64152
rect 10138 63316 10140 63336
rect 10140 63316 10192 63336
rect 10192 63316 10194 63336
rect 10138 63280 10194 63316
rect 10138 62464 10194 62520
rect 10138 61784 10194 61840
rect 10138 60968 10194 61024
rect 10138 60288 10194 60344
rect 10138 59472 10194 59528
rect 10138 58656 10194 58712
rect 10138 55664 10194 55720
rect 10046 54052 10102 54088
rect 10046 54032 10048 54052
rect 10048 54032 10100 54052
rect 10100 54032 10102 54052
rect 10046 53388 10048 53408
rect 10048 53388 10100 53408
rect 10100 53388 10102 53408
rect 10046 53352 10102 53388
rect 10046 52536 10102 52592
rect 10046 51756 10048 51776
rect 10048 51756 10100 51776
rect 10100 51756 10102 51776
rect 10046 51720 10102 51756
rect 10046 51040 10102 51096
rect 10046 50224 10102 50280
rect 10046 48728 10102 48784
rect 10046 47948 10048 47968
rect 10048 47948 10100 47968
rect 10100 47948 10102 47968
rect 10046 47912 10102 47948
rect 10046 47096 10102 47152
rect 10046 46436 10102 46472
rect 10046 46416 10048 46436
rect 10048 46416 10100 46436
rect 10100 46416 10102 46436
rect 9116 43002 9172 43004
rect 9196 43002 9252 43004
rect 9276 43002 9332 43004
rect 9356 43002 9412 43004
rect 9116 42950 9162 43002
rect 9162 42950 9172 43002
rect 9196 42950 9226 43002
rect 9226 42950 9238 43002
rect 9238 42950 9252 43002
rect 9276 42950 9290 43002
rect 9290 42950 9302 43002
rect 9302 42950 9332 43002
rect 9356 42950 9366 43002
rect 9366 42950 9412 43002
rect 9116 42948 9172 42950
rect 9196 42948 9252 42950
rect 9276 42948 9332 42950
rect 9356 42948 9412 42950
rect 9116 41914 9172 41916
rect 9196 41914 9252 41916
rect 9276 41914 9332 41916
rect 9356 41914 9412 41916
rect 9116 41862 9162 41914
rect 9162 41862 9172 41914
rect 9196 41862 9226 41914
rect 9226 41862 9238 41914
rect 9238 41862 9252 41914
rect 9276 41862 9290 41914
rect 9290 41862 9302 41914
rect 9302 41862 9332 41914
rect 9356 41862 9366 41914
rect 9366 41862 9412 41914
rect 9116 41860 9172 41862
rect 9196 41860 9252 41862
rect 9276 41860 9332 41862
rect 9356 41860 9412 41862
rect 7484 41370 7540 41372
rect 7564 41370 7620 41372
rect 7644 41370 7700 41372
rect 7724 41370 7780 41372
rect 7484 41318 7530 41370
rect 7530 41318 7540 41370
rect 7564 41318 7594 41370
rect 7594 41318 7606 41370
rect 7606 41318 7620 41370
rect 7644 41318 7658 41370
rect 7658 41318 7670 41370
rect 7670 41318 7700 41370
rect 7724 41318 7734 41370
rect 7734 41318 7780 41370
rect 7484 41316 7540 41318
rect 7564 41316 7620 41318
rect 7644 41316 7700 41318
rect 7724 41316 7780 41318
rect 9116 40826 9172 40828
rect 9196 40826 9252 40828
rect 9276 40826 9332 40828
rect 9356 40826 9412 40828
rect 9116 40774 9162 40826
rect 9162 40774 9172 40826
rect 9196 40774 9226 40826
rect 9226 40774 9238 40826
rect 9238 40774 9252 40826
rect 9276 40774 9290 40826
rect 9290 40774 9302 40826
rect 9302 40774 9332 40826
rect 9356 40774 9366 40826
rect 9366 40774 9412 40826
rect 9116 40772 9172 40774
rect 9196 40772 9252 40774
rect 9276 40772 9332 40774
rect 9356 40772 9412 40774
rect 7484 40282 7540 40284
rect 7564 40282 7620 40284
rect 7644 40282 7700 40284
rect 7724 40282 7780 40284
rect 7484 40230 7530 40282
rect 7530 40230 7540 40282
rect 7564 40230 7594 40282
rect 7594 40230 7606 40282
rect 7606 40230 7620 40282
rect 7644 40230 7658 40282
rect 7658 40230 7670 40282
rect 7670 40230 7700 40282
rect 7724 40230 7734 40282
rect 7734 40230 7780 40282
rect 7484 40228 7540 40230
rect 7564 40228 7620 40230
rect 7644 40228 7700 40230
rect 7724 40228 7780 40230
rect 9116 39738 9172 39740
rect 9196 39738 9252 39740
rect 9276 39738 9332 39740
rect 9356 39738 9412 39740
rect 9116 39686 9162 39738
rect 9162 39686 9172 39738
rect 9196 39686 9226 39738
rect 9226 39686 9238 39738
rect 9238 39686 9252 39738
rect 9276 39686 9290 39738
rect 9290 39686 9302 39738
rect 9302 39686 9332 39738
rect 9356 39686 9366 39738
rect 9366 39686 9412 39738
rect 9116 39684 9172 39686
rect 9196 39684 9252 39686
rect 9276 39684 9332 39686
rect 9356 39684 9412 39686
rect 10046 45600 10102 45656
rect 10046 44784 10102 44840
rect 10046 44140 10048 44160
rect 10048 44140 10100 44160
rect 10100 44140 10102 44160
rect 10046 44104 10102 44140
rect 10046 43288 10102 43344
rect 10046 42508 10048 42528
rect 10048 42508 10100 42528
rect 10100 42508 10102 42528
rect 10046 42472 10102 42508
rect 10046 41792 10102 41848
rect 10046 40996 10102 41032
rect 10046 40976 10048 40996
rect 10048 40976 10100 40996
rect 10100 40976 10102 40996
rect 10046 40332 10048 40352
rect 10048 40332 10100 40352
rect 10100 40332 10102 40352
rect 10046 40296 10102 40332
rect 7484 39194 7540 39196
rect 7564 39194 7620 39196
rect 7644 39194 7700 39196
rect 7724 39194 7780 39196
rect 7484 39142 7530 39194
rect 7530 39142 7540 39194
rect 7564 39142 7594 39194
rect 7594 39142 7606 39194
rect 7606 39142 7620 39194
rect 7644 39142 7658 39194
rect 7658 39142 7670 39194
rect 7670 39142 7700 39194
rect 7724 39142 7734 39194
rect 7734 39142 7780 39194
rect 7484 39140 7540 39142
rect 7564 39140 7620 39142
rect 7644 39140 7700 39142
rect 7724 39140 7780 39142
rect 9116 38650 9172 38652
rect 9196 38650 9252 38652
rect 9276 38650 9332 38652
rect 9356 38650 9412 38652
rect 9116 38598 9162 38650
rect 9162 38598 9172 38650
rect 9196 38598 9226 38650
rect 9226 38598 9238 38650
rect 9238 38598 9252 38650
rect 9276 38598 9290 38650
rect 9290 38598 9302 38650
rect 9302 38598 9332 38650
rect 9356 38598 9366 38650
rect 9366 38598 9412 38650
rect 9116 38596 9172 38598
rect 9196 38596 9252 38598
rect 9276 38596 9332 38598
rect 9356 38596 9412 38598
rect 7484 38106 7540 38108
rect 7564 38106 7620 38108
rect 7644 38106 7700 38108
rect 7724 38106 7780 38108
rect 7484 38054 7530 38106
rect 7530 38054 7540 38106
rect 7564 38054 7594 38106
rect 7594 38054 7606 38106
rect 7606 38054 7620 38106
rect 7644 38054 7658 38106
rect 7658 38054 7670 38106
rect 7670 38054 7700 38106
rect 7724 38054 7734 38106
rect 7734 38054 7780 38106
rect 7484 38052 7540 38054
rect 7564 38052 7620 38054
rect 7644 38052 7700 38054
rect 7724 38052 7780 38054
rect 9116 37562 9172 37564
rect 9196 37562 9252 37564
rect 9276 37562 9332 37564
rect 9356 37562 9412 37564
rect 9116 37510 9162 37562
rect 9162 37510 9172 37562
rect 9196 37510 9226 37562
rect 9226 37510 9238 37562
rect 9238 37510 9252 37562
rect 9276 37510 9290 37562
rect 9290 37510 9302 37562
rect 9302 37510 9332 37562
rect 9356 37510 9366 37562
rect 9366 37510 9412 37562
rect 9116 37508 9172 37510
rect 9196 37508 9252 37510
rect 9276 37508 9332 37510
rect 9356 37508 9412 37510
rect 7484 37018 7540 37020
rect 7564 37018 7620 37020
rect 7644 37018 7700 37020
rect 7724 37018 7780 37020
rect 7484 36966 7530 37018
rect 7530 36966 7540 37018
rect 7564 36966 7594 37018
rect 7594 36966 7606 37018
rect 7606 36966 7620 37018
rect 7644 36966 7658 37018
rect 7658 36966 7670 37018
rect 7670 36966 7700 37018
rect 7724 36966 7734 37018
rect 7734 36966 7780 37018
rect 7484 36964 7540 36966
rect 7564 36964 7620 36966
rect 7644 36964 7700 36966
rect 7724 36964 7780 36966
rect 9116 36474 9172 36476
rect 9196 36474 9252 36476
rect 9276 36474 9332 36476
rect 9356 36474 9412 36476
rect 9116 36422 9162 36474
rect 9162 36422 9172 36474
rect 9196 36422 9226 36474
rect 9226 36422 9238 36474
rect 9238 36422 9252 36474
rect 9276 36422 9290 36474
rect 9290 36422 9302 36474
rect 9302 36422 9332 36474
rect 9356 36422 9366 36474
rect 9366 36422 9412 36474
rect 9116 36420 9172 36422
rect 9196 36420 9252 36422
rect 9276 36420 9332 36422
rect 9356 36420 9412 36422
rect 10046 39480 10102 39536
rect 10046 38700 10048 38720
rect 10048 38700 10100 38720
rect 10100 38700 10102 38720
rect 10046 38664 10102 38700
rect 7484 35930 7540 35932
rect 7564 35930 7620 35932
rect 7644 35930 7700 35932
rect 7724 35930 7780 35932
rect 7484 35878 7530 35930
rect 7530 35878 7540 35930
rect 7564 35878 7594 35930
rect 7594 35878 7606 35930
rect 7606 35878 7620 35930
rect 7644 35878 7658 35930
rect 7658 35878 7670 35930
rect 7670 35878 7700 35930
rect 7724 35878 7734 35930
rect 7734 35878 7780 35930
rect 7484 35876 7540 35878
rect 7564 35876 7620 35878
rect 7644 35876 7700 35878
rect 7724 35876 7780 35878
rect 9116 35386 9172 35388
rect 9196 35386 9252 35388
rect 9276 35386 9332 35388
rect 9356 35386 9412 35388
rect 9116 35334 9162 35386
rect 9162 35334 9172 35386
rect 9196 35334 9226 35386
rect 9226 35334 9238 35386
rect 9238 35334 9252 35386
rect 9276 35334 9290 35386
rect 9290 35334 9302 35386
rect 9302 35334 9332 35386
rect 9356 35334 9366 35386
rect 9366 35334 9412 35386
rect 9116 35332 9172 35334
rect 9196 35332 9252 35334
rect 9276 35332 9332 35334
rect 9356 35332 9412 35334
rect 7484 34842 7540 34844
rect 7564 34842 7620 34844
rect 7644 34842 7700 34844
rect 7724 34842 7780 34844
rect 7484 34790 7530 34842
rect 7530 34790 7540 34842
rect 7564 34790 7594 34842
rect 7594 34790 7606 34842
rect 7606 34790 7620 34842
rect 7644 34790 7658 34842
rect 7658 34790 7670 34842
rect 7670 34790 7700 34842
rect 7724 34790 7734 34842
rect 7734 34790 7780 34842
rect 7484 34788 7540 34790
rect 7564 34788 7620 34790
rect 7644 34788 7700 34790
rect 7724 34788 7780 34790
rect 9116 34298 9172 34300
rect 9196 34298 9252 34300
rect 9276 34298 9332 34300
rect 9356 34298 9412 34300
rect 9116 34246 9162 34298
rect 9162 34246 9172 34298
rect 9196 34246 9226 34298
rect 9226 34246 9238 34298
rect 9238 34246 9252 34298
rect 9276 34246 9290 34298
rect 9290 34246 9302 34298
rect 9302 34246 9332 34298
rect 9356 34246 9366 34298
rect 9366 34246 9412 34298
rect 9116 34244 9172 34246
rect 9196 34244 9252 34246
rect 9276 34244 9332 34246
rect 9356 34244 9412 34246
rect 9586 34040 9642 34096
rect 7484 33754 7540 33756
rect 7564 33754 7620 33756
rect 7644 33754 7700 33756
rect 7724 33754 7780 33756
rect 7484 33702 7530 33754
rect 7530 33702 7540 33754
rect 7564 33702 7594 33754
rect 7594 33702 7606 33754
rect 7606 33702 7620 33754
rect 7644 33702 7658 33754
rect 7658 33702 7670 33754
rect 7670 33702 7700 33754
rect 7724 33702 7734 33754
rect 7734 33702 7780 33754
rect 7484 33700 7540 33702
rect 7564 33700 7620 33702
rect 7644 33700 7700 33702
rect 7724 33700 7780 33702
rect 9116 33210 9172 33212
rect 9196 33210 9252 33212
rect 9276 33210 9332 33212
rect 9356 33210 9412 33212
rect 9116 33158 9162 33210
rect 9162 33158 9172 33210
rect 9196 33158 9226 33210
rect 9226 33158 9238 33210
rect 9238 33158 9252 33210
rect 9276 33158 9290 33210
rect 9290 33158 9302 33210
rect 9302 33158 9332 33210
rect 9356 33158 9366 33210
rect 9366 33158 9412 33210
rect 9116 33156 9172 33158
rect 9196 33156 9252 33158
rect 9276 33156 9332 33158
rect 9356 33156 9412 33158
rect 7484 32666 7540 32668
rect 7564 32666 7620 32668
rect 7644 32666 7700 32668
rect 7724 32666 7780 32668
rect 7484 32614 7530 32666
rect 7530 32614 7540 32666
rect 7564 32614 7594 32666
rect 7594 32614 7606 32666
rect 7606 32614 7620 32666
rect 7644 32614 7658 32666
rect 7658 32614 7670 32666
rect 7670 32614 7700 32666
rect 7724 32614 7734 32666
rect 7734 32614 7780 32666
rect 7484 32612 7540 32614
rect 7564 32612 7620 32614
rect 7644 32612 7700 32614
rect 7724 32612 7780 32614
rect 9116 32122 9172 32124
rect 9196 32122 9252 32124
rect 9276 32122 9332 32124
rect 9356 32122 9412 32124
rect 9116 32070 9162 32122
rect 9162 32070 9172 32122
rect 9196 32070 9226 32122
rect 9226 32070 9238 32122
rect 9238 32070 9252 32122
rect 9276 32070 9290 32122
rect 9290 32070 9302 32122
rect 9302 32070 9332 32122
rect 9356 32070 9366 32122
rect 9366 32070 9412 32122
rect 9116 32068 9172 32070
rect 9196 32068 9252 32070
rect 9276 32068 9332 32070
rect 9356 32068 9412 32070
rect 10046 37984 10102 38040
rect 10046 37168 10102 37224
rect 10046 36352 10102 36408
rect 10046 35672 10102 35728
rect 10046 34892 10048 34912
rect 10048 34892 10100 34912
rect 10100 34892 10102 34912
rect 10046 34856 10102 34892
rect 10046 33380 10102 33416
rect 10046 33360 10048 33380
rect 10048 33360 10100 33380
rect 10100 33360 10102 33380
rect 10046 32544 10102 32600
rect 10046 31728 10102 31784
rect 7484 31578 7540 31580
rect 7564 31578 7620 31580
rect 7644 31578 7700 31580
rect 7724 31578 7780 31580
rect 7484 31526 7530 31578
rect 7530 31526 7540 31578
rect 7564 31526 7594 31578
rect 7594 31526 7606 31578
rect 7606 31526 7620 31578
rect 7644 31526 7658 31578
rect 7658 31526 7670 31578
rect 7670 31526 7700 31578
rect 7724 31526 7734 31578
rect 7734 31526 7780 31578
rect 7484 31524 7540 31526
rect 7564 31524 7620 31526
rect 7644 31524 7700 31526
rect 7724 31524 7780 31526
rect 9116 31034 9172 31036
rect 9196 31034 9252 31036
rect 9276 31034 9332 31036
rect 9356 31034 9412 31036
rect 9116 30982 9162 31034
rect 9162 30982 9172 31034
rect 9196 30982 9226 31034
rect 9226 30982 9238 31034
rect 9238 30982 9252 31034
rect 9276 30982 9290 31034
rect 9290 30982 9302 31034
rect 9302 30982 9332 31034
rect 9356 30982 9366 31034
rect 9366 30982 9412 31034
rect 9116 30980 9172 30982
rect 9196 30980 9252 30982
rect 9276 30980 9332 30982
rect 9356 30980 9412 30982
rect 7484 30490 7540 30492
rect 7564 30490 7620 30492
rect 7644 30490 7700 30492
rect 7724 30490 7780 30492
rect 7484 30438 7530 30490
rect 7530 30438 7540 30490
rect 7564 30438 7594 30490
rect 7594 30438 7606 30490
rect 7606 30438 7620 30490
rect 7644 30438 7658 30490
rect 7658 30438 7670 30490
rect 7670 30438 7700 30490
rect 7724 30438 7734 30490
rect 7734 30438 7780 30490
rect 7484 30436 7540 30438
rect 7564 30436 7620 30438
rect 7644 30436 7700 30438
rect 7724 30436 7780 30438
rect 10046 31084 10048 31104
rect 10048 31084 10100 31104
rect 10100 31084 10102 31104
rect 10046 31048 10102 31084
rect 10046 30232 10102 30288
rect 9116 29946 9172 29948
rect 9196 29946 9252 29948
rect 9276 29946 9332 29948
rect 9356 29946 9412 29948
rect 9116 29894 9162 29946
rect 9162 29894 9172 29946
rect 9196 29894 9226 29946
rect 9226 29894 9238 29946
rect 9238 29894 9252 29946
rect 9276 29894 9290 29946
rect 9290 29894 9302 29946
rect 9302 29894 9332 29946
rect 9356 29894 9366 29946
rect 9366 29894 9412 29946
rect 9116 29892 9172 29894
rect 9196 29892 9252 29894
rect 9276 29892 9332 29894
rect 9356 29892 9412 29894
rect 7484 29402 7540 29404
rect 7564 29402 7620 29404
rect 7644 29402 7700 29404
rect 7724 29402 7780 29404
rect 7484 29350 7530 29402
rect 7530 29350 7540 29402
rect 7564 29350 7594 29402
rect 7594 29350 7606 29402
rect 7606 29350 7620 29402
rect 7644 29350 7658 29402
rect 7658 29350 7670 29402
rect 7670 29350 7700 29402
rect 7724 29350 7734 29402
rect 7734 29350 7780 29402
rect 7484 29348 7540 29350
rect 7564 29348 7620 29350
rect 7644 29348 7700 29350
rect 7724 29348 7780 29350
rect 7484 28314 7540 28316
rect 7564 28314 7620 28316
rect 7644 28314 7700 28316
rect 7724 28314 7780 28316
rect 7484 28262 7530 28314
rect 7530 28262 7540 28314
rect 7564 28262 7594 28314
rect 7594 28262 7606 28314
rect 7606 28262 7620 28314
rect 7644 28262 7658 28314
rect 7658 28262 7670 28314
rect 7670 28262 7700 28314
rect 7724 28262 7734 28314
rect 7734 28262 7780 28314
rect 7484 28260 7540 28262
rect 7564 28260 7620 28262
rect 7644 28260 7700 28262
rect 7724 28260 7780 28262
rect 7484 27226 7540 27228
rect 7564 27226 7620 27228
rect 7644 27226 7700 27228
rect 7724 27226 7780 27228
rect 7484 27174 7530 27226
rect 7530 27174 7540 27226
rect 7564 27174 7594 27226
rect 7594 27174 7606 27226
rect 7606 27174 7620 27226
rect 7644 27174 7658 27226
rect 7658 27174 7670 27226
rect 7670 27174 7700 27226
rect 7724 27174 7734 27226
rect 7734 27174 7780 27226
rect 7484 27172 7540 27174
rect 7564 27172 7620 27174
rect 7644 27172 7700 27174
rect 7724 27172 7780 27174
rect 7484 26138 7540 26140
rect 7564 26138 7620 26140
rect 7644 26138 7700 26140
rect 7724 26138 7780 26140
rect 7484 26086 7530 26138
rect 7530 26086 7540 26138
rect 7564 26086 7594 26138
rect 7594 26086 7606 26138
rect 7606 26086 7620 26138
rect 7644 26086 7658 26138
rect 7658 26086 7670 26138
rect 7670 26086 7700 26138
rect 7724 26086 7734 26138
rect 7734 26086 7780 26138
rect 7484 26084 7540 26086
rect 7564 26084 7620 26086
rect 7644 26084 7700 26086
rect 7724 26084 7780 26086
rect 5852 25594 5908 25596
rect 5932 25594 5988 25596
rect 6012 25594 6068 25596
rect 6092 25594 6148 25596
rect 5852 25542 5898 25594
rect 5898 25542 5908 25594
rect 5932 25542 5962 25594
rect 5962 25542 5974 25594
rect 5974 25542 5988 25594
rect 6012 25542 6026 25594
rect 6026 25542 6038 25594
rect 6038 25542 6068 25594
rect 6092 25542 6102 25594
rect 6102 25542 6148 25594
rect 5852 25540 5908 25542
rect 5932 25540 5988 25542
rect 6012 25540 6068 25542
rect 6092 25540 6148 25542
rect 7484 25050 7540 25052
rect 7564 25050 7620 25052
rect 7644 25050 7700 25052
rect 7724 25050 7780 25052
rect 7484 24998 7530 25050
rect 7530 24998 7540 25050
rect 7564 24998 7594 25050
rect 7594 24998 7606 25050
rect 7606 24998 7620 25050
rect 7644 24998 7658 25050
rect 7658 24998 7670 25050
rect 7670 24998 7700 25050
rect 7724 24998 7734 25050
rect 7734 24998 7780 25050
rect 7484 24996 7540 24998
rect 7564 24996 7620 24998
rect 7644 24996 7700 24998
rect 7724 24996 7780 24998
rect 5852 24506 5908 24508
rect 5932 24506 5988 24508
rect 6012 24506 6068 24508
rect 6092 24506 6148 24508
rect 5852 24454 5898 24506
rect 5898 24454 5908 24506
rect 5932 24454 5962 24506
rect 5962 24454 5974 24506
rect 5974 24454 5988 24506
rect 6012 24454 6026 24506
rect 6026 24454 6038 24506
rect 6038 24454 6068 24506
rect 6092 24454 6102 24506
rect 6102 24454 6148 24506
rect 5852 24452 5908 24454
rect 5932 24452 5988 24454
rect 6012 24452 6068 24454
rect 6092 24452 6148 24454
rect 7484 23962 7540 23964
rect 7564 23962 7620 23964
rect 7644 23962 7700 23964
rect 7724 23962 7780 23964
rect 7484 23910 7530 23962
rect 7530 23910 7540 23962
rect 7564 23910 7594 23962
rect 7594 23910 7606 23962
rect 7606 23910 7620 23962
rect 7644 23910 7658 23962
rect 7658 23910 7670 23962
rect 7670 23910 7700 23962
rect 7724 23910 7734 23962
rect 7734 23910 7780 23962
rect 7484 23908 7540 23910
rect 7564 23908 7620 23910
rect 7644 23908 7700 23910
rect 7724 23908 7780 23910
rect 5852 23418 5908 23420
rect 5932 23418 5988 23420
rect 6012 23418 6068 23420
rect 6092 23418 6148 23420
rect 5852 23366 5898 23418
rect 5898 23366 5908 23418
rect 5932 23366 5962 23418
rect 5962 23366 5974 23418
rect 5974 23366 5988 23418
rect 6012 23366 6026 23418
rect 6026 23366 6038 23418
rect 6038 23366 6068 23418
rect 6092 23366 6102 23418
rect 6102 23366 6148 23418
rect 5852 23364 5908 23366
rect 5932 23364 5988 23366
rect 6012 23364 6068 23366
rect 6092 23364 6148 23366
rect 7484 22874 7540 22876
rect 7564 22874 7620 22876
rect 7644 22874 7700 22876
rect 7724 22874 7780 22876
rect 7484 22822 7530 22874
rect 7530 22822 7540 22874
rect 7564 22822 7594 22874
rect 7594 22822 7606 22874
rect 7606 22822 7620 22874
rect 7644 22822 7658 22874
rect 7658 22822 7670 22874
rect 7670 22822 7700 22874
rect 7724 22822 7734 22874
rect 7734 22822 7780 22874
rect 7484 22820 7540 22822
rect 7564 22820 7620 22822
rect 7644 22820 7700 22822
rect 7724 22820 7780 22822
rect 5852 22330 5908 22332
rect 5932 22330 5988 22332
rect 6012 22330 6068 22332
rect 6092 22330 6148 22332
rect 5852 22278 5898 22330
rect 5898 22278 5908 22330
rect 5932 22278 5962 22330
rect 5962 22278 5974 22330
rect 5974 22278 5988 22330
rect 6012 22278 6026 22330
rect 6026 22278 6038 22330
rect 6038 22278 6068 22330
rect 6092 22278 6102 22330
rect 6102 22278 6148 22330
rect 5852 22276 5908 22278
rect 5932 22276 5988 22278
rect 6012 22276 6068 22278
rect 6092 22276 6148 22278
rect 7484 21786 7540 21788
rect 7564 21786 7620 21788
rect 7644 21786 7700 21788
rect 7724 21786 7780 21788
rect 7484 21734 7530 21786
rect 7530 21734 7540 21786
rect 7564 21734 7594 21786
rect 7594 21734 7606 21786
rect 7606 21734 7620 21786
rect 7644 21734 7658 21786
rect 7658 21734 7670 21786
rect 7670 21734 7700 21786
rect 7724 21734 7734 21786
rect 7734 21734 7780 21786
rect 7484 21732 7540 21734
rect 7564 21732 7620 21734
rect 7644 21732 7700 21734
rect 7724 21732 7780 21734
rect 5852 21242 5908 21244
rect 5932 21242 5988 21244
rect 6012 21242 6068 21244
rect 6092 21242 6148 21244
rect 5852 21190 5898 21242
rect 5898 21190 5908 21242
rect 5932 21190 5962 21242
rect 5962 21190 5974 21242
rect 5974 21190 5988 21242
rect 6012 21190 6026 21242
rect 6026 21190 6038 21242
rect 6038 21190 6068 21242
rect 6092 21190 6102 21242
rect 6102 21190 6148 21242
rect 5852 21188 5908 21190
rect 5932 21188 5988 21190
rect 6012 21188 6068 21190
rect 6092 21188 6148 21190
rect 7484 20698 7540 20700
rect 7564 20698 7620 20700
rect 7644 20698 7700 20700
rect 7724 20698 7780 20700
rect 7484 20646 7530 20698
rect 7530 20646 7540 20698
rect 7564 20646 7594 20698
rect 7594 20646 7606 20698
rect 7606 20646 7620 20698
rect 7644 20646 7658 20698
rect 7658 20646 7670 20698
rect 7670 20646 7700 20698
rect 7724 20646 7734 20698
rect 7734 20646 7780 20698
rect 7484 20644 7540 20646
rect 7564 20644 7620 20646
rect 7644 20644 7700 20646
rect 7724 20644 7780 20646
rect 10138 29416 10194 29472
rect 9116 28858 9172 28860
rect 9196 28858 9252 28860
rect 9276 28858 9332 28860
rect 9356 28858 9412 28860
rect 9116 28806 9162 28858
rect 9162 28806 9172 28858
rect 9196 28806 9226 28858
rect 9226 28806 9238 28858
rect 9238 28806 9252 28858
rect 9276 28806 9290 28858
rect 9290 28806 9302 28858
rect 9302 28806 9332 28858
rect 9356 28806 9366 28858
rect 9366 28806 9412 28858
rect 9116 28804 9172 28806
rect 9196 28804 9252 28806
rect 9276 28804 9332 28806
rect 9356 28804 9412 28806
rect 10138 28736 10194 28792
rect 9954 27956 9956 27976
rect 9956 27956 10008 27976
rect 10008 27956 10010 27976
rect 9954 27920 10010 27956
rect 9116 27770 9172 27772
rect 9196 27770 9252 27772
rect 9276 27770 9332 27772
rect 9356 27770 9412 27772
rect 9116 27718 9162 27770
rect 9162 27718 9172 27770
rect 9196 27718 9226 27770
rect 9226 27718 9238 27770
rect 9238 27718 9252 27770
rect 9276 27718 9290 27770
rect 9290 27718 9302 27770
rect 9302 27718 9332 27770
rect 9356 27718 9366 27770
rect 9366 27718 9412 27770
rect 9116 27716 9172 27718
rect 9196 27716 9252 27718
rect 9276 27716 9332 27718
rect 9356 27716 9412 27718
rect 9954 27104 10010 27160
rect 9116 26682 9172 26684
rect 9196 26682 9252 26684
rect 9276 26682 9332 26684
rect 9356 26682 9412 26684
rect 9116 26630 9162 26682
rect 9162 26630 9172 26682
rect 9196 26630 9226 26682
rect 9226 26630 9238 26682
rect 9238 26630 9252 26682
rect 9276 26630 9290 26682
rect 9290 26630 9302 26682
rect 9302 26630 9332 26682
rect 9356 26630 9366 26682
rect 9366 26630 9412 26682
rect 9116 26628 9172 26630
rect 9196 26628 9252 26630
rect 9276 26628 9332 26630
rect 9356 26628 9412 26630
rect 10138 26424 10194 26480
rect 10138 25644 10140 25664
rect 10140 25644 10192 25664
rect 10192 25644 10194 25664
rect 10138 25608 10194 25644
rect 9116 25594 9172 25596
rect 9196 25594 9252 25596
rect 9276 25594 9332 25596
rect 9356 25594 9412 25596
rect 9116 25542 9162 25594
rect 9162 25542 9172 25594
rect 9196 25542 9226 25594
rect 9226 25542 9238 25594
rect 9238 25542 9252 25594
rect 9276 25542 9290 25594
rect 9290 25542 9302 25594
rect 9302 25542 9332 25594
rect 9356 25542 9366 25594
rect 9366 25542 9412 25594
rect 9116 25540 9172 25542
rect 9196 25540 9252 25542
rect 9276 25540 9332 25542
rect 9356 25540 9412 25542
rect 10138 24792 10194 24848
rect 9116 24506 9172 24508
rect 9196 24506 9252 24508
rect 9276 24506 9332 24508
rect 9356 24506 9412 24508
rect 9116 24454 9162 24506
rect 9162 24454 9172 24506
rect 9196 24454 9226 24506
rect 9226 24454 9238 24506
rect 9238 24454 9252 24506
rect 9276 24454 9290 24506
rect 9290 24454 9302 24506
rect 9302 24454 9332 24506
rect 9356 24454 9366 24506
rect 9366 24454 9412 24506
rect 9116 24452 9172 24454
rect 9196 24452 9252 24454
rect 9276 24452 9332 24454
rect 9356 24452 9412 24454
rect 10138 24148 10140 24168
rect 10140 24148 10192 24168
rect 10192 24148 10194 24168
rect 10138 24112 10194 24148
rect 9116 23418 9172 23420
rect 9196 23418 9252 23420
rect 9276 23418 9332 23420
rect 9356 23418 9412 23420
rect 9116 23366 9162 23418
rect 9162 23366 9172 23418
rect 9196 23366 9226 23418
rect 9226 23366 9238 23418
rect 9238 23366 9252 23418
rect 9276 23366 9290 23418
rect 9290 23366 9302 23418
rect 9302 23366 9332 23418
rect 9356 23366 9366 23418
rect 9366 23366 9412 23418
rect 9116 23364 9172 23366
rect 9196 23364 9252 23366
rect 9276 23364 9332 23366
rect 9356 23364 9412 23366
rect 10138 23296 10194 23352
rect 10138 22500 10194 22536
rect 10138 22480 10140 22500
rect 10140 22480 10192 22500
rect 10192 22480 10194 22500
rect 9116 22330 9172 22332
rect 9196 22330 9252 22332
rect 9276 22330 9332 22332
rect 9356 22330 9412 22332
rect 9116 22278 9162 22330
rect 9162 22278 9172 22330
rect 9196 22278 9226 22330
rect 9226 22278 9238 22330
rect 9238 22278 9252 22330
rect 9276 22278 9290 22330
rect 9290 22278 9302 22330
rect 9302 22278 9332 22330
rect 9356 22278 9366 22330
rect 9366 22278 9412 22330
rect 9116 22276 9172 22278
rect 9196 22276 9252 22278
rect 9276 22276 9332 22278
rect 9356 22276 9412 22278
rect 10138 21800 10194 21856
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 9276 21242 9332 21244
rect 9356 21242 9412 21244
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9238 21242
rect 9238 21190 9252 21242
rect 9276 21190 9290 21242
rect 9290 21190 9302 21242
rect 9302 21190 9332 21242
rect 9356 21190 9366 21242
rect 9366 21190 9412 21242
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 9276 21188 9332 21190
rect 9356 21188 9412 21190
rect 10138 20984 10194 21040
rect 5852 20154 5908 20156
rect 5932 20154 5988 20156
rect 6012 20154 6068 20156
rect 6092 20154 6148 20156
rect 5852 20102 5898 20154
rect 5898 20102 5908 20154
rect 5932 20102 5962 20154
rect 5962 20102 5974 20154
rect 5974 20102 5988 20154
rect 6012 20102 6026 20154
rect 6026 20102 6038 20154
rect 6038 20102 6068 20154
rect 6092 20102 6102 20154
rect 6102 20102 6148 20154
rect 5852 20100 5908 20102
rect 5932 20100 5988 20102
rect 6012 20100 6068 20102
rect 6092 20100 6148 20102
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 9276 20154 9332 20156
rect 9356 20154 9412 20156
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9238 20154
rect 9238 20102 9252 20154
rect 9276 20102 9290 20154
rect 9290 20102 9302 20154
rect 9302 20102 9332 20154
rect 9356 20102 9366 20154
rect 9366 20102 9412 20154
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 9276 20100 9332 20102
rect 9356 20100 9412 20102
rect 7484 19610 7540 19612
rect 7564 19610 7620 19612
rect 7644 19610 7700 19612
rect 7724 19610 7780 19612
rect 7484 19558 7530 19610
rect 7530 19558 7540 19610
rect 7564 19558 7594 19610
rect 7594 19558 7606 19610
rect 7606 19558 7620 19610
rect 7644 19558 7658 19610
rect 7658 19558 7670 19610
rect 7670 19558 7700 19610
rect 7724 19558 7734 19610
rect 7734 19558 7780 19610
rect 7484 19556 7540 19558
rect 7564 19556 7620 19558
rect 7644 19556 7700 19558
rect 7724 19556 7780 19558
rect 5852 19066 5908 19068
rect 5932 19066 5988 19068
rect 6012 19066 6068 19068
rect 6092 19066 6148 19068
rect 5852 19014 5898 19066
rect 5898 19014 5908 19066
rect 5932 19014 5962 19066
rect 5962 19014 5974 19066
rect 5974 19014 5988 19066
rect 6012 19014 6026 19066
rect 6026 19014 6038 19066
rect 6038 19014 6068 19066
rect 6092 19014 6102 19066
rect 6102 19014 6148 19066
rect 5852 19012 5908 19014
rect 5932 19012 5988 19014
rect 6012 19012 6068 19014
rect 6092 19012 6148 19014
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 9276 19066 9332 19068
rect 9356 19066 9412 19068
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9238 19066
rect 9238 19014 9252 19066
rect 9276 19014 9290 19066
rect 9290 19014 9302 19066
rect 9302 19014 9332 19066
rect 9356 19014 9366 19066
rect 9366 19014 9412 19066
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 9276 19012 9332 19014
rect 9356 19012 9412 19014
rect 7484 18522 7540 18524
rect 7564 18522 7620 18524
rect 7644 18522 7700 18524
rect 7724 18522 7780 18524
rect 7484 18470 7530 18522
rect 7530 18470 7540 18522
rect 7564 18470 7594 18522
rect 7594 18470 7606 18522
rect 7606 18470 7620 18522
rect 7644 18470 7658 18522
rect 7658 18470 7670 18522
rect 7670 18470 7700 18522
rect 7724 18470 7734 18522
rect 7734 18470 7780 18522
rect 7484 18468 7540 18470
rect 7564 18468 7620 18470
rect 7644 18468 7700 18470
rect 7724 18468 7780 18470
rect 5852 17978 5908 17980
rect 5932 17978 5988 17980
rect 6012 17978 6068 17980
rect 6092 17978 6148 17980
rect 5852 17926 5898 17978
rect 5898 17926 5908 17978
rect 5932 17926 5962 17978
rect 5962 17926 5974 17978
rect 5974 17926 5988 17978
rect 6012 17926 6026 17978
rect 6026 17926 6038 17978
rect 6038 17926 6068 17978
rect 6092 17926 6102 17978
rect 6102 17926 6148 17978
rect 5852 17924 5908 17926
rect 5932 17924 5988 17926
rect 6012 17924 6068 17926
rect 6092 17924 6148 17926
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 9276 17978 9332 17980
rect 9356 17978 9412 17980
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9238 17978
rect 9238 17926 9252 17978
rect 9276 17926 9290 17978
rect 9290 17926 9302 17978
rect 9302 17926 9332 17978
rect 9356 17926 9366 17978
rect 9366 17926 9412 17978
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 9276 17924 9332 17926
rect 9356 17924 9412 17926
rect 7484 17434 7540 17436
rect 7564 17434 7620 17436
rect 7644 17434 7700 17436
rect 7724 17434 7780 17436
rect 7484 17382 7530 17434
rect 7530 17382 7540 17434
rect 7564 17382 7594 17434
rect 7594 17382 7606 17434
rect 7606 17382 7620 17434
rect 7644 17382 7658 17434
rect 7658 17382 7670 17434
rect 7670 17382 7700 17434
rect 7724 17382 7734 17434
rect 7734 17382 7780 17434
rect 7484 17380 7540 17382
rect 7564 17380 7620 17382
rect 7644 17380 7700 17382
rect 7724 17380 7780 17382
rect 5852 16890 5908 16892
rect 5932 16890 5988 16892
rect 6012 16890 6068 16892
rect 6092 16890 6148 16892
rect 5852 16838 5898 16890
rect 5898 16838 5908 16890
rect 5932 16838 5962 16890
rect 5962 16838 5974 16890
rect 5974 16838 5988 16890
rect 6012 16838 6026 16890
rect 6026 16838 6038 16890
rect 6038 16838 6068 16890
rect 6092 16838 6102 16890
rect 6102 16838 6148 16890
rect 5852 16836 5908 16838
rect 5932 16836 5988 16838
rect 6012 16836 6068 16838
rect 6092 16836 6148 16838
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 9276 16890 9332 16892
rect 9356 16890 9412 16892
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9238 16890
rect 9238 16838 9252 16890
rect 9276 16838 9290 16890
rect 9290 16838 9302 16890
rect 9302 16838 9332 16890
rect 9356 16838 9366 16890
rect 9366 16838 9412 16890
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 9276 16836 9332 16838
rect 9356 16836 9412 16838
rect 7484 16346 7540 16348
rect 7564 16346 7620 16348
rect 7644 16346 7700 16348
rect 7724 16346 7780 16348
rect 7484 16294 7530 16346
rect 7530 16294 7540 16346
rect 7564 16294 7594 16346
rect 7594 16294 7606 16346
rect 7606 16294 7620 16346
rect 7644 16294 7658 16346
rect 7658 16294 7670 16346
rect 7670 16294 7700 16346
rect 7724 16294 7734 16346
rect 7734 16294 7780 16346
rect 7484 16292 7540 16294
rect 7564 16292 7620 16294
rect 7644 16292 7700 16294
rect 7724 16292 7780 16294
rect 5852 15802 5908 15804
rect 5932 15802 5988 15804
rect 6012 15802 6068 15804
rect 6092 15802 6148 15804
rect 5852 15750 5898 15802
rect 5898 15750 5908 15802
rect 5932 15750 5962 15802
rect 5962 15750 5974 15802
rect 5974 15750 5988 15802
rect 6012 15750 6026 15802
rect 6026 15750 6038 15802
rect 6038 15750 6068 15802
rect 6092 15750 6102 15802
rect 6102 15750 6148 15802
rect 5852 15748 5908 15750
rect 5932 15748 5988 15750
rect 6012 15748 6068 15750
rect 6092 15748 6148 15750
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 9276 15802 9332 15804
rect 9356 15802 9412 15804
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9238 15802
rect 9238 15750 9252 15802
rect 9276 15750 9290 15802
rect 9290 15750 9302 15802
rect 9302 15750 9332 15802
rect 9356 15750 9366 15802
rect 9366 15750 9412 15802
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 9276 15748 9332 15750
rect 9356 15748 9412 15750
rect 7484 15258 7540 15260
rect 7564 15258 7620 15260
rect 7644 15258 7700 15260
rect 7724 15258 7780 15260
rect 7484 15206 7530 15258
rect 7530 15206 7540 15258
rect 7564 15206 7594 15258
rect 7594 15206 7606 15258
rect 7606 15206 7620 15258
rect 7644 15206 7658 15258
rect 7658 15206 7670 15258
rect 7670 15206 7700 15258
rect 7724 15206 7734 15258
rect 7734 15206 7780 15258
rect 7484 15204 7540 15206
rect 7564 15204 7620 15206
rect 7644 15204 7700 15206
rect 7724 15204 7780 15206
rect 5852 14714 5908 14716
rect 5932 14714 5988 14716
rect 6012 14714 6068 14716
rect 6092 14714 6148 14716
rect 5852 14662 5898 14714
rect 5898 14662 5908 14714
rect 5932 14662 5962 14714
rect 5962 14662 5974 14714
rect 5974 14662 5988 14714
rect 6012 14662 6026 14714
rect 6026 14662 6038 14714
rect 6038 14662 6068 14714
rect 6092 14662 6102 14714
rect 6102 14662 6148 14714
rect 5852 14660 5908 14662
rect 5932 14660 5988 14662
rect 6012 14660 6068 14662
rect 6092 14660 6148 14662
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 9276 14714 9332 14716
rect 9356 14714 9412 14716
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9238 14714
rect 9238 14662 9252 14714
rect 9276 14662 9290 14714
rect 9290 14662 9302 14714
rect 9302 14662 9332 14714
rect 9356 14662 9366 14714
rect 9366 14662 9412 14714
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 9276 14660 9332 14662
rect 9356 14660 9412 14662
rect 7484 14170 7540 14172
rect 7564 14170 7620 14172
rect 7644 14170 7700 14172
rect 7724 14170 7780 14172
rect 7484 14118 7530 14170
rect 7530 14118 7540 14170
rect 7564 14118 7594 14170
rect 7594 14118 7606 14170
rect 7606 14118 7620 14170
rect 7644 14118 7658 14170
rect 7658 14118 7670 14170
rect 7670 14118 7700 14170
rect 7724 14118 7734 14170
rect 7734 14118 7780 14170
rect 7484 14116 7540 14118
rect 7564 14116 7620 14118
rect 7644 14116 7700 14118
rect 7724 14116 7780 14118
rect 5852 13626 5908 13628
rect 5932 13626 5988 13628
rect 6012 13626 6068 13628
rect 6092 13626 6148 13628
rect 5852 13574 5898 13626
rect 5898 13574 5908 13626
rect 5932 13574 5962 13626
rect 5962 13574 5974 13626
rect 5974 13574 5988 13626
rect 6012 13574 6026 13626
rect 6026 13574 6038 13626
rect 6038 13574 6068 13626
rect 6092 13574 6102 13626
rect 6102 13574 6148 13626
rect 5852 13572 5908 13574
rect 5932 13572 5988 13574
rect 6012 13572 6068 13574
rect 6092 13572 6148 13574
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 9276 13626 9332 13628
rect 9356 13626 9412 13628
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9238 13626
rect 9238 13574 9252 13626
rect 9276 13574 9290 13626
rect 9290 13574 9302 13626
rect 9302 13574 9332 13626
rect 9356 13574 9366 13626
rect 9366 13574 9412 13626
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 9276 13572 9332 13574
rect 9356 13572 9412 13574
rect 9586 13368 9642 13424
rect 7484 13082 7540 13084
rect 7564 13082 7620 13084
rect 7644 13082 7700 13084
rect 7724 13082 7780 13084
rect 7484 13030 7530 13082
rect 7530 13030 7540 13082
rect 7564 13030 7594 13082
rect 7594 13030 7606 13082
rect 7606 13030 7620 13082
rect 7644 13030 7658 13082
rect 7658 13030 7670 13082
rect 7670 13030 7700 13082
rect 7724 13030 7734 13082
rect 7734 13030 7780 13082
rect 7484 13028 7540 13030
rect 7564 13028 7620 13030
rect 7644 13028 7700 13030
rect 7724 13028 7780 13030
rect 10046 20324 10102 20360
rect 10046 20304 10048 20324
rect 10048 20304 10100 20324
rect 10100 20304 10102 20324
rect 10046 19488 10102 19544
rect 10046 18672 10102 18728
rect 10046 18028 10048 18048
rect 10048 18028 10100 18048
rect 10100 18028 10102 18048
rect 10046 17992 10102 18028
rect 10046 17176 10102 17232
rect 10046 16396 10048 16416
rect 10048 16396 10100 16416
rect 10100 16396 10102 16416
rect 10046 16360 10102 16396
rect 10046 15680 10102 15736
rect 5852 12538 5908 12540
rect 5932 12538 5988 12540
rect 6012 12538 6068 12540
rect 6092 12538 6148 12540
rect 5852 12486 5898 12538
rect 5898 12486 5908 12538
rect 5932 12486 5962 12538
rect 5962 12486 5974 12538
rect 5974 12486 5988 12538
rect 6012 12486 6026 12538
rect 6026 12486 6038 12538
rect 6038 12486 6068 12538
rect 6092 12486 6102 12538
rect 6102 12486 6148 12538
rect 5852 12484 5908 12486
rect 5932 12484 5988 12486
rect 6012 12484 6068 12486
rect 6092 12484 6148 12486
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 9276 12538 9332 12540
rect 9356 12538 9412 12540
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9238 12538
rect 9238 12486 9252 12538
rect 9276 12486 9290 12538
rect 9290 12486 9302 12538
rect 9302 12486 9332 12538
rect 9356 12486 9366 12538
rect 9366 12486 9412 12538
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 9276 12484 9332 12486
rect 9356 12484 9412 12486
rect 10046 14884 10102 14920
rect 10046 14864 10048 14884
rect 10048 14864 10100 14884
rect 10100 14864 10102 14884
rect 10046 14048 10102 14104
rect 10046 12588 10048 12608
rect 10048 12588 10100 12608
rect 10100 12588 10102 12608
rect 10046 12552 10102 12588
rect 7484 11994 7540 11996
rect 7564 11994 7620 11996
rect 7644 11994 7700 11996
rect 7724 11994 7780 11996
rect 7484 11942 7530 11994
rect 7530 11942 7540 11994
rect 7564 11942 7594 11994
rect 7594 11942 7606 11994
rect 7606 11942 7620 11994
rect 7644 11942 7658 11994
rect 7658 11942 7670 11994
rect 7670 11942 7700 11994
rect 7724 11942 7734 11994
rect 7734 11942 7780 11994
rect 7484 11940 7540 11942
rect 7564 11940 7620 11942
rect 7644 11940 7700 11942
rect 7724 11940 7780 11942
rect 10046 11736 10102 11792
rect 5852 11450 5908 11452
rect 5932 11450 5988 11452
rect 6012 11450 6068 11452
rect 6092 11450 6148 11452
rect 5852 11398 5898 11450
rect 5898 11398 5908 11450
rect 5932 11398 5962 11450
rect 5962 11398 5974 11450
rect 5974 11398 5988 11450
rect 6012 11398 6026 11450
rect 6026 11398 6038 11450
rect 6038 11398 6068 11450
rect 6092 11398 6102 11450
rect 6102 11398 6148 11450
rect 5852 11396 5908 11398
rect 5932 11396 5988 11398
rect 6012 11396 6068 11398
rect 6092 11396 6148 11398
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 9276 11450 9332 11452
rect 9356 11450 9412 11452
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9238 11450
rect 9238 11398 9252 11450
rect 9276 11398 9290 11450
rect 9290 11398 9302 11450
rect 9302 11398 9332 11450
rect 9356 11398 9366 11450
rect 9366 11398 9412 11450
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 9276 11396 9332 11398
rect 9356 11396 9412 11398
rect 10046 11056 10102 11112
rect 7484 10906 7540 10908
rect 7564 10906 7620 10908
rect 7644 10906 7700 10908
rect 7724 10906 7780 10908
rect 7484 10854 7530 10906
rect 7530 10854 7540 10906
rect 7564 10854 7594 10906
rect 7594 10854 7606 10906
rect 7606 10854 7620 10906
rect 7644 10854 7658 10906
rect 7658 10854 7670 10906
rect 7670 10854 7700 10906
rect 7724 10854 7734 10906
rect 7734 10854 7780 10906
rect 7484 10852 7540 10854
rect 7564 10852 7620 10854
rect 7644 10852 7700 10854
rect 7724 10852 7780 10854
rect 5852 10362 5908 10364
rect 5932 10362 5988 10364
rect 6012 10362 6068 10364
rect 6092 10362 6148 10364
rect 5852 10310 5898 10362
rect 5898 10310 5908 10362
rect 5932 10310 5962 10362
rect 5962 10310 5974 10362
rect 5974 10310 5988 10362
rect 6012 10310 6026 10362
rect 6026 10310 6038 10362
rect 6038 10310 6068 10362
rect 6092 10310 6102 10362
rect 6102 10310 6148 10362
rect 5852 10308 5908 10310
rect 5932 10308 5988 10310
rect 6012 10308 6068 10310
rect 6092 10308 6148 10310
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 9276 10362 9332 10364
rect 9356 10362 9412 10364
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9238 10362
rect 9238 10310 9252 10362
rect 9276 10310 9290 10362
rect 9290 10310 9302 10362
rect 9302 10310 9332 10362
rect 9356 10310 9366 10362
rect 9366 10310 9412 10362
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 9276 10308 9332 10310
rect 9356 10308 9412 10310
rect 10046 10240 10102 10296
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4266 9818
rect 4266 9766 4276 9818
rect 4300 9766 4330 9818
rect 4330 9766 4342 9818
rect 4342 9766 4356 9818
rect 4380 9766 4394 9818
rect 4394 9766 4406 9818
rect 4406 9766 4436 9818
rect 4460 9766 4470 9818
rect 4470 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 7484 9818 7540 9820
rect 7564 9818 7620 9820
rect 7644 9818 7700 9820
rect 7724 9818 7780 9820
rect 7484 9766 7530 9818
rect 7530 9766 7540 9818
rect 7564 9766 7594 9818
rect 7594 9766 7606 9818
rect 7606 9766 7620 9818
rect 7644 9766 7658 9818
rect 7658 9766 7670 9818
rect 7670 9766 7700 9818
rect 7724 9766 7734 9818
rect 7734 9766 7780 9818
rect 7484 9764 7540 9766
rect 7564 9764 7620 9766
rect 7644 9764 7700 9766
rect 7724 9764 7780 9766
rect 10046 9444 10102 9480
rect 10046 9424 10048 9444
rect 10048 9424 10100 9444
rect 10100 9424 10102 9444
rect 5852 9274 5908 9276
rect 5932 9274 5988 9276
rect 6012 9274 6068 9276
rect 6092 9274 6148 9276
rect 5852 9222 5898 9274
rect 5898 9222 5908 9274
rect 5932 9222 5962 9274
rect 5962 9222 5974 9274
rect 5974 9222 5988 9274
rect 6012 9222 6026 9274
rect 6026 9222 6038 9274
rect 6038 9222 6068 9274
rect 6092 9222 6102 9274
rect 6102 9222 6148 9274
rect 5852 9220 5908 9222
rect 5932 9220 5988 9222
rect 6012 9220 6068 9222
rect 6092 9220 6148 9222
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 9276 9274 9332 9276
rect 9356 9274 9412 9276
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9238 9274
rect 9238 9222 9252 9274
rect 9276 9222 9290 9274
rect 9290 9222 9302 9274
rect 9302 9222 9332 9274
rect 9356 9222 9366 9274
rect 9366 9222 9412 9274
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 9276 9220 9332 9222
rect 9356 9220 9412 9222
rect 10046 8780 10048 8800
rect 10048 8780 10100 8800
rect 10100 8780 10102 8800
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4266 8730
rect 4266 8678 4276 8730
rect 4300 8678 4330 8730
rect 4330 8678 4342 8730
rect 4342 8678 4356 8730
rect 4380 8678 4394 8730
rect 4394 8678 4406 8730
rect 4406 8678 4436 8730
rect 4460 8678 4470 8730
rect 4470 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 7484 8730 7540 8732
rect 7564 8730 7620 8732
rect 7644 8730 7700 8732
rect 7724 8730 7780 8732
rect 7484 8678 7530 8730
rect 7530 8678 7540 8730
rect 7564 8678 7594 8730
rect 7594 8678 7606 8730
rect 7606 8678 7620 8730
rect 7644 8678 7658 8730
rect 7658 8678 7670 8730
rect 7670 8678 7700 8730
rect 7724 8678 7734 8730
rect 7734 8678 7780 8730
rect 7484 8676 7540 8678
rect 7564 8676 7620 8678
rect 7644 8676 7700 8678
rect 7724 8676 7780 8678
rect 10046 8744 10102 8780
rect 5852 8186 5908 8188
rect 5932 8186 5988 8188
rect 6012 8186 6068 8188
rect 6092 8186 6148 8188
rect 5852 8134 5898 8186
rect 5898 8134 5908 8186
rect 5932 8134 5962 8186
rect 5962 8134 5974 8186
rect 5974 8134 5988 8186
rect 6012 8134 6026 8186
rect 6026 8134 6038 8186
rect 6038 8134 6068 8186
rect 6092 8134 6102 8186
rect 6102 8134 6148 8186
rect 5852 8132 5908 8134
rect 5932 8132 5988 8134
rect 6012 8132 6068 8134
rect 6092 8132 6148 8134
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 9276 8186 9332 8188
rect 9356 8186 9412 8188
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9238 8186
rect 9238 8134 9252 8186
rect 9276 8134 9290 8186
rect 9290 8134 9302 8186
rect 9302 8134 9332 8186
rect 9356 8134 9366 8186
rect 9366 8134 9412 8186
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 9276 8132 9332 8134
rect 9356 8132 9412 8134
rect 10046 7928 10102 7984
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4266 7642
rect 4266 7590 4276 7642
rect 4300 7590 4330 7642
rect 4330 7590 4342 7642
rect 4342 7590 4356 7642
rect 4380 7590 4394 7642
rect 4394 7590 4406 7642
rect 4406 7590 4436 7642
rect 4460 7590 4470 7642
rect 4470 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 7484 7642 7540 7644
rect 7564 7642 7620 7644
rect 7644 7642 7700 7644
rect 7724 7642 7780 7644
rect 7484 7590 7530 7642
rect 7530 7590 7540 7642
rect 7564 7590 7594 7642
rect 7594 7590 7606 7642
rect 7606 7590 7620 7642
rect 7644 7590 7658 7642
rect 7658 7590 7670 7642
rect 7670 7590 7700 7642
rect 7724 7590 7734 7642
rect 7734 7590 7780 7642
rect 7484 7588 7540 7590
rect 7564 7588 7620 7590
rect 7644 7588 7700 7590
rect 7724 7588 7780 7590
rect 3974 4820 4030 4856
rect 3974 4800 3976 4820
rect 3976 4800 4028 4820
rect 4028 4800 4030 4820
rect 5852 7098 5908 7100
rect 5932 7098 5988 7100
rect 6012 7098 6068 7100
rect 6092 7098 6148 7100
rect 5852 7046 5898 7098
rect 5898 7046 5908 7098
rect 5932 7046 5962 7098
rect 5962 7046 5974 7098
rect 5974 7046 5988 7098
rect 6012 7046 6026 7098
rect 6026 7046 6038 7098
rect 6038 7046 6068 7098
rect 6092 7046 6102 7098
rect 6102 7046 6148 7098
rect 5852 7044 5908 7046
rect 5932 7044 5988 7046
rect 6012 7044 6068 7046
rect 6092 7044 6148 7046
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 9276 7098 9332 7100
rect 9356 7098 9412 7100
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9238 7098
rect 9238 7046 9252 7098
rect 9276 7046 9290 7098
rect 9290 7046 9302 7098
rect 9302 7046 9332 7098
rect 9356 7046 9366 7098
rect 9366 7046 9412 7098
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 9276 7044 9332 7046
rect 9356 7044 9412 7046
rect 10046 7148 10048 7168
rect 10048 7148 10100 7168
rect 10100 7148 10102 7168
rect 10046 7112 10102 7148
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4266 6554
rect 4266 6502 4276 6554
rect 4300 6502 4330 6554
rect 4330 6502 4342 6554
rect 4342 6502 4356 6554
rect 4380 6502 4394 6554
rect 4394 6502 4406 6554
rect 4406 6502 4436 6554
rect 4460 6502 4470 6554
rect 4470 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 7484 6554 7540 6556
rect 7564 6554 7620 6556
rect 7644 6554 7700 6556
rect 7724 6554 7780 6556
rect 7484 6502 7530 6554
rect 7530 6502 7540 6554
rect 7564 6502 7594 6554
rect 7594 6502 7606 6554
rect 7606 6502 7620 6554
rect 7644 6502 7658 6554
rect 7658 6502 7670 6554
rect 7670 6502 7700 6554
rect 7724 6502 7734 6554
rect 7734 6502 7780 6554
rect 7484 6500 7540 6502
rect 7564 6500 7620 6502
rect 7644 6500 7700 6502
rect 7724 6500 7780 6502
rect 5852 6010 5908 6012
rect 5932 6010 5988 6012
rect 6012 6010 6068 6012
rect 6092 6010 6148 6012
rect 5852 5958 5898 6010
rect 5898 5958 5908 6010
rect 5932 5958 5962 6010
rect 5962 5958 5974 6010
rect 5974 5958 5988 6010
rect 6012 5958 6026 6010
rect 6026 5958 6038 6010
rect 6038 5958 6068 6010
rect 6092 5958 6102 6010
rect 6102 5958 6148 6010
rect 5852 5956 5908 5958
rect 5932 5956 5988 5958
rect 6012 5956 6068 5958
rect 6092 5956 6148 5958
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 9276 6010 9332 6012
rect 9356 6010 9412 6012
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9238 6010
rect 9238 5958 9252 6010
rect 9276 5958 9290 6010
rect 9290 5958 9302 6010
rect 9302 5958 9332 6010
rect 9356 5958 9366 6010
rect 9366 5958 9412 6010
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 9276 5956 9332 5958
rect 9356 5956 9412 5958
rect 10046 6432 10102 6488
rect 10046 5616 10102 5672
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4266 5466
rect 4266 5414 4276 5466
rect 4300 5414 4330 5466
rect 4330 5414 4342 5466
rect 4342 5414 4356 5466
rect 4380 5414 4394 5466
rect 4394 5414 4406 5466
rect 4406 5414 4436 5466
rect 4460 5414 4470 5466
rect 4470 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 7484 5466 7540 5468
rect 7564 5466 7620 5468
rect 7644 5466 7700 5468
rect 7724 5466 7780 5468
rect 7484 5414 7530 5466
rect 7530 5414 7540 5466
rect 7564 5414 7594 5466
rect 7594 5414 7606 5466
rect 7606 5414 7620 5466
rect 7644 5414 7658 5466
rect 7658 5414 7670 5466
rect 7670 5414 7700 5466
rect 7724 5414 7734 5466
rect 7734 5414 7780 5466
rect 7484 5412 7540 5414
rect 7564 5412 7620 5414
rect 7644 5412 7700 5414
rect 7724 5412 7780 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4266 4378
rect 4266 4326 4276 4378
rect 4300 4326 4330 4378
rect 4330 4326 4342 4378
rect 4342 4326 4356 4378
rect 4380 4326 4394 4378
rect 4394 4326 4406 4378
rect 4406 4326 4436 4378
rect 4460 4326 4470 4378
rect 4470 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 5852 4922 5908 4924
rect 5932 4922 5988 4924
rect 6012 4922 6068 4924
rect 6092 4922 6148 4924
rect 5852 4870 5898 4922
rect 5898 4870 5908 4922
rect 5932 4870 5962 4922
rect 5962 4870 5974 4922
rect 5974 4870 5988 4922
rect 6012 4870 6026 4922
rect 6026 4870 6038 4922
rect 6038 4870 6068 4922
rect 6092 4870 6102 4922
rect 6102 4870 6148 4922
rect 5852 4868 5908 4870
rect 5932 4868 5988 4870
rect 6012 4868 6068 4870
rect 6092 4868 6148 4870
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 9276 4922 9332 4924
rect 9356 4922 9412 4924
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9238 4922
rect 9238 4870 9252 4922
rect 9276 4870 9290 4922
rect 9290 4870 9302 4922
rect 9302 4870 9332 4922
rect 9356 4870 9366 4922
rect 9366 4870 9412 4922
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 9276 4868 9332 4870
rect 9356 4868 9412 4870
rect 10046 4800 10102 4856
rect 7484 4378 7540 4380
rect 7564 4378 7620 4380
rect 7644 4378 7700 4380
rect 7724 4378 7780 4380
rect 7484 4326 7530 4378
rect 7530 4326 7540 4378
rect 7564 4326 7594 4378
rect 7594 4326 7606 4378
rect 7606 4326 7620 4378
rect 7644 4326 7658 4378
rect 7658 4326 7670 4378
rect 7670 4326 7700 4378
rect 7724 4326 7734 4378
rect 7734 4326 7780 4378
rect 7484 4324 7540 4326
rect 7564 4324 7620 4326
rect 7644 4324 7700 4326
rect 7724 4324 7780 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4266 3290
rect 4266 3238 4276 3290
rect 4300 3238 4330 3290
rect 4330 3238 4342 3290
rect 4342 3238 4356 3290
rect 4380 3238 4394 3290
rect 4394 3238 4406 3290
rect 4406 3238 4436 3290
rect 4460 3238 4470 3290
rect 4470 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4066 2488 4122 2544
rect 5852 3834 5908 3836
rect 5932 3834 5988 3836
rect 6012 3834 6068 3836
rect 6092 3834 6148 3836
rect 5852 3782 5898 3834
rect 5898 3782 5908 3834
rect 5932 3782 5962 3834
rect 5962 3782 5974 3834
rect 5974 3782 5988 3834
rect 6012 3782 6026 3834
rect 6026 3782 6038 3834
rect 6038 3782 6068 3834
rect 6092 3782 6102 3834
rect 6102 3782 6148 3834
rect 5852 3780 5908 3782
rect 5932 3780 5988 3782
rect 6012 3780 6068 3782
rect 6092 3780 6148 3782
rect 7484 3290 7540 3292
rect 7564 3290 7620 3292
rect 7644 3290 7700 3292
rect 7724 3290 7780 3292
rect 7484 3238 7530 3290
rect 7530 3238 7540 3290
rect 7564 3238 7594 3290
rect 7594 3238 7606 3290
rect 7606 3238 7620 3290
rect 7644 3238 7658 3290
rect 7658 3238 7670 3290
rect 7670 3238 7700 3290
rect 7724 3238 7734 3290
rect 7734 3238 7780 3290
rect 7484 3236 7540 3238
rect 7564 3236 7620 3238
rect 7644 3236 7700 3238
rect 7724 3236 7780 3238
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 9276 3834 9332 3836
rect 9356 3834 9412 3836
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9238 3834
rect 9238 3782 9252 3834
rect 9276 3782 9290 3834
rect 9290 3782 9302 3834
rect 9302 3782 9332 3834
rect 9356 3782 9366 3834
rect 9366 3782 9412 3834
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 9276 3780 9332 3782
rect 9356 3780 9412 3782
rect 10046 4120 10102 4176
rect 10046 3340 10048 3360
rect 10048 3340 10100 3360
rect 10100 3340 10102 3360
rect 10046 3304 10102 3340
rect 5852 2746 5908 2748
rect 5932 2746 5988 2748
rect 6012 2746 6068 2748
rect 6092 2746 6148 2748
rect 5852 2694 5898 2746
rect 5898 2694 5908 2746
rect 5932 2694 5962 2746
rect 5962 2694 5974 2746
rect 5974 2694 5988 2746
rect 6012 2694 6026 2746
rect 6026 2694 6038 2746
rect 6038 2694 6068 2746
rect 6092 2694 6102 2746
rect 6102 2694 6148 2746
rect 5852 2692 5908 2694
rect 5932 2692 5988 2694
rect 6012 2692 6068 2694
rect 6092 2692 6148 2694
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 9276 2746 9332 2748
rect 9356 2746 9412 2748
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9238 2746
rect 9238 2694 9252 2746
rect 9276 2694 9290 2746
rect 9290 2694 9302 2746
rect 9302 2694 9332 2746
rect 9356 2694 9366 2746
rect 9366 2694 9412 2746
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 9276 2692 9332 2694
rect 9356 2692 9412 2694
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4266 2202
rect 4266 2150 4276 2202
rect 4300 2150 4330 2202
rect 4330 2150 4342 2202
rect 4342 2150 4356 2202
rect 4380 2150 4394 2202
rect 4394 2150 4406 2202
rect 4406 2150 4436 2202
rect 4460 2150 4470 2202
rect 4470 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 4066 1808 4122 1864
rect 3974 1400 4030 1456
rect 7484 2202 7540 2204
rect 7564 2202 7620 2204
rect 7644 2202 7700 2204
rect 7724 2202 7780 2204
rect 7484 2150 7530 2202
rect 7530 2150 7540 2202
rect 7564 2150 7594 2202
rect 7594 2150 7606 2202
rect 7606 2150 7620 2202
rect 7644 2150 7658 2202
rect 7658 2150 7670 2202
rect 7670 2150 7700 2202
rect 7724 2150 7734 2202
rect 7734 2150 7780 2202
rect 7484 2148 7540 2150
rect 7564 2148 7620 2150
rect 7644 2148 7700 2150
rect 7724 2148 7780 2150
rect 2870 584 2926 640
rect 1398 176 1454 232
rect 10046 2488 10102 2544
rect 9494 1808 9550 1864
rect 9586 992 9642 1048
rect 9310 312 9366 368
<< metal3 >>
rect 0 79658 800 79688
rect 2957 79658 3023 79661
rect 0 79656 3023 79658
rect 0 79600 2962 79656
rect 3018 79600 3023 79656
rect 0 79598 3023 79600
rect 0 79568 800 79598
rect 2957 79595 3023 79598
rect 9949 79522 10015 79525
rect 11200 79522 12000 79552
rect 9949 79520 12000 79522
rect 9949 79464 9954 79520
rect 10010 79464 12000 79520
rect 9949 79462 12000 79464
rect 9949 79459 10015 79462
rect 11200 79432 12000 79462
rect 0 79250 800 79280
rect 1393 79250 1459 79253
rect 0 79248 1459 79250
rect 0 79192 1398 79248
rect 1454 79192 1459 79248
rect 0 79190 1459 79192
rect 0 79160 800 79190
rect 1393 79187 1459 79190
rect 0 78842 800 78872
rect 3693 78842 3759 78845
rect 0 78840 3759 78842
rect 0 78784 3698 78840
rect 3754 78784 3759 78840
rect 0 78782 3759 78784
rect 0 78752 800 78782
rect 3693 78779 3759 78782
rect 9581 78706 9647 78709
rect 11200 78706 12000 78736
rect 9581 78704 12000 78706
rect 9581 78648 9586 78704
rect 9642 78648 12000 78704
rect 9581 78646 12000 78648
rect 9581 78643 9647 78646
rect 11200 78616 12000 78646
rect 0 78434 800 78464
rect 4061 78434 4127 78437
rect 0 78432 4127 78434
rect 0 78376 4066 78432
rect 4122 78376 4127 78432
rect 0 78374 4127 78376
rect 0 78344 800 78374
rect 4061 78371 4127 78374
rect 0 78026 800 78056
rect 3417 78026 3483 78029
rect 0 78024 3483 78026
rect 0 77968 3422 78024
rect 3478 77968 3483 78024
rect 0 77966 3483 77968
rect 0 77936 800 77966
rect 3417 77963 3483 77966
rect 9489 78026 9555 78029
rect 11200 78026 12000 78056
rect 9489 78024 12000 78026
rect 9489 77968 9494 78024
rect 9550 77968 12000 78024
rect 9489 77966 12000 77968
rect 9489 77963 9555 77966
rect 11200 77936 12000 77966
rect 2576 77824 2896 77825
rect 2576 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2576 77759 2896 77760
rect 5840 77824 6160 77825
rect 5840 77760 5848 77824
rect 5912 77760 5928 77824
rect 5992 77760 6008 77824
rect 6072 77760 6088 77824
rect 6152 77760 6160 77824
rect 5840 77759 6160 77760
rect 9104 77824 9424 77825
rect 9104 77760 9112 77824
rect 9176 77760 9192 77824
rect 9256 77760 9272 77824
rect 9336 77760 9352 77824
rect 9416 77760 9424 77824
rect 9104 77759 9424 77760
rect 0 77618 800 77648
rect 3969 77618 4035 77621
rect 0 77616 4035 77618
rect 0 77560 3974 77616
rect 4030 77560 4035 77616
rect 0 77558 4035 77560
rect 0 77528 800 77558
rect 3969 77555 4035 77558
rect 4208 77280 4528 77281
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 77215 4528 77216
rect 7472 77280 7792 77281
rect 7472 77216 7480 77280
rect 7544 77216 7560 77280
rect 7624 77216 7640 77280
rect 7704 77216 7720 77280
rect 7784 77216 7792 77280
rect 7472 77215 7792 77216
rect 9397 77210 9463 77213
rect 11200 77210 12000 77240
rect 9397 77208 12000 77210
rect 9397 77152 9402 77208
rect 9458 77152 12000 77208
rect 9397 77150 12000 77152
rect 9397 77147 9463 77150
rect 11200 77120 12000 77150
rect 0 77074 800 77104
rect 2957 77074 3023 77077
rect 0 77072 3023 77074
rect 0 77016 2962 77072
rect 3018 77016 3023 77072
rect 0 77014 3023 77016
rect 0 76984 800 77014
rect 2957 77011 3023 77014
rect 2576 76736 2896 76737
rect 0 76666 800 76696
rect 2576 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2576 76671 2896 76672
rect 5840 76736 6160 76737
rect 5840 76672 5848 76736
rect 5912 76672 5928 76736
rect 5992 76672 6008 76736
rect 6072 76672 6088 76736
rect 6152 76672 6160 76736
rect 5840 76671 6160 76672
rect 9104 76736 9424 76737
rect 9104 76672 9112 76736
rect 9176 76672 9192 76736
rect 9256 76672 9272 76736
rect 9336 76672 9352 76736
rect 9416 76672 9424 76736
rect 9104 76671 9424 76672
rect 0 76606 1778 76666
rect 0 76576 800 76606
rect 1718 76530 1778 76606
rect 3325 76530 3391 76533
rect 1718 76528 3391 76530
rect 1718 76472 3330 76528
rect 3386 76472 3391 76528
rect 1718 76470 3391 76472
rect 3325 76467 3391 76470
rect 10133 76394 10199 76397
rect 11200 76394 12000 76424
rect 10133 76392 12000 76394
rect 10133 76336 10138 76392
rect 10194 76336 12000 76392
rect 10133 76334 12000 76336
rect 10133 76331 10199 76334
rect 11200 76304 12000 76334
rect 0 76258 800 76288
rect 3969 76258 4035 76261
rect 0 76256 4035 76258
rect 0 76200 3974 76256
rect 4030 76200 4035 76256
rect 0 76198 4035 76200
rect 0 76168 800 76198
rect 3969 76195 4035 76198
rect 4208 76192 4528 76193
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 76127 4528 76128
rect 7472 76192 7792 76193
rect 7472 76128 7480 76192
rect 7544 76128 7560 76192
rect 7624 76128 7640 76192
rect 7704 76128 7720 76192
rect 7784 76128 7792 76192
rect 7472 76127 7792 76128
rect 0 75850 800 75880
rect 2497 75850 2563 75853
rect 0 75848 2563 75850
rect 0 75792 2502 75848
rect 2558 75792 2563 75848
rect 0 75790 2563 75792
rect 0 75760 800 75790
rect 2497 75787 2563 75790
rect 10133 75714 10199 75717
rect 11200 75714 12000 75744
rect 10133 75712 12000 75714
rect 10133 75656 10138 75712
rect 10194 75656 12000 75712
rect 10133 75654 12000 75656
rect 10133 75651 10199 75654
rect 2576 75648 2896 75649
rect 2576 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2576 75583 2896 75584
rect 5840 75648 6160 75649
rect 5840 75584 5848 75648
rect 5912 75584 5928 75648
rect 5992 75584 6008 75648
rect 6072 75584 6088 75648
rect 6152 75584 6160 75648
rect 5840 75583 6160 75584
rect 9104 75648 9424 75649
rect 9104 75584 9112 75648
rect 9176 75584 9192 75648
rect 9256 75584 9272 75648
rect 9336 75584 9352 75648
rect 9416 75584 9424 75648
rect 11200 75624 12000 75654
rect 9104 75583 9424 75584
rect 0 75442 800 75472
rect 3693 75442 3759 75445
rect 0 75440 3759 75442
rect 0 75384 3698 75440
rect 3754 75384 3759 75440
rect 0 75382 3759 75384
rect 0 75352 800 75382
rect 3693 75379 3759 75382
rect 4208 75104 4528 75105
rect 0 75034 800 75064
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 75039 4528 75040
rect 7472 75104 7792 75105
rect 7472 75040 7480 75104
rect 7544 75040 7560 75104
rect 7624 75040 7640 75104
rect 7704 75040 7720 75104
rect 7784 75040 7792 75104
rect 7472 75039 7792 75040
rect 1393 75034 1459 75037
rect 0 75032 1459 75034
rect 0 74976 1398 75032
rect 1454 74976 1459 75032
rect 0 74974 1459 74976
rect 0 74944 800 74974
rect 1393 74971 1459 74974
rect 2497 75034 2563 75037
rect 3918 75034 3924 75036
rect 2497 75032 3924 75034
rect 2497 74976 2502 75032
rect 2558 74976 3924 75032
rect 2497 74974 3924 74976
rect 2497 74971 2563 74974
rect 3918 74972 3924 74974
rect 3988 74972 3994 75036
rect 10133 74898 10199 74901
rect 11200 74898 12000 74928
rect 10133 74896 12000 74898
rect 10133 74840 10138 74896
rect 10194 74840 12000 74896
rect 10133 74838 12000 74840
rect 10133 74835 10199 74838
rect 11200 74808 12000 74838
rect 0 74626 800 74656
rect 1577 74626 1643 74629
rect 0 74624 1643 74626
rect 0 74568 1582 74624
rect 1638 74568 1643 74624
rect 0 74566 1643 74568
rect 0 74536 800 74566
rect 1577 74563 1643 74566
rect 2576 74560 2896 74561
rect 2576 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2576 74495 2896 74496
rect 5840 74560 6160 74561
rect 5840 74496 5848 74560
rect 5912 74496 5928 74560
rect 5992 74496 6008 74560
rect 6072 74496 6088 74560
rect 6152 74496 6160 74560
rect 5840 74495 6160 74496
rect 9104 74560 9424 74561
rect 9104 74496 9112 74560
rect 9176 74496 9192 74560
rect 9256 74496 9272 74560
rect 9336 74496 9352 74560
rect 9416 74496 9424 74560
rect 9104 74495 9424 74496
rect 0 74082 800 74112
rect 2957 74082 3023 74085
rect 0 74080 3023 74082
rect 0 74024 2962 74080
rect 3018 74024 3023 74080
rect 0 74022 3023 74024
rect 0 73992 800 74022
rect 2957 74019 3023 74022
rect 10133 74082 10199 74085
rect 11200 74082 12000 74112
rect 10133 74080 12000 74082
rect 10133 74024 10138 74080
rect 10194 74024 12000 74080
rect 10133 74022 12000 74024
rect 10133 74019 10199 74022
rect 4208 74016 4528 74017
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 73951 4528 73952
rect 7472 74016 7792 74017
rect 7472 73952 7480 74016
rect 7544 73952 7560 74016
rect 7624 73952 7640 74016
rect 7704 73952 7720 74016
rect 7784 73952 7792 74016
rect 11200 73992 12000 74022
rect 7472 73951 7792 73952
rect 0 73674 800 73704
rect 2865 73674 2931 73677
rect 0 73672 2931 73674
rect 0 73616 2870 73672
rect 2926 73616 2931 73672
rect 0 73614 2931 73616
rect 0 73584 800 73614
rect 2865 73611 2931 73614
rect 2576 73472 2896 73473
rect 2576 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2576 73407 2896 73408
rect 5840 73472 6160 73473
rect 5840 73408 5848 73472
rect 5912 73408 5928 73472
rect 5992 73408 6008 73472
rect 6072 73408 6088 73472
rect 6152 73408 6160 73472
rect 5840 73407 6160 73408
rect 9104 73472 9424 73473
rect 9104 73408 9112 73472
rect 9176 73408 9192 73472
rect 9256 73408 9272 73472
rect 9336 73408 9352 73472
rect 9416 73408 9424 73472
rect 9104 73407 9424 73408
rect 10133 73402 10199 73405
rect 11200 73402 12000 73432
rect 10133 73400 12000 73402
rect 10133 73344 10138 73400
rect 10194 73344 12000 73400
rect 10133 73342 12000 73344
rect 10133 73339 10199 73342
rect 11200 73312 12000 73342
rect 0 73266 800 73296
rect 2221 73266 2287 73269
rect 0 73264 2287 73266
rect 0 73208 2226 73264
rect 2282 73208 2287 73264
rect 0 73206 2287 73208
rect 0 73176 800 73206
rect 2221 73203 2287 73206
rect 4208 72928 4528 72929
rect 0 72858 800 72888
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 72863 4528 72864
rect 7472 72928 7792 72929
rect 7472 72864 7480 72928
rect 7544 72864 7560 72928
rect 7624 72864 7640 72928
rect 7704 72864 7720 72928
rect 7784 72864 7792 72928
rect 7472 72863 7792 72864
rect 1393 72858 1459 72861
rect 0 72856 1459 72858
rect 0 72800 1398 72856
rect 1454 72800 1459 72856
rect 0 72798 1459 72800
rect 0 72768 800 72798
rect 1393 72795 1459 72798
rect 1117 72722 1183 72725
rect 2681 72722 2747 72725
rect 1117 72720 2747 72722
rect 1117 72664 1122 72720
rect 1178 72664 2686 72720
rect 2742 72664 2747 72720
rect 1117 72662 2747 72664
rect 1117 72659 1183 72662
rect 2681 72659 2747 72662
rect 10133 72586 10199 72589
rect 11200 72586 12000 72616
rect 10133 72584 12000 72586
rect 10133 72528 10138 72584
rect 10194 72528 12000 72584
rect 10133 72526 12000 72528
rect 10133 72523 10199 72526
rect 11200 72496 12000 72526
rect 0 72450 800 72480
rect 1577 72450 1643 72453
rect 0 72448 1643 72450
rect 0 72392 1582 72448
rect 1638 72392 1643 72448
rect 0 72390 1643 72392
rect 0 72360 800 72390
rect 1577 72387 1643 72390
rect 2576 72384 2896 72385
rect 2576 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2576 72319 2896 72320
rect 5840 72384 6160 72385
rect 5840 72320 5848 72384
rect 5912 72320 5928 72384
rect 5992 72320 6008 72384
rect 6072 72320 6088 72384
rect 6152 72320 6160 72384
rect 5840 72319 6160 72320
rect 9104 72384 9424 72385
rect 9104 72320 9112 72384
rect 9176 72320 9192 72384
rect 9256 72320 9272 72384
rect 9336 72320 9352 72384
rect 9416 72320 9424 72384
rect 9104 72319 9424 72320
rect 0 72042 800 72072
rect 2865 72042 2931 72045
rect 0 72040 2931 72042
rect 0 71984 2870 72040
rect 2926 71984 2931 72040
rect 0 71982 2931 71984
rect 0 71952 800 71982
rect 2865 71979 2931 71982
rect 4208 71840 4528 71841
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 71775 4528 71776
rect 7472 71840 7792 71841
rect 7472 71776 7480 71840
rect 7544 71776 7560 71840
rect 7624 71776 7640 71840
rect 7704 71776 7720 71840
rect 7784 71776 7792 71840
rect 7472 71775 7792 71776
rect 10133 71770 10199 71773
rect 11200 71770 12000 71800
rect 10133 71768 12000 71770
rect 10133 71712 10138 71768
rect 10194 71712 12000 71768
rect 10133 71710 12000 71712
rect 10133 71707 10199 71710
rect 11200 71680 12000 71710
rect 0 71634 800 71664
rect 2221 71634 2287 71637
rect 0 71632 2287 71634
rect 0 71576 2226 71632
rect 2282 71576 2287 71632
rect 0 71574 2287 71576
rect 0 71544 800 71574
rect 2221 71571 2287 71574
rect 2576 71296 2896 71297
rect 2576 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2576 71231 2896 71232
rect 5840 71296 6160 71297
rect 5840 71232 5848 71296
rect 5912 71232 5928 71296
rect 5992 71232 6008 71296
rect 6072 71232 6088 71296
rect 6152 71232 6160 71296
rect 5840 71231 6160 71232
rect 9104 71296 9424 71297
rect 9104 71232 9112 71296
rect 9176 71232 9192 71296
rect 9256 71232 9272 71296
rect 9336 71232 9352 71296
rect 9416 71232 9424 71296
rect 9104 71231 9424 71232
rect 0 71090 800 71120
rect 1577 71090 1643 71093
rect 0 71088 1643 71090
rect 0 71032 1582 71088
rect 1638 71032 1643 71088
rect 0 71030 1643 71032
rect 0 71000 800 71030
rect 1577 71027 1643 71030
rect 10133 71090 10199 71093
rect 11200 71090 12000 71120
rect 10133 71088 12000 71090
rect 10133 71032 10138 71088
rect 10194 71032 12000 71088
rect 10133 71030 12000 71032
rect 10133 71027 10199 71030
rect 11200 71000 12000 71030
rect 4208 70752 4528 70753
rect 0 70682 800 70712
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 70687 4528 70688
rect 7472 70752 7792 70753
rect 7472 70688 7480 70752
rect 7544 70688 7560 70752
rect 7624 70688 7640 70752
rect 7704 70688 7720 70752
rect 7784 70688 7792 70752
rect 7472 70687 7792 70688
rect 1577 70682 1643 70685
rect 0 70680 1643 70682
rect 0 70624 1582 70680
rect 1638 70624 1643 70680
rect 0 70622 1643 70624
rect 0 70592 800 70622
rect 1577 70619 1643 70622
rect 0 70274 800 70304
rect 1577 70274 1643 70277
rect 0 70272 1643 70274
rect 0 70216 1582 70272
rect 1638 70216 1643 70272
rect 0 70214 1643 70216
rect 0 70184 800 70214
rect 1577 70211 1643 70214
rect 10133 70274 10199 70277
rect 11200 70274 12000 70304
rect 10133 70272 12000 70274
rect 10133 70216 10138 70272
rect 10194 70216 12000 70272
rect 10133 70214 12000 70216
rect 10133 70211 10199 70214
rect 2576 70208 2896 70209
rect 2576 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2576 70143 2896 70144
rect 5840 70208 6160 70209
rect 5840 70144 5848 70208
rect 5912 70144 5928 70208
rect 5992 70144 6008 70208
rect 6072 70144 6088 70208
rect 6152 70144 6160 70208
rect 5840 70143 6160 70144
rect 9104 70208 9424 70209
rect 9104 70144 9112 70208
rect 9176 70144 9192 70208
rect 9256 70144 9272 70208
rect 9336 70144 9352 70208
rect 9416 70144 9424 70208
rect 11200 70184 12000 70214
rect 9104 70143 9424 70144
rect 0 69866 800 69896
rect 2037 69866 2103 69869
rect 0 69864 2103 69866
rect 0 69808 2042 69864
rect 2098 69808 2103 69864
rect 0 69806 2103 69808
rect 0 69776 800 69806
rect 2037 69803 2103 69806
rect 4208 69664 4528 69665
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 69599 4528 69600
rect 7472 69664 7792 69665
rect 7472 69600 7480 69664
rect 7544 69600 7560 69664
rect 7624 69600 7640 69664
rect 7704 69600 7720 69664
rect 7784 69600 7792 69664
rect 7472 69599 7792 69600
rect 0 69458 800 69488
rect 2865 69458 2931 69461
rect 0 69456 2931 69458
rect 0 69400 2870 69456
rect 2926 69400 2931 69456
rect 0 69398 2931 69400
rect 0 69368 800 69398
rect 2865 69395 2931 69398
rect 10133 69458 10199 69461
rect 11200 69458 12000 69488
rect 10133 69456 12000 69458
rect 10133 69400 10138 69456
rect 10194 69400 12000 69456
rect 10133 69398 12000 69400
rect 10133 69395 10199 69398
rect 11200 69368 12000 69398
rect 2262 69260 2268 69324
rect 2332 69322 2338 69324
rect 2681 69322 2747 69325
rect 2332 69320 2747 69322
rect 2332 69264 2686 69320
rect 2742 69264 2747 69320
rect 2332 69262 2747 69264
rect 2332 69260 2338 69262
rect 2681 69259 2747 69262
rect 2576 69120 2896 69121
rect 0 69050 800 69080
rect 2576 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2576 69055 2896 69056
rect 5840 69120 6160 69121
rect 5840 69056 5848 69120
rect 5912 69056 5928 69120
rect 5992 69056 6008 69120
rect 6072 69056 6088 69120
rect 6152 69056 6160 69120
rect 5840 69055 6160 69056
rect 9104 69120 9424 69121
rect 9104 69056 9112 69120
rect 9176 69056 9192 69120
rect 9256 69056 9272 69120
rect 9336 69056 9352 69120
rect 9416 69056 9424 69120
rect 9104 69055 9424 69056
rect 2221 69050 2287 69053
rect 0 69048 2287 69050
rect 0 68992 2226 69048
rect 2282 68992 2287 69048
rect 0 68990 2287 68992
rect 0 68960 800 68990
rect 2221 68987 2287 68990
rect 10133 68778 10199 68781
rect 11200 68778 12000 68808
rect 10133 68776 12000 68778
rect 10133 68720 10138 68776
rect 10194 68720 12000 68776
rect 10133 68718 12000 68720
rect 10133 68715 10199 68718
rect 11200 68688 12000 68718
rect 0 68642 800 68672
rect 2957 68642 3023 68645
rect 0 68640 3023 68642
rect 0 68584 2962 68640
rect 3018 68584 3023 68640
rect 0 68582 3023 68584
rect 0 68552 800 68582
rect 2957 68579 3023 68582
rect 4208 68576 4528 68577
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 68511 4528 68512
rect 7472 68576 7792 68577
rect 7472 68512 7480 68576
rect 7544 68512 7560 68576
rect 7624 68512 7640 68576
rect 7704 68512 7720 68576
rect 7784 68512 7792 68576
rect 7472 68511 7792 68512
rect 0 68098 800 68128
rect 1577 68098 1643 68101
rect 0 68096 1643 68098
rect 0 68040 1582 68096
rect 1638 68040 1643 68096
rect 0 68038 1643 68040
rect 0 68008 800 68038
rect 1577 68035 1643 68038
rect 2576 68032 2896 68033
rect 2576 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2576 67967 2896 67968
rect 5840 68032 6160 68033
rect 5840 67968 5848 68032
rect 5912 67968 5928 68032
rect 5992 67968 6008 68032
rect 6072 67968 6088 68032
rect 6152 67968 6160 68032
rect 5840 67967 6160 67968
rect 9104 68032 9424 68033
rect 9104 67968 9112 68032
rect 9176 67968 9192 68032
rect 9256 67968 9272 68032
rect 9336 67968 9352 68032
rect 9416 67968 9424 68032
rect 9104 67967 9424 67968
rect 10133 67962 10199 67965
rect 11200 67962 12000 67992
rect 10133 67960 12000 67962
rect 10133 67904 10138 67960
rect 10194 67904 12000 67960
rect 10133 67902 12000 67904
rect 10133 67899 10199 67902
rect 11200 67872 12000 67902
rect 0 67690 800 67720
rect 1301 67690 1367 67693
rect 0 67688 1367 67690
rect 0 67632 1306 67688
rect 1362 67632 1367 67688
rect 0 67630 1367 67632
rect 0 67600 800 67630
rect 1301 67627 1367 67630
rect 1669 67692 1735 67693
rect 1669 67688 1716 67692
rect 1780 67690 1786 67692
rect 1669 67632 1674 67688
rect 1669 67628 1716 67632
rect 1780 67630 1826 67690
rect 1780 67628 1786 67630
rect 1669 67627 1735 67628
rect 4208 67488 4528 67489
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 67423 4528 67424
rect 7472 67488 7792 67489
rect 7472 67424 7480 67488
rect 7544 67424 7560 67488
rect 7624 67424 7640 67488
rect 7704 67424 7720 67488
rect 7784 67424 7792 67488
rect 7472 67423 7792 67424
rect 2078 67356 2084 67420
rect 2148 67418 2154 67420
rect 2221 67418 2287 67421
rect 2148 67416 2287 67418
rect 2148 67360 2226 67416
rect 2282 67360 2287 67416
rect 2148 67358 2287 67360
rect 2148 67356 2154 67358
rect 2221 67355 2287 67358
rect 0 67282 800 67312
rect 1393 67282 1459 67285
rect 0 67280 1459 67282
rect 0 67224 1398 67280
rect 1454 67224 1459 67280
rect 0 67222 1459 67224
rect 0 67192 800 67222
rect 1393 67219 1459 67222
rect 10133 67146 10199 67149
rect 11200 67146 12000 67176
rect 10133 67144 12000 67146
rect 10133 67088 10138 67144
rect 10194 67088 12000 67144
rect 10133 67086 12000 67088
rect 10133 67083 10199 67086
rect 11200 67056 12000 67086
rect 2576 66944 2896 66945
rect 0 66874 800 66904
rect 2576 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2576 66879 2896 66880
rect 5840 66944 6160 66945
rect 5840 66880 5848 66944
rect 5912 66880 5928 66944
rect 5992 66880 6008 66944
rect 6072 66880 6088 66944
rect 6152 66880 6160 66944
rect 5840 66879 6160 66880
rect 9104 66944 9424 66945
rect 9104 66880 9112 66944
rect 9176 66880 9192 66944
rect 9256 66880 9272 66944
rect 9336 66880 9352 66944
rect 9416 66880 9424 66944
rect 9104 66879 9424 66880
rect 1393 66874 1459 66877
rect 0 66872 1459 66874
rect 0 66816 1398 66872
rect 1454 66816 1459 66872
rect 0 66814 1459 66816
rect 0 66784 800 66814
rect 1393 66811 1459 66814
rect 0 66466 800 66496
rect 3049 66466 3115 66469
rect 0 66464 3115 66466
rect 0 66408 3054 66464
rect 3110 66408 3115 66464
rect 0 66406 3115 66408
rect 0 66376 800 66406
rect 3049 66403 3115 66406
rect 10133 66466 10199 66469
rect 11200 66466 12000 66496
rect 10133 66464 12000 66466
rect 10133 66408 10138 66464
rect 10194 66408 12000 66464
rect 10133 66406 12000 66408
rect 10133 66403 10199 66406
rect 4208 66400 4528 66401
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 66335 4528 66336
rect 7472 66400 7792 66401
rect 7472 66336 7480 66400
rect 7544 66336 7560 66400
rect 7624 66336 7640 66400
rect 7704 66336 7720 66400
rect 7784 66336 7792 66400
rect 11200 66376 12000 66406
rect 7472 66335 7792 66336
rect 1577 66194 1643 66197
rect 5441 66194 5507 66197
rect 1577 66192 5507 66194
rect 1577 66136 1582 66192
rect 1638 66136 5446 66192
rect 5502 66136 5507 66192
rect 1577 66134 5507 66136
rect 1577 66131 1643 66134
rect 5441 66131 5507 66134
rect 0 66058 800 66088
rect 1577 66058 1643 66061
rect 0 66056 1643 66058
rect 0 66000 1582 66056
rect 1638 66000 1643 66056
rect 0 65998 1643 66000
rect 0 65968 800 65998
rect 1577 65995 1643 65998
rect 2576 65856 2896 65857
rect 2576 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2576 65791 2896 65792
rect 5840 65856 6160 65857
rect 5840 65792 5848 65856
rect 5912 65792 5928 65856
rect 5992 65792 6008 65856
rect 6072 65792 6088 65856
rect 6152 65792 6160 65856
rect 5840 65791 6160 65792
rect 9104 65856 9424 65857
rect 9104 65792 9112 65856
rect 9176 65792 9192 65856
rect 9256 65792 9272 65856
rect 9336 65792 9352 65856
rect 9416 65792 9424 65856
rect 9104 65791 9424 65792
rect 0 65650 800 65680
rect 2957 65650 3023 65653
rect 0 65648 3023 65650
rect 0 65592 2962 65648
rect 3018 65592 3023 65648
rect 0 65590 3023 65592
rect 0 65560 800 65590
rect 2957 65587 3023 65590
rect 10133 65650 10199 65653
rect 11200 65650 12000 65680
rect 10133 65648 12000 65650
rect 10133 65592 10138 65648
rect 10194 65592 12000 65648
rect 10133 65590 12000 65592
rect 10133 65587 10199 65590
rect 11200 65560 12000 65590
rect 4208 65312 4528 65313
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 65247 4528 65248
rect 7472 65312 7792 65313
rect 7472 65248 7480 65312
rect 7544 65248 7560 65312
rect 7624 65248 7640 65312
rect 7704 65248 7720 65312
rect 7784 65248 7792 65312
rect 7472 65247 7792 65248
rect 0 65106 800 65136
rect 3969 65106 4035 65109
rect 0 65104 4035 65106
rect 0 65048 3974 65104
rect 4030 65048 4035 65104
rect 0 65046 4035 65048
rect 0 65016 800 65046
rect 3969 65043 4035 65046
rect 1342 64908 1348 64972
rect 1412 64970 1418 64972
rect 1485 64970 1551 64973
rect 1412 64968 1551 64970
rect 1412 64912 1490 64968
rect 1546 64912 1551 64968
rect 1412 64910 1551 64912
rect 1412 64908 1418 64910
rect 1485 64907 1551 64910
rect 10133 64834 10199 64837
rect 11200 64834 12000 64864
rect 10133 64832 12000 64834
rect 10133 64776 10138 64832
rect 10194 64776 12000 64832
rect 10133 64774 12000 64776
rect 10133 64771 10199 64774
rect 2576 64768 2896 64769
rect 0 64698 800 64728
rect 2576 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2576 64703 2896 64704
rect 5840 64768 6160 64769
rect 5840 64704 5848 64768
rect 5912 64704 5928 64768
rect 5992 64704 6008 64768
rect 6072 64704 6088 64768
rect 6152 64704 6160 64768
rect 5840 64703 6160 64704
rect 9104 64768 9424 64769
rect 9104 64704 9112 64768
rect 9176 64704 9192 64768
rect 9256 64704 9272 64768
rect 9336 64704 9352 64768
rect 9416 64704 9424 64768
rect 11200 64744 12000 64774
rect 9104 64703 9424 64704
rect 0 64638 1410 64698
rect 0 64608 800 64638
rect 1350 64562 1410 64638
rect 3049 64562 3115 64565
rect 1350 64560 3115 64562
rect 1350 64504 3054 64560
rect 3110 64504 3115 64560
rect 1350 64502 3115 64504
rect 3049 64499 3115 64502
rect 0 64290 800 64320
rect 3049 64290 3115 64293
rect 0 64288 3115 64290
rect 0 64232 3054 64288
rect 3110 64232 3115 64288
rect 0 64230 3115 64232
rect 0 64200 800 64230
rect 3049 64227 3115 64230
rect 4208 64224 4528 64225
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 64159 4528 64160
rect 7472 64224 7792 64225
rect 7472 64160 7480 64224
rect 7544 64160 7560 64224
rect 7624 64160 7640 64224
rect 7704 64160 7720 64224
rect 7784 64160 7792 64224
rect 7472 64159 7792 64160
rect 2221 64156 2287 64157
rect 2221 64154 2268 64156
rect 2176 64152 2268 64154
rect 2176 64096 2226 64152
rect 2176 64094 2268 64096
rect 2221 64092 2268 64094
rect 2332 64092 2338 64156
rect 10133 64154 10199 64157
rect 11200 64154 12000 64184
rect 10133 64152 12000 64154
rect 10133 64096 10138 64152
rect 10194 64096 12000 64152
rect 10133 64094 12000 64096
rect 2221 64091 2287 64092
rect 10133 64091 10199 64094
rect 11200 64064 12000 64094
rect 0 63882 800 63912
rect 3049 63882 3115 63885
rect 0 63880 3115 63882
rect 0 63824 3054 63880
rect 3110 63824 3115 63880
rect 0 63822 3115 63824
rect 0 63792 800 63822
rect 3049 63819 3115 63822
rect 2576 63680 2896 63681
rect 2576 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2576 63615 2896 63616
rect 5840 63680 6160 63681
rect 5840 63616 5848 63680
rect 5912 63616 5928 63680
rect 5992 63616 6008 63680
rect 6072 63616 6088 63680
rect 6152 63616 6160 63680
rect 5840 63615 6160 63616
rect 9104 63680 9424 63681
rect 9104 63616 9112 63680
rect 9176 63616 9192 63680
rect 9256 63616 9272 63680
rect 9336 63616 9352 63680
rect 9416 63616 9424 63680
rect 9104 63615 9424 63616
rect 0 63474 800 63504
rect 1669 63474 1735 63477
rect 0 63472 1735 63474
rect 0 63416 1674 63472
rect 1730 63416 1735 63472
rect 0 63414 1735 63416
rect 0 63384 800 63414
rect 1669 63411 1735 63414
rect 3233 63474 3299 63477
rect 3550 63474 3556 63476
rect 3233 63472 3556 63474
rect 3233 63416 3238 63472
rect 3294 63416 3556 63472
rect 3233 63414 3556 63416
rect 3233 63411 3299 63414
rect 3550 63412 3556 63414
rect 3620 63412 3626 63476
rect 10133 63338 10199 63341
rect 11200 63338 12000 63368
rect 10133 63336 12000 63338
rect 10133 63280 10138 63336
rect 10194 63280 12000 63336
rect 10133 63278 12000 63280
rect 10133 63275 10199 63278
rect 11200 63248 12000 63278
rect 4208 63136 4528 63137
rect 0 63066 800 63096
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 63071 4528 63072
rect 7472 63136 7792 63137
rect 7472 63072 7480 63136
rect 7544 63072 7560 63136
rect 7624 63072 7640 63136
rect 7704 63072 7720 63136
rect 7784 63072 7792 63136
rect 7472 63071 7792 63072
rect 1577 63066 1643 63069
rect 0 63064 1643 63066
rect 0 63008 1582 63064
rect 1638 63008 1643 63064
rect 0 63006 1643 63008
rect 0 62976 800 63006
rect 1577 63003 1643 63006
rect 1894 62868 1900 62932
rect 1964 62930 1970 62932
rect 2865 62930 2931 62933
rect 1964 62928 2931 62930
rect 1964 62872 2870 62928
rect 2926 62872 2931 62928
rect 1964 62870 2931 62872
rect 1964 62868 1970 62870
rect 2865 62867 2931 62870
rect 0 62658 800 62688
rect 2313 62658 2379 62661
rect 0 62656 2379 62658
rect 0 62600 2318 62656
rect 2374 62600 2379 62656
rect 0 62598 2379 62600
rect 0 62568 800 62598
rect 2313 62595 2379 62598
rect 2576 62592 2896 62593
rect 2576 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2576 62527 2896 62528
rect 5840 62592 6160 62593
rect 5840 62528 5848 62592
rect 5912 62528 5928 62592
rect 5992 62528 6008 62592
rect 6072 62528 6088 62592
rect 6152 62528 6160 62592
rect 5840 62527 6160 62528
rect 9104 62592 9424 62593
rect 9104 62528 9112 62592
rect 9176 62528 9192 62592
rect 9256 62528 9272 62592
rect 9336 62528 9352 62592
rect 9416 62528 9424 62592
rect 9104 62527 9424 62528
rect 10133 62522 10199 62525
rect 11200 62522 12000 62552
rect 10133 62520 12000 62522
rect 10133 62464 10138 62520
rect 10194 62464 12000 62520
rect 10133 62462 12000 62464
rect 10133 62459 10199 62462
rect 11200 62432 12000 62462
rect 1526 62188 1532 62252
rect 1596 62250 1602 62252
rect 1669 62250 1735 62253
rect 1596 62248 1735 62250
rect 1596 62192 1674 62248
rect 1730 62192 1735 62248
rect 1596 62190 1735 62192
rect 1596 62188 1602 62190
rect 1669 62187 1735 62190
rect 0 62114 800 62144
rect 1393 62114 1459 62117
rect 0 62112 1459 62114
rect 0 62056 1398 62112
rect 1454 62056 1459 62112
rect 0 62054 1459 62056
rect 0 62024 800 62054
rect 1393 62051 1459 62054
rect 4208 62048 4528 62049
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 61983 4528 61984
rect 7472 62048 7792 62049
rect 7472 61984 7480 62048
rect 7544 61984 7560 62048
rect 7624 61984 7640 62048
rect 7704 61984 7720 62048
rect 7784 61984 7792 62048
rect 7472 61983 7792 61984
rect 2681 61842 2747 61845
rect 3366 61842 3372 61844
rect 2681 61840 3372 61842
rect 2681 61784 2686 61840
rect 2742 61784 3372 61840
rect 2681 61782 3372 61784
rect 2681 61779 2747 61782
rect 3366 61780 3372 61782
rect 3436 61842 3442 61844
rect 3693 61842 3759 61845
rect 3436 61840 3759 61842
rect 3436 61784 3698 61840
rect 3754 61784 3759 61840
rect 3436 61782 3759 61784
rect 3436 61780 3442 61782
rect 3693 61779 3759 61782
rect 10133 61842 10199 61845
rect 11200 61842 12000 61872
rect 10133 61840 12000 61842
rect 10133 61784 10138 61840
rect 10194 61784 12000 61840
rect 10133 61782 12000 61784
rect 10133 61779 10199 61782
rect 11200 61752 12000 61782
rect 0 61706 800 61736
rect 3693 61706 3759 61709
rect 0 61704 3759 61706
rect 0 61648 3698 61704
rect 3754 61648 3759 61704
rect 0 61646 3759 61648
rect 0 61616 800 61646
rect 3693 61643 3759 61646
rect 2576 61504 2896 61505
rect 2576 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2576 61439 2896 61440
rect 5840 61504 6160 61505
rect 5840 61440 5848 61504
rect 5912 61440 5928 61504
rect 5992 61440 6008 61504
rect 6072 61440 6088 61504
rect 6152 61440 6160 61504
rect 5840 61439 6160 61440
rect 9104 61504 9424 61505
rect 9104 61440 9112 61504
rect 9176 61440 9192 61504
rect 9256 61440 9272 61504
rect 9336 61440 9352 61504
rect 9416 61440 9424 61504
rect 9104 61439 9424 61440
rect 1577 61432 1643 61437
rect 1577 61376 1582 61432
rect 1638 61376 1643 61432
rect 1577 61371 1643 61376
rect 3785 61434 3851 61437
rect 3969 61434 4035 61437
rect 3785 61432 4035 61434
rect 3785 61376 3790 61432
rect 3846 61376 3974 61432
rect 4030 61376 4035 61432
rect 3785 61374 4035 61376
rect 3785 61371 3851 61374
rect 3969 61371 4035 61374
rect 0 61298 800 61328
rect 1580 61298 1640 61371
rect 0 61238 1640 61298
rect 1761 61298 1827 61301
rect 2262 61298 2268 61300
rect 1761 61296 2268 61298
rect 1761 61240 1766 61296
rect 1822 61240 2268 61296
rect 1761 61238 2268 61240
rect 0 61208 800 61238
rect 1761 61235 1827 61238
rect 2262 61236 2268 61238
rect 2332 61236 2338 61300
rect 2078 61100 2084 61164
rect 2148 61162 2154 61164
rect 2148 61102 2514 61162
rect 2148 61100 2154 61102
rect 2454 61029 2514 61102
rect 1945 61026 2011 61029
rect 2078 61026 2084 61028
rect 1945 61024 2084 61026
rect 1945 60968 1950 61024
rect 2006 60968 2084 61024
rect 1945 60966 2084 60968
rect 1945 60963 2011 60966
rect 2078 60964 2084 60966
rect 2148 60964 2154 61028
rect 2454 61024 2563 61029
rect 2454 60968 2502 61024
rect 2558 60968 2563 61024
rect 2454 60966 2563 60968
rect 2497 60963 2563 60966
rect 3182 60964 3188 61028
rect 3252 61026 3258 61028
rect 3417 61026 3483 61029
rect 3252 61024 3483 61026
rect 3252 60968 3422 61024
rect 3478 60968 3483 61024
rect 3252 60966 3483 60968
rect 3252 60964 3258 60966
rect 3417 60963 3483 60966
rect 10133 61026 10199 61029
rect 11200 61026 12000 61056
rect 10133 61024 12000 61026
rect 10133 60968 10138 61024
rect 10194 60968 12000 61024
rect 10133 60966 12000 60968
rect 10133 60963 10199 60966
rect 4208 60960 4528 60961
rect 0 60890 800 60920
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 60895 4528 60896
rect 7472 60960 7792 60961
rect 7472 60896 7480 60960
rect 7544 60896 7560 60960
rect 7624 60896 7640 60960
rect 7704 60896 7720 60960
rect 7784 60896 7792 60960
rect 11200 60936 12000 60966
rect 7472 60895 7792 60896
rect 2773 60890 2839 60893
rect 0 60888 2839 60890
rect 0 60832 2778 60888
rect 2834 60832 2839 60888
rect 0 60830 2839 60832
rect 0 60800 800 60830
rect 2773 60827 2839 60830
rect 2998 60828 3004 60892
rect 3068 60890 3074 60892
rect 3233 60890 3299 60893
rect 3068 60888 3299 60890
rect 3068 60832 3238 60888
rect 3294 60832 3299 60888
rect 3068 60830 3299 60832
rect 3068 60828 3074 60830
rect 3233 60827 3299 60830
rect 2313 60754 2379 60757
rect 1166 60752 2379 60754
rect 1166 60696 2318 60752
rect 2374 60696 2379 60752
rect 1166 60694 2379 60696
rect 933 60618 999 60621
rect 1166 60618 1226 60694
rect 2313 60691 2379 60694
rect 2957 60754 3023 60757
rect 3233 60754 3299 60757
rect 2957 60752 3299 60754
rect 2957 60696 2962 60752
rect 3018 60696 3238 60752
rect 3294 60696 3299 60752
rect 2957 60694 3299 60696
rect 2957 60691 3023 60694
rect 3233 60691 3299 60694
rect 2957 60618 3023 60621
rect 933 60616 1226 60618
rect 933 60560 938 60616
rect 994 60560 1226 60616
rect 933 60558 1226 60560
rect 1350 60616 3023 60618
rect 1350 60560 2962 60616
rect 3018 60560 3023 60616
rect 1350 60558 3023 60560
rect 933 60555 999 60558
rect 0 60482 800 60512
rect 1350 60482 1410 60558
rect 2957 60555 3023 60558
rect 3734 60556 3740 60620
rect 3804 60618 3810 60620
rect 4061 60618 4127 60621
rect 3804 60616 4127 60618
rect 3804 60560 4066 60616
rect 4122 60560 4127 60616
rect 3804 60558 4127 60560
rect 3804 60556 3810 60558
rect 4061 60555 4127 60558
rect 0 60422 1410 60482
rect 0 60392 800 60422
rect 2998 60420 3004 60484
rect 3068 60482 3074 60484
rect 4061 60482 4127 60485
rect 3068 60480 4127 60482
rect 3068 60424 4066 60480
rect 4122 60424 4127 60480
rect 3068 60422 4127 60424
rect 3068 60420 3074 60422
rect 4061 60419 4127 60422
rect 2576 60416 2896 60417
rect 2576 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2576 60351 2896 60352
rect 5840 60416 6160 60417
rect 5840 60352 5848 60416
rect 5912 60352 5928 60416
rect 5992 60352 6008 60416
rect 6072 60352 6088 60416
rect 6152 60352 6160 60416
rect 5840 60351 6160 60352
rect 9104 60416 9424 60417
rect 9104 60352 9112 60416
rect 9176 60352 9192 60416
rect 9256 60352 9272 60416
rect 9336 60352 9352 60416
rect 9416 60352 9424 60416
rect 9104 60351 9424 60352
rect 3049 60346 3115 60349
rect 3366 60346 3372 60348
rect 3049 60344 3372 60346
rect 3049 60288 3054 60344
rect 3110 60288 3372 60344
rect 3049 60286 3372 60288
rect 3049 60283 3115 60286
rect 3366 60284 3372 60286
rect 3436 60284 3442 60348
rect 10133 60346 10199 60349
rect 11200 60346 12000 60376
rect 10133 60344 12000 60346
rect 10133 60288 10138 60344
rect 10194 60288 12000 60344
rect 10133 60286 12000 60288
rect 10133 60283 10199 60286
rect 11200 60256 12000 60286
rect 0 60074 800 60104
rect 2313 60074 2379 60077
rect 6177 60074 6243 60077
rect 0 60072 2379 60074
rect 0 60016 2318 60072
rect 2374 60016 2379 60072
rect 0 60014 2379 60016
rect 0 59984 800 60014
rect 2313 60011 2379 60014
rect 2454 60072 6243 60074
rect 2454 60016 6182 60072
rect 6238 60016 6243 60072
rect 2454 60014 6243 60016
rect 2313 59938 2379 59941
rect 2454 59938 2514 60014
rect 6177 60011 6243 60014
rect 2313 59936 2514 59938
rect 2313 59880 2318 59936
rect 2374 59880 2514 59936
rect 2313 59878 2514 59880
rect 2313 59875 2379 59878
rect 4208 59872 4528 59873
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 59807 4528 59808
rect 7472 59872 7792 59873
rect 7472 59808 7480 59872
rect 7544 59808 7560 59872
rect 7624 59808 7640 59872
rect 7704 59808 7720 59872
rect 7784 59808 7792 59872
rect 7472 59807 7792 59808
rect 0 59666 800 59696
rect 2773 59666 2839 59669
rect 0 59664 2839 59666
rect 0 59608 2778 59664
rect 2834 59608 2839 59664
rect 0 59606 2839 59608
rect 0 59576 800 59606
rect 2773 59603 2839 59606
rect 2129 59530 2195 59533
rect 2262 59530 2268 59532
rect 2129 59528 2268 59530
rect 2129 59472 2134 59528
rect 2190 59472 2268 59528
rect 2129 59470 2268 59472
rect 2129 59467 2195 59470
rect 2262 59468 2268 59470
rect 2332 59530 2338 59532
rect 2589 59530 2655 59533
rect 2332 59528 2655 59530
rect 2332 59472 2594 59528
rect 2650 59472 2655 59528
rect 2332 59470 2655 59472
rect 2332 59468 2338 59470
rect 2589 59467 2655 59470
rect 10133 59530 10199 59533
rect 11200 59530 12000 59560
rect 10133 59528 12000 59530
rect 10133 59472 10138 59528
rect 10194 59472 12000 59528
rect 10133 59470 12000 59472
rect 10133 59467 10199 59470
rect 11200 59440 12000 59470
rect 2576 59328 2896 59329
rect 2576 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2576 59263 2896 59264
rect 5840 59328 6160 59329
rect 5840 59264 5848 59328
rect 5912 59264 5928 59328
rect 5992 59264 6008 59328
rect 6072 59264 6088 59328
rect 6152 59264 6160 59328
rect 5840 59263 6160 59264
rect 9104 59328 9424 59329
rect 9104 59264 9112 59328
rect 9176 59264 9192 59328
rect 9256 59264 9272 59328
rect 9336 59264 9352 59328
rect 9416 59264 9424 59328
rect 9104 59263 9424 59264
rect 0 59122 800 59152
rect 1577 59122 1643 59125
rect 0 59120 1643 59122
rect 0 59064 1582 59120
rect 1638 59064 1643 59120
rect 0 59062 1643 59064
rect 0 59032 800 59062
rect 1577 59059 1643 59062
rect 1117 58986 1183 58989
rect 5073 58986 5139 58989
rect 1117 58984 5139 58986
rect 1117 58928 1122 58984
rect 1178 58928 5078 58984
rect 5134 58928 5139 58984
rect 1117 58926 5139 58928
rect 1117 58923 1183 58926
rect 5073 58923 5139 58926
rect 1117 58850 1183 58853
rect 2221 58850 2287 58853
rect 1117 58848 2287 58850
rect 1117 58792 1122 58848
rect 1178 58792 2226 58848
rect 2282 58792 2287 58848
rect 1117 58790 2287 58792
rect 1117 58787 1183 58790
rect 2221 58787 2287 58790
rect 4208 58784 4528 58785
rect 0 58714 800 58744
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 58719 4528 58720
rect 7472 58784 7792 58785
rect 7472 58720 7480 58784
rect 7544 58720 7560 58784
rect 7624 58720 7640 58784
rect 7704 58720 7720 58784
rect 7784 58720 7792 58784
rect 7472 58719 7792 58720
rect 3969 58714 4035 58717
rect 0 58712 4035 58714
rect 0 58656 3974 58712
rect 4030 58656 4035 58712
rect 0 58654 4035 58656
rect 0 58624 800 58654
rect 3969 58651 4035 58654
rect 10133 58714 10199 58717
rect 11200 58714 12000 58744
rect 10133 58712 12000 58714
rect 10133 58656 10138 58712
rect 10194 58656 12000 58712
rect 10133 58654 12000 58656
rect 10133 58651 10199 58654
rect 11200 58624 12000 58654
rect 2681 58578 2747 58581
rect 3550 58578 3556 58580
rect 2681 58576 3556 58578
rect 2681 58520 2686 58576
rect 2742 58520 3556 58576
rect 2681 58518 3556 58520
rect 2681 58515 2747 58518
rect 3550 58516 3556 58518
rect 3620 58516 3626 58580
rect 3509 58442 3575 58445
rect 1350 58440 3575 58442
rect 1350 58384 3514 58440
rect 3570 58384 3575 58440
rect 1350 58382 3575 58384
rect 0 58306 800 58336
rect 1350 58306 1410 58382
rect 3509 58379 3575 58382
rect 0 58246 1410 58306
rect 0 58216 800 58246
rect 2576 58240 2896 58241
rect 2576 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2576 58175 2896 58176
rect 5840 58240 6160 58241
rect 5840 58176 5848 58240
rect 5912 58176 5928 58240
rect 5992 58176 6008 58240
rect 6072 58176 6088 58240
rect 6152 58176 6160 58240
rect 5840 58175 6160 58176
rect 9104 58240 9424 58241
rect 9104 58176 9112 58240
rect 9176 58176 9192 58240
rect 9256 58176 9272 58240
rect 9336 58176 9352 58240
rect 9416 58176 9424 58240
rect 9104 58175 9424 58176
rect 9489 58034 9555 58037
rect 11200 58034 12000 58064
rect 9489 58032 12000 58034
rect 9489 57976 9494 58032
rect 9550 57976 12000 58032
rect 9489 57974 12000 57976
rect 9489 57971 9555 57974
rect 11200 57944 12000 57974
rect 0 57898 800 57928
rect 2589 57898 2655 57901
rect 0 57896 2655 57898
rect 0 57840 2594 57896
rect 2650 57840 2655 57896
rect 0 57838 2655 57840
rect 0 57808 800 57838
rect 2589 57835 2655 57838
rect 4208 57696 4528 57697
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 57631 4528 57632
rect 7472 57696 7792 57697
rect 7472 57632 7480 57696
rect 7544 57632 7560 57696
rect 7624 57632 7640 57696
rect 7704 57632 7720 57696
rect 7784 57632 7792 57696
rect 7472 57631 7792 57632
rect 2262 57564 2268 57628
rect 2332 57626 2338 57628
rect 2405 57626 2471 57629
rect 2332 57624 2471 57626
rect 2332 57568 2410 57624
rect 2466 57568 2471 57624
rect 2332 57566 2471 57568
rect 2332 57564 2338 57566
rect 2405 57563 2471 57566
rect 0 57490 800 57520
rect 1393 57490 1459 57493
rect 0 57488 1459 57490
rect 0 57432 1398 57488
rect 1454 57432 1459 57488
rect 0 57430 1459 57432
rect 0 57400 800 57430
rect 1393 57427 1459 57430
rect 1945 57490 2011 57493
rect 5574 57490 5580 57492
rect 1945 57488 5580 57490
rect 1945 57432 1950 57488
rect 2006 57432 5580 57488
rect 1945 57430 5580 57432
rect 1945 57427 2011 57430
rect 5574 57428 5580 57430
rect 5644 57428 5650 57492
rect 2262 57292 2268 57356
rect 2332 57354 2338 57356
rect 2681 57354 2747 57357
rect 2332 57352 2747 57354
rect 2332 57296 2686 57352
rect 2742 57296 2747 57352
rect 2332 57294 2747 57296
rect 2332 57292 2338 57294
rect 2681 57291 2747 57294
rect 9489 57218 9555 57221
rect 11200 57218 12000 57248
rect 9489 57216 12000 57218
rect 9489 57160 9494 57216
rect 9550 57160 12000 57216
rect 9489 57158 12000 57160
rect 9489 57155 9555 57158
rect 2576 57152 2896 57153
rect 0 57082 800 57112
rect 2576 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2576 57087 2896 57088
rect 5840 57152 6160 57153
rect 5840 57088 5848 57152
rect 5912 57088 5928 57152
rect 5992 57088 6008 57152
rect 6072 57088 6088 57152
rect 6152 57088 6160 57152
rect 5840 57087 6160 57088
rect 9104 57152 9424 57153
rect 9104 57088 9112 57152
rect 9176 57088 9192 57152
rect 9256 57088 9272 57152
rect 9336 57088 9352 57152
rect 9416 57088 9424 57152
rect 11200 57128 12000 57158
rect 9104 57087 9424 57088
rect 1577 57082 1643 57085
rect 0 57080 1643 57082
rect 0 57024 1582 57080
rect 1638 57024 1643 57080
rect 0 57022 1643 57024
rect 0 56992 800 57022
rect 1577 57019 1643 57022
rect 0 56674 800 56704
rect 1669 56674 1735 56677
rect 0 56672 1735 56674
rect 0 56616 1674 56672
rect 1730 56616 1735 56672
rect 0 56614 1735 56616
rect 0 56584 800 56614
rect 1669 56611 1735 56614
rect 4208 56608 4528 56609
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 56543 4528 56544
rect 7472 56608 7792 56609
rect 7472 56544 7480 56608
rect 7544 56544 7560 56608
rect 7624 56544 7640 56608
rect 7704 56544 7720 56608
rect 7784 56544 7792 56608
rect 7472 56543 7792 56544
rect 54 56340 60 56404
rect 124 56402 130 56404
rect 1117 56402 1183 56405
rect 124 56400 1183 56402
rect 124 56344 1122 56400
rect 1178 56344 1183 56400
rect 124 56342 1183 56344
rect 124 56340 130 56342
rect 1117 56339 1183 56342
rect 9305 56402 9371 56405
rect 11200 56402 12000 56432
rect 9305 56400 12000 56402
rect 9305 56344 9310 56400
rect 9366 56344 12000 56400
rect 9305 56342 12000 56344
rect 9305 56339 9371 56342
rect 11200 56312 12000 56342
rect 2681 56266 2747 56269
rect 1350 56264 2747 56266
rect 1350 56208 2686 56264
rect 2742 56208 2747 56264
rect 1350 56206 2747 56208
rect 0 56130 800 56160
rect 1350 56130 1410 56206
rect 2681 56203 2747 56206
rect 0 56070 1410 56130
rect 0 56040 800 56070
rect 2576 56064 2896 56065
rect 2576 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2576 55999 2896 56000
rect 5840 56064 6160 56065
rect 5840 56000 5848 56064
rect 5912 56000 5928 56064
rect 5992 56000 6008 56064
rect 6072 56000 6088 56064
rect 6152 56000 6160 56064
rect 5840 55999 6160 56000
rect 9104 56064 9424 56065
rect 9104 56000 9112 56064
rect 9176 56000 9192 56064
rect 9256 56000 9272 56064
rect 9336 56000 9352 56064
rect 9416 56000 9424 56064
rect 9104 55999 9424 56000
rect 3509 55858 3575 55861
rect 3374 55856 3575 55858
rect 3374 55800 3514 55856
rect 3570 55800 3575 55856
rect 3374 55798 3575 55800
rect 0 55722 800 55752
rect 2313 55722 2379 55725
rect 0 55720 2379 55722
rect 0 55664 2318 55720
rect 2374 55664 2379 55720
rect 0 55662 2379 55664
rect 0 55632 800 55662
rect 2313 55659 2379 55662
rect 2865 55722 2931 55725
rect 3374 55724 3434 55798
rect 3509 55795 3575 55798
rect 3366 55722 3372 55724
rect 2865 55720 3372 55722
rect 2865 55664 2870 55720
rect 2926 55664 3372 55720
rect 2865 55662 3372 55664
rect 2865 55659 2931 55662
rect 3366 55660 3372 55662
rect 3436 55660 3442 55724
rect 4153 55722 4219 55725
rect 4654 55722 4660 55724
rect 4153 55720 4660 55722
rect 4153 55664 4158 55720
rect 4214 55664 4660 55720
rect 4153 55662 4660 55664
rect 4153 55659 4219 55662
rect 4654 55660 4660 55662
rect 4724 55660 4730 55724
rect 10133 55722 10199 55725
rect 11200 55722 12000 55752
rect 10133 55720 12000 55722
rect 10133 55664 10138 55720
rect 10194 55664 12000 55720
rect 10133 55662 12000 55664
rect 10133 55659 10199 55662
rect 11200 55632 12000 55662
rect 4208 55520 4528 55521
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 55455 4528 55456
rect 7472 55520 7792 55521
rect 7472 55456 7480 55520
rect 7544 55456 7560 55520
rect 7624 55456 7640 55520
rect 7704 55456 7720 55520
rect 7784 55456 7792 55520
rect 7472 55455 7792 55456
rect 1158 55388 1164 55452
rect 1228 55450 1234 55452
rect 1577 55450 1643 55453
rect 1228 55448 1643 55450
rect 1228 55392 1582 55448
rect 1638 55392 1643 55448
rect 1228 55390 1643 55392
rect 1228 55388 1234 55390
rect 1577 55387 1643 55390
rect 1761 55450 1827 55453
rect 1761 55448 3112 55450
rect 1761 55392 1766 55448
rect 1822 55392 3112 55448
rect 1761 55390 3112 55392
rect 1761 55387 1827 55390
rect 0 55314 800 55344
rect 3052 55317 3112 55390
rect 2313 55314 2379 55317
rect 0 55312 2379 55314
rect 0 55256 2318 55312
rect 2374 55256 2379 55312
rect 0 55254 2379 55256
rect 0 55224 800 55254
rect 2313 55251 2379 55254
rect 3049 55312 3115 55317
rect 3049 55256 3054 55312
rect 3110 55256 3115 55312
rect 3049 55251 3115 55256
rect 974 55116 980 55180
rect 1044 55178 1050 55180
rect 1301 55178 1367 55181
rect 1044 55176 1367 55178
rect 1044 55120 1306 55176
rect 1362 55120 1367 55176
rect 1044 55118 1367 55120
rect 1044 55116 1050 55118
rect 1301 55115 1367 55118
rect 2078 55116 2084 55180
rect 2148 55178 2154 55180
rect 2998 55178 3004 55180
rect 2148 55118 3004 55178
rect 2148 55116 2154 55118
rect 2998 55116 3004 55118
rect 3068 55116 3074 55180
rect 4337 55178 4403 55181
rect 4654 55178 4660 55180
rect 4337 55176 4660 55178
rect 4337 55120 4342 55176
rect 4398 55120 4660 55176
rect 4337 55118 4660 55120
rect 4337 55115 4403 55118
rect 4654 55116 4660 55118
rect 4724 55116 4730 55180
rect 3509 55042 3575 55045
rect 3374 55040 3575 55042
rect 3374 54984 3514 55040
rect 3570 54984 3575 55040
rect 3374 54982 3575 54984
rect 2576 54976 2896 54977
rect 0 54906 800 54936
rect 2576 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2576 54911 2896 54912
rect 1158 54906 1164 54908
rect 0 54846 1164 54906
rect 0 54816 800 54846
rect 1158 54844 1164 54846
rect 1228 54844 1234 54908
rect 974 54708 980 54772
rect 1044 54770 1050 54772
rect 3374 54770 3434 54982
rect 3509 54979 3575 54982
rect 5840 54976 6160 54977
rect 5840 54912 5848 54976
rect 5912 54912 5928 54976
rect 5992 54912 6008 54976
rect 6072 54912 6088 54976
rect 6152 54912 6160 54976
rect 5840 54911 6160 54912
rect 9104 54976 9424 54977
rect 9104 54912 9112 54976
rect 9176 54912 9192 54976
rect 9256 54912 9272 54976
rect 9336 54912 9352 54976
rect 9416 54912 9424 54976
rect 9104 54911 9424 54912
rect 9581 54906 9647 54909
rect 11200 54906 12000 54936
rect 9581 54904 12000 54906
rect 9581 54848 9586 54904
rect 9642 54848 12000 54904
rect 9581 54846 12000 54848
rect 9581 54843 9647 54846
rect 11200 54816 12000 54846
rect 1044 54710 3434 54770
rect 1044 54708 1050 54710
rect 0 54498 800 54528
rect 2773 54498 2839 54501
rect 0 54496 2839 54498
rect 0 54440 2778 54496
rect 2834 54440 2839 54496
rect 0 54438 2839 54440
rect 0 54408 800 54438
rect 2773 54435 2839 54438
rect 4208 54432 4528 54433
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 54367 4528 54368
rect 7472 54432 7792 54433
rect 7472 54368 7480 54432
rect 7544 54368 7560 54432
rect 7624 54368 7640 54432
rect 7704 54368 7720 54432
rect 7784 54368 7792 54432
rect 7472 54367 7792 54368
rect 1761 54362 1827 54365
rect 2078 54362 2084 54364
rect 1761 54360 2084 54362
rect 1761 54304 1766 54360
rect 1822 54304 2084 54360
rect 1761 54302 2084 54304
rect 1761 54299 1827 54302
rect 2078 54300 2084 54302
rect 2148 54300 2154 54364
rect 0 54090 800 54120
rect 1485 54090 1551 54093
rect 0 54088 1551 54090
rect 0 54032 1490 54088
rect 1546 54032 1551 54088
rect 0 54030 1551 54032
rect 0 54000 800 54030
rect 1485 54027 1551 54030
rect 10041 54090 10107 54093
rect 11200 54090 12000 54120
rect 10041 54088 12000 54090
rect 10041 54032 10046 54088
rect 10102 54032 12000 54088
rect 10041 54030 12000 54032
rect 10041 54027 10107 54030
rect 11200 54000 12000 54030
rect 2576 53888 2896 53889
rect 2576 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2576 53823 2896 53824
rect 5840 53888 6160 53889
rect 5840 53824 5848 53888
rect 5912 53824 5928 53888
rect 5992 53824 6008 53888
rect 6072 53824 6088 53888
rect 6152 53824 6160 53888
rect 5840 53823 6160 53824
rect 9104 53888 9424 53889
rect 9104 53824 9112 53888
rect 9176 53824 9192 53888
rect 9256 53824 9272 53888
rect 9336 53824 9352 53888
rect 9416 53824 9424 53888
rect 9104 53823 9424 53824
rect 0 53682 800 53712
rect 2037 53682 2103 53685
rect 0 53680 2103 53682
rect 0 53624 2042 53680
rect 2098 53624 2103 53680
rect 0 53622 2103 53624
rect 0 53592 800 53622
rect 2037 53619 2103 53622
rect 3182 53484 3188 53548
rect 3252 53546 3258 53548
rect 4838 53546 4844 53548
rect 3252 53486 4844 53546
rect 3252 53484 3258 53486
rect 4838 53484 4844 53486
rect 4908 53484 4914 53548
rect 473 53410 539 53413
rect 3182 53410 3188 53412
rect 473 53408 3188 53410
rect 473 53352 478 53408
rect 534 53352 3188 53408
rect 473 53350 3188 53352
rect 473 53347 539 53350
rect 3182 53348 3188 53350
rect 3252 53348 3258 53412
rect 10041 53410 10107 53413
rect 11200 53410 12000 53440
rect 10041 53408 12000 53410
rect 10041 53352 10046 53408
rect 10102 53352 12000 53408
rect 10041 53350 12000 53352
rect 10041 53347 10107 53350
rect 4208 53344 4528 53345
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 53279 4528 53280
rect 7472 53344 7792 53345
rect 7472 53280 7480 53344
rect 7544 53280 7560 53344
rect 7624 53280 7640 53344
rect 7704 53280 7720 53344
rect 7784 53280 7792 53344
rect 11200 53320 12000 53350
rect 7472 53279 7792 53280
rect 0 53138 800 53168
rect 2313 53138 2379 53141
rect 0 53136 2379 53138
rect 0 53080 2318 53136
rect 2374 53080 2379 53136
rect 0 53078 2379 53080
rect 0 53048 800 53078
rect 2313 53075 2379 53078
rect 2589 53002 2655 53005
rect 2132 53000 2655 53002
rect 2132 52944 2594 53000
rect 2650 52944 2655 53000
rect 2132 52942 2655 52944
rect 0 52730 800 52760
rect 2132 52733 2192 52942
rect 2589 52939 2655 52942
rect 4654 52804 4660 52868
rect 4724 52866 4730 52868
rect 4797 52866 4863 52869
rect 4724 52864 4863 52866
rect 4724 52808 4802 52864
rect 4858 52808 4863 52864
rect 4724 52806 4863 52808
rect 4724 52804 4730 52806
rect 4797 52803 4863 52806
rect 2576 52800 2896 52801
rect 2576 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2576 52735 2896 52736
rect 5840 52800 6160 52801
rect 5840 52736 5848 52800
rect 5912 52736 5928 52800
rect 5992 52736 6008 52800
rect 6072 52736 6088 52800
rect 6152 52736 6160 52800
rect 5840 52735 6160 52736
rect 9104 52800 9424 52801
rect 9104 52736 9112 52800
rect 9176 52736 9192 52800
rect 9256 52736 9272 52800
rect 9336 52736 9352 52800
rect 9416 52736 9424 52800
rect 9104 52735 9424 52736
rect 1393 52730 1459 52733
rect 0 52728 1459 52730
rect 0 52672 1398 52728
rect 1454 52672 1459 52728
rect 0 52670 1459 52672
rect 0 52640 800 52670
rect 1393 52667 1459 52670
rect 2129 52728 2195 52733
rect 2129 52672 2134 52728
rect 2190 52672 2195 52728
rect 2129 52667 2195 52672
rect 3734 52668 3740 52732
rect 3804 52730 3810 52732
rect 4153 52730 4219 52733
rect 5349 52732 5415 52733
rect 5349 52730 5396 52732
rect 3804 52728 4219 52730
rect 3804 52672 4158 52728
rect 4214 52672 4219 52728
rect 3804 52670 4219 52672
rect 5304 52728 5396 52730
rect 5304 52672 5354 52728
rect 5304 52670 5396 52672
rect 3804 52668 3810 52670
rect 4153 52667 4219 52670
rect 5349 52668 5396 52670
rect 5460 52668 5466 52732
rect 5349 52667 5415 52668
rect 10041 52594 10107 52597
rect 11200 52594 12000 52624
rect 10041 52592 12000 52594
rect 10041 52536 10046 52592
rect 10102 52536 12000 52592
rect 10041 52534 12000 52536
rect 10041 52531 10107 52534
rect 11200 52504 12000 52534
rect 0 52322 800 52352
rect 1577 52322 1643 52325
rect 0 52320 1643 52322
rect 0 52264 1582 52320
rect 1638 52264 1643 52320
rect 0 52262 1643 52264
rect 0 52232 800 52262
rect 1577 52259 1643 52262
rect 4208 52256 4528 52257
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 52191 4528 52192
rect 7472 52256 7792 52257
rect 7472 52192 7480 52256
rect 7544 52192 7560 52256
rect 7624 52192 7640 52256
rect 7704 52192 7720 52256
rect 7784 52192 7792 52256
rect 7472 52191 7792 52192
rect 1577 52186 1643 52189
rect 1534 52184 1643 52186
rect 1534 52128 1582 52184
rect 1638 52128 1643 52184
rect 1534 52123 1643 52128
rect 5206 52124 5212 52188
rect 5276 52186 5282 52188
rect 5349 52186 5415 52189
rect 5276 52184 5415 52186
rect 5276 52128 5354 52184
rect 5410 52128 5415 52184
rect 5276 52126 5415 52128
rect 5276 52124 5282 52126
rect 5349 52123 5415 52126
rect 1534 52050 1594 52123
rect 798 51990 1594 52050
rect 798 51944 858 51990
rect 0 51854 858 51944
rect 2865 51914 2931 51917
rect 2865 51912 3066 51914
rect 2865 51856 2870 51912
rect 2926 51856 3066 51912
rect 2865 51854 3066 51856
rect 0 51824 800 51854
rect 2865 51851 2931 51854
rect 2576 51712 2896 51713
rect 2576 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2576 51647 2896 51648
rect 974 51580 980 51644
rect 1044 51642 1050 51644
rect 1301 51642 1367 51645
rect 1044 51640 1367 51642
rect 1044 51584 1306 51640
rect 1362 51584 1367 51640
rect 1044 51582 1367 51584
rect 1044 51580 1050 51582
rect 1301 51579 1367 51582
rect 0 51506 800 51536
rect 3006 51506 3066 51854
rect 10041 51778 10107 51781
rect 11200 51778 12000 51808
rect 10041 51776 12000 51778
rect 10041 51720 10046 51776
rect 10102 51720 12000 51776
rect 10041 51718 12000 51720
rect 10041 51715 10107 51718
rect 5840 51712 6160 51713
rect 5840 51648 5848 51712
rect 5912 51648 5928 51712
rect 5992 51648 6008 51712
rect 6072 51648 6088 51712
rect 6152 51648 6160 51712
rect 5840 51647 6160 51648
rect 9104 51712 9424 51713
rect 9104 51648 9112 51712
rect 9176 51648 9192 51712
rect 9256 51648 9272 51712
rect 9336 51648 9352 51712
rect 9416 51648 9424 51712
rect 11200 51688 12000 51718
rect 9104 51647 9424 51648
rect 3233 51642 3299 51645
rect 0 51446 3066 51506
rect 3190 51640 3299 51642
rect 3190 51584 3238 51640
rect 3294 51584 3299 51640
rect 3190 51579 3299 51584
rect 0 51416 800 51446
rect 1158 51308 1164 51372
rect 1228 51370 1234 51372
rect 1761 51370 1827 51373
rect 1228 51368 1827 51370
rect 1228 51312 1766 51368
rect 1822 51312 1827 51368
rect 1228 51310 1827 51312
rect 1228 51308 1234 51310
rect 1761 51307 1827 51310
rect 2078 51308 2084 51372
rect 2148 51370 2154 51372
rect 2148 51310 2514 51370
rect 2148 51308 2154 51310
rect 1301 51234 1367 51237
rect 1166 51232 1367 51234
rect 1166 51176 1306 51232
rect 1362 51176 1367 51232
rect 1166 51174 1367 51176
rect 0 51098 800 51128
rect 1166 51098 1226 51174
rect 1301 51171 1367 51174
rect 1761 51234 1827 51237
rect 2129 51234 2195 51237
rect 1761 51232 2195 51234
rect 1761 51176 1766 51232
rect 1822 51176 2134 51232
rect 2190 51176 2195 51232
rect 1761 51174 2195 51176
rect 1761 51171 1827 51174
rect 2129 51171 2195 51174
rect 1669 51098 1735 51101
rect 0 51038 1226 51098
rect 1534 51096 1735 51098
rect 1534 51040 1674 51096
rect 1730 51040 1735 51096
rect 1534 51038 1735 51040
rect 0 51008 800 51038
rect 974 50900 980 50964
rect 1044 50962 1050 50964
rect 1209 50962 1275 50965
rect 1393 50962 1459 50965
rect 1044 50960 1275 50962
rect 1044 50904 1214 50960
rect 1270 50904 1275 50960
rect 1044 50902 1275 50904
rect 1044 50900 1050 50902
rect 1209 50899 1275 50902
rect 1350 50960 1459 50962
rect 1350 50904 1398 50960
rect 1454 50904 1459 50960
rect 1350 50899 1459 50904
rect 974 50764 980 50828
rect 1044 50826 1050 50828
rect 1350 50826 1410 50899
rect 1044 50766 1410 50826
rect 1534 50826 1594 51038
rect 1669 51035 1735 51038
rect 2129 50826 2195 50829
rect 1534 50824 2195 50826
rect 1534 50768 2134 50824
rect 2190 50768 2195 50824
rect 1534 50766 2195 50768
rect 1044 50764 1050 50766
rect 2129 50763 2195 50766
rect 0 50690 800 50720
rect 1117 50690 1183 50693
rect 0 50688 1183 50690
rect 0 50632 1122 50688
rect 1178 50632 1183 50688
rect 0 50630 1183 50632
rect 0 50600 800 50630
rect 1117 50627 1183 50630
rect 105 50420 171 50421
rect 54 50356 60 50420
rect 124 50418 171 50420
rect 1669 50420 1735 50421
rect 124 50416 216 50418
rect 166 50360 216 50416
rect 124 50358 216 50360
rect 1669 50416 1716 50420
rect 1780 50418 1786 50420
rect 2454 50418 2514 51310
rect 3190 51234 3250 51579
rect 4613 51508 4679 51509
rect 4613 51506 4660 51508
rect 4568 51504 4660 51506
rect 4568 51448 4618 51504
rect 4568 51446 4660 51448
rect 4613 51444 4660 51446
rect 4724 51444 4730 51508
rect 4613 51443 4679 51444
rect 3366 51308 3372 51372
rect 3436 51370 3442 51372
rect 3601 51370 3667 51373
rect 3436 51368 3667 51370
rect 3436 51312 3606 51368
rect 3662 51312 3667 51368
rect 3436 51310 3667 51312
rect 3436 51308 3442 51310
rect 3601 51307 3667 51310
rect 3366 51234 3372 51236
rect 3190 51174 3372 51234
rect 3366 51172 3372 51174
rect 3436 51172 3442 51236
rect 4208 51168 4528 51169
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 51103 4528 51104
rect 7472 51168 7792 51169
rect 7472 51104 7480 51168
rect 7544 51104 7560 51168
rect 7624 51104 7640 51168
rect 7704 51104 7720 51168
rect 7784 51104 7792 51168
rect 7472 51103 7792 51104
rect 10041 51098 10107 51101
rect 11200 51098 12000 51128
rect 10041 51096 12000 51098
rect 5022 51028 5028 51092
rect 5092 51090 5098 51092
rect 5349 51090 5415 51093
rect 5092 51088 5415 51090
rect 5092 51032 5354 51088
rect 5410 51032 5415 51088
rect 10041 51040 10046 51096
rect 10102 51040 12000 51096
rect 10041 51038 12000 51040
rect 10041 51035 10107 51038
rect 5092 51030 5415 51032
rect 5092 51028 5098 51030
rect 5349 51027 5415 51030
rect 11200 51008 12000 51038
rect 3141 50962 3207 50965
rect 3366 50962 3372 50964
rect 3141 50960 3372 50962
rect 3141 50904 3146 50960
rect 3202 50904 3372 50960
rect 3141 50902 3372 50904
rect 3141 50899 3207 50902
rect 3366 50900 3372 50902
rect 3436 50900 3442 50964
rect 3550 50900 3556 50964
rect 3620 50962 3626 50964
rect 4061 50962 4127 50965
rect 3620 50960 4127 50962
rect 3620 50904 4066 50960
rect 4122 50904 4127 50960
rect 3620 50902 4127 50904
rect 3620 50900 3626 50902
rect 4061 50899 4127 50902
rect 4981 50962 5047 50965
rect 4981 50960 5090 50962
rect 4981 50904 4986 50960
rect 5042 50904 5090 50960
rect 4981 50899 5090 50904
rect 4613 50826 4679 50829
rect 5030 50826 5090 50899
rect 4613 50824 5090 50826
rect 4613 50768 4618 50824
rect 4674 50768 5090 50824
rect 4613 50766 5090 50768
rect 4613 50763 4679 50766
rect 5206 50764 5212 50828
rect 5276 50826 5282 50828
rect 5349 50826 5415 50829
rect 5276 50824 5415 50826
rect 5276 50768 5354 50824
rect 5410 50768 5415 50824
rect 5276 50766 5415 50768
rect 5276 50764 5282 50766
rect 5349 50763 5415 50766
rect 4654 50628 4660 50692
rect 4724 50690 4730 50692
rect 4797 50690 4863 50693
rect 4724 50688 4863 50690
rect 4724 50632 4802 50688
rect 4858 50632 4863 50688
rect 4724 50630 4863 50632
rect 4724 50628 4730 50630
rect 4797 50627 4863 50630
rect 5073 50690 5139 50693
rect 5390 50690 5396 50692
rect 5073 50688 5396 50690
rect 5073 50632 5078 50688
rect 5134 50632 5396 50688
rect 5073 50630 5396 50632
rect 5073 50627 5139 50630
rect 5390 50628 5396 50630
rect 5460 50628 5466 50692
rect 2576 50624 2896 50625
rect 2576 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2576 50559 2896 50560
rect 5840 50624 6160 50625
rect 5840 50560 5848 50624
rect 5912 50560 5928 50624
rect 5992 50560 6008 50624
rect 6072 50560 6088 50624
rect 6152 50560 6160 50624
rect 5840 50559 6160 50560
rect 9104 50624 9424 50625
rect 9104 50560 9112 50624
rect 9176 50560 9192 50624
rect 9256 50560 9272 50624
rect 9336 50560 9352 50624
rect 9416 50560 9424 50624
rect 9104 50559 9424 50560
rect 4654 50418 4660 50420
rect 1669 50360 1674 50416
rect 124 50356 171 50358
rect 105 50355 171 50356
rect 1669 50356 1716 50360
rect 1780 50358 1826 50418
rect 2454 50358 4660 50418
rect 1780 50356 1786 50358
rect 4654 50356 4660 50358
rect 4724 50356 4730 50420
rect 1669 50355 1735 50356
rect 1485 50280 1551 50285
rect 1485 50224 1490 50280
rect 1546 50224 1551 50280
rect 1485 50219 1551 50224
rect 1710 50220 1716 50284
rect 1780 50282 1786 50284
rect 4838 50282 4844 50284
rect 1780 50222 4844 50282
rect 1780 50220 1786 50222
rect 4838 50220 4844 50222
rect 4908 50220 4914 50284
rect 10041 50282 10107 50285
rect 11200 50282 12000 50312
rect 10041 50280 12000 50282
rect 10041 50224 10046 50280
rect 10102 50224 12000 50280
rect 10041 50222 12000 50224
rect 10041 50219 10107 50222
rect 0 50146 800 50176
rect 1488 50146 1548 50219
rect 11200 50192 12000 50222
rect 0 50086 1548 50146
rect 2957 50146 3023 50149
rect 3366 50146 3372 50148
rect 2957 50144 3372 50146
rect 2957 50088 2962 50144
rect 3018 50088 3372 50144
rect 2957 50086 3372 50088
rect 0 50056 800 50086
rect 2957 50083 3023 50086
rect 3366 50084 3372 50086
rect 3436 50084 3442 50148
rect 4208 50080 4528 50081
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 50015 4528 50016
rect 7472 50080 7792 50081
rect 7472 50016 7480 50080
rect 7544 50016 7560 50080
rect 7624 50016 7640 50080
rect 7704 50016 7720 50080
rect 7784 50016 7792 50080
rect 7472 50015 7792 50016
rect 3785 50012 3851 50013
rect 3734 50010 3740 50012
rect 3694 49950 3740 50010
rect 3804 50008 3851 50012
rect 3846 49952 3851 50008
rect 3734 49948 3740 49950
rect 3804 49948 3851 49952
rect 3785 49947 3851 49948
rect 1117 49874 1183 49877
rect 6545 49874 6611 49877
rect 1117 49872 6611 49874
rect 1117 49816 1122 49872
rect 1178 49816 6550 49872
rect 6606 49816 6611 49872
rect 1117 49814 6611 49816
rect 1117 49811 1183 49814
rect 6545 49811 6611 49814
rect 0 49738 800 49768
rect 2773 49738 2839 49741
rect 0 49736 2839 49738
rect 0 49680 2778 49736
rect 2834 49680 2839 49736
rect 0 49678 2839 49680
rect 0 49648 800 49678
rect 2773 49675 2839 49678
rect 3509 49600 3575 49605
rect 3509 49544 3514 49600
rect 3570 49544 3575 49600
rect 3509 49539 3575 49544
rect 2576 49536 2896 49537
rect 2576 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2576 49471 2896 49472
rect 0 49330 800 49360
rect 2497 49330 2563 49333
rect 0 49328 2563 49330
rect 0 49272 2502 49328
rect 2558 49272 2563 49328
rect 0 49270 2563 49272
rect 0 49240 800 49270
rect 2497 49267 2563 49270
rect 2773 49330 2839 49333
rect 3512 49330 3572 49539
rect 5840 49536 6160 49537
rect 5840 49472 5848 49536
rect 5912 49472 5928 49536
rect 5992 49472 6008 49536
rect 6072 49472 6088 49536
rect 6152 49472 6160 49536
rect 5840 49471 6160 49472
rect 9104 49536 9424 49537
rect 9104 49472 9112 49536
rect 9176 49472 9192 49536
rect 9256 49472 9272 49536
rect 9336 49472 9352 49536
rect 9416 49472 9424 49536
rect 9104 49471 9424 49472
rect 9581 49466 9647 49469
rect 11200 49466 12000 49496
rect 9581 49464 12000 49466
rect 9581 49408 9586 49464
rect 9642 49408 12000 49464
rect 9581 49406 12000 49408
rect 9581 49403 9647 49406
rect 11200 49376 12000 49406
rect 2773 49328 3572 49330
rect 2773 49272 2778 49328
rect 2834 49272 3572 49328
rect 2773 49270 3572 49272
rect 4521 49330 4587 49333
rect 5206 49330 5212 49332
rect 4521 49328 5212 49330
rect 4521 49272 4526 49328
rect 4582 49272 5212 49328
rect 4521 49270 5212 49272
rect 2773 49267 2839 49270
rect 4521 49267 4587 49270
rect 5206 49268 5212 49270
rect 5276 49268 5282 49332
rect 2262 49132 2268 49196
rect 2332 49194 2338 49196
rect 2589 49194 2655 49197
rect 2332 49192 2655 49194
rect 2332 49136 2594 49192
rect 2650 49136 2655 49192
rect 2332 49134 2655 49136
rect 2332 49132 2338 49134
rect 2589 49131 2655 49134
rect 2865 49194 2931 49197
rect 5390 49194 5396 49196
rect 2865 49192 5396 49194
rect 2865 49136 2870 49192
rect 2926 49136 5396 49192
rect 2865 49134 5396 49136
rect 2865 49131 2931 49134
rect 5390 49132 5396 49134
rect 5460 49132 5466 49196
rect 2497 49058 2563 49061
rect 3141 49058 3207 49061
rect 2497 49056 3207 49058
rect 2497 49000 2502 49056
rect 2558 49000 3146 49056
rect 3202 49000 3207 49056
rect 2497 48998 3207 49000
rect 2497 48995 2563 48998
rect 3141 48995 3207 48998
rect 4208 48992 4528 48993
rect 0 48922 800 48952
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 48927 4528 48928
rect 7472 48992 7792 48993
rect 7472 48928 7480 48992
rect 7544 48928 7560 48992
rect 7624 48928 7640 48992
rect 7704 48928 7720 48992
rect 7784 48928 7792 48992
rect 7472 48927 7792 48928
rect 2313 48922 2379 48925
rect 0 48920 2379 48922
rect 0 48864 2318 48920
rect 2374 48864 2379 48920
rect 0 48862 2379 48864
rect 0 48832 800 48862
rect 2313 48859 2379 48862
rect 3325 48786 3391 48789
rect 3190 48784 3391 48786
rect 3190 48728 3330 48784
rect 3386 48728 3391 48784
rect 3190 48726 3391 48728
rect 2957 48648 3023 48653
rect 2957 48592 2962 48648
rect 3018 48592 3023 48648
rect 2957 48587 3023 48592
rect 0 48514 800 48544
rect 1393 48514 1459 48517
rect 0 48512 1459 48514
rect 0 48456 1398 48512
rect 1454 48456 1459 48512
rect 0 48454 1459 48456
rect 0 48424 800 48454
rect 1393 48451 1459 48454
rect 2576 48448 2896 48449
rect 2576 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2576 48383 2896 48384
rect 1117 48380 1183 48381
rect 1117 48376 1164 48380
rect 1228 48378 1234 48380
rect 1117 48320 1122 48376
rect 1117 48316 1164 48320
rect 1228 48318 1274 48378
rect 1228 48316 1234 48318
rect 1117 48315 1183 48316
rect 1761 48242 1827 48245
rect 1894 48242 1900 48244
rect 1761 48240 1900 48242
rect 1761 48184 1766 48240
rect 1822 48184 1900 48240
rect 1761 48182 1900 48184
rect 1761 48179 1827 48182
rect 1894 48180 1900 48182
rect 1964 48180 1970 48244
rect 2405 48240 2471 48245
rect 2405 48184 2410 48240
rect 2466 48184 2471 48240
rect 2405 48179 2471 48184
rect 2773 48242 2839 48245
rect 2960 48242 3020 48587
rect 2773 48240 3020 48242
rect 2773 48184 2778 48240
rect 2834 48184 3020 48240
rect 2773 48182 3020 48184
rect 2773 48179 2839 48182
rect 0 48106 800 48136
rect 1577 48106 1643 48109
rect 0 48104 1643 48106
rect 0 48048 1582 48104
rect 1638 48048 1643 48104
rect 0 48046 1643 48048
rect 0 48016 800 48046
rect 1577 48043 1643 48046
rect 1894 48044 1900 48108
rect 1964 48106 1970 48108
rect 2408 48106 2468 48179
rect 1964 48046 2468 48106
rect 3190 48106 3250 48726
rect 3325 48723 3391 48726
rect 10041 48786 10107 48789
rect 11200 48786 12000 48816
rect 10041 48784 12000 48786
rect 10041 48728 10046 48784
rect 10102 48728 12000 48784
rect 10041 48726 12000 48728
rect 10041 48723 10107 48726
rect 11200 48696 12000 48726
rect 4521 48514 4587 48517
rect 5574 48514 5580 48516
rect 4521 48512 5580 48514
rect 4521 48456 4526 48512
rect 4582 48456 5580 48512
rect 4521 48454 5580 48456
rect 4521 48451 4587 48454
rect 5574 48452 5580 48454
rect 5644 48452 5650 48516
rect 5840 48448 6160 48449
rect 5840 48384 5848 48448
rect 5912 48384 5928 48448
rect 5992 48384 6008 48448
rect 6072 48384 6088 48448
rect 6152 48384 6160 48448
rect 5840 48383 6160 48384
rect 9104 48448 9424 48449
rect 9104 48384 9112 48448
rect 9176 48384 9192 48448
rect 9256 48384 9272 48448
rect 9336 48384 9352 48448
rect 9416 48384 9424 48448
rect 9104 48383 9424 48384
rect 3785 48244 3851 48245
rect 3734 48180 3740 48244
rect 3804 48242 3851 48244
rect 3804 48240 3896 48242
rect 3846 48184 3896 48240
rect 3804 48182 3896 48184
rect 3804 48180 3851 48182
rect 3785 48179 3851 48180
rect 3325 48106 3391 48109
rect 4521 48106 4587 48109
rect 3190 48104 3391 48106
rect 3190 48048 3330 48104
rect 3386 48048 3391 48104
rect 3190 48046 3391 48048
rect 1964 48044 1970 48046
rect 3325 48043 3391 48046
rect 3972 48104 4587 48106
rect 3972 48048 4526 48104
rect 4582 48048 4587 48104
rect 3972 48046 4587 48048
rect 2262 47908 2268 47972
rect 2332 47970 2338 47972
rect 2405 47970 2471 47973
rect 3972 47970 4032 48046
rect 4521 48043 4587 48046
rect 2332 47968 4032 47970
rect 2332 47912 2410 47968
rect 2466 47912 4032 47968
rect 2332 47910 4032 47912
rect 10041 47970 10107 47973
rect 11200 47970 12000 48000
rect 10041 47968 12000 47970
rect 10041 47912 10046 47968
rect 10102 47912 12000 47968
rect 10041 47910 12000 47912
rect 2332 47908 2338 47910
rect 2405 47907 2471 47910
rect 10041 47907 10107 47910
rect 4208 47904 4528 47905
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 47839 4528 47840
rect 7472 47904 7792 47905
rect 7472 47840 7480 47904
rect 7544 47840 7560 47904
rect 7624 47840 7640 47904
rect 7704 47840 7720 47904
rect 7784 47840 7792 47904
rect 11200 47880 12000 47910
rect 7472 47839 7792 47840
rect 2400 47772 2406 47836
rect 2470 47834 2476 47836
rect 2681 47834 2747 47837
rect 2470 47832 2747 47834
rect 2470 47776 2686 47832
rect 2742 47776 2747 47832
rect 2470 47774 2747 47776
rect 2470 47772 2476 47774
rect 2681 47771 2747 47774
rect 3509 47834 3575 47837
rect 3734 47834 3740 47836
rect 3509 47832 3740 47834
rect 3509 47776 3514 47832
rect 3570 47776 3740 47832
rect 3509 47774 3740 47776
rect 3509 47771 3575 47774
rect 3734 47772 3740 47774
rect 3804 47772 3810 47836
rect 0 47698 800 47728
rect 1577 47698 1643 47701
rect 0 47696 1643 47698
rect 0 47640 1582 47696
rect 1638 47640 1643 47696
rect 0 47638 1643 47640
rect 0 47608 800 47638
rect 1577 47635 1643 47638
rect 3141 47698 3207 47701
rect 3141 47696 3250 47698
rect 3141 47640 3146 47696
rect 3202 47640 3250 47696
rect 3141 47635 3250 47640
rect 238 47364 244 47428
rect 308 47426 314 47428
rect 1393 47426 1459 47429
rect 308 47424 1459 47426
rect 308 47368 1398 47424
rect 1454 47368 1459 47424
rect 308 47366 1459 47368
rect 308 47364 314 47366
rect 1393 47363 1459 47366
rect 2576 47360 2896 47361
rect 2576 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2576 47295 2896 47296
rect 3190 47290 3250 47635
rect 4613 47562 4679 47565
rect 6310 47562 6316 47564
rect 4613 47560 6316 47562
rect 4613 47504 4618 47560
rect 4674 47504 6316 47560
rect 4613 47502 6316 47504
rect 4613 47499 4679 47502
rect 6310 47500 6316 47502
rect 6380 47500 6386 47564
rect 5840 47360 6160 47361
rect 5840 47296 5848 47360
rect 5912 47296 5928 47360
rect 5992 47296 6008 47360
rect 6072 47296 6088 47360
rect 6152 47296 6160 47360
rect 5840 47295 6160 47296
rect 9104 47360 9424 47361
rect 9104 47296 9112 47360
rect 9176 47296 9192 47360
rect 9256 47296 9272 47360
rect 9336 47296 9352 47360
rect 9416 47296 9424 47360
rect 9104 47295 9424 47296
rect 3325 47290 3391 47293
rect 3190 47288 3391 47290
rect 3190 47232 3330 47288
rect 3386 47232 3391 47288
rect 3190 47230 3391 47232
rect 3325 47227 3391 47230
rect 0 47154 800 47184
rect 3693 47154 3759 47157
rect 0 47152 3759 47154
rect 0 47096 3698 47152
rect 3754 47096 3759 47152
rect 0 47094 3759 47096
rect 0 47064 800 47094
rect 3693 47091 3759 47094
rect 3877 47154 3943 47157
rect 5574 47154 5580 47156
rect 3877 47152 5580 47154
rect 3877 47096 3882 47152
rect 3938 47096 5580 47152
rect 3877 47094 5580 47096
rect 3877 47091 3943 47094
rect 5574 47092 5580 47094
rect 5644 47092 5650 47156
rect 10041 47154 10107 47157
rect 11200 47154 12000 47184
rect 10041 47152 12000 47154
rect 10041 47096 10046 47152
rect 10102 47096 12000 47152
rect 10041 47094 12000 47096
rect 10041 47091 10107 47094
rect 11200 47064 12000 47094
rect 4521 47018 4587 47021
rect 4838 47018 4844 47020
rect 4521 47016 4844 47018
rect 4521 46960 4526 47016
rect 4582 46960 4844 47016
rect 4521 46958 4844 46960
rect 4521 46955 4587 46958
rect 4838 46956 4844 46958
rect 4908 46956 4914 47020
rect 1526 46820 1532 46884
rect 1596 46882 1602 46884
rect 1669 46882 1735 46885
rect 1596 46880 1735 46882
rect 1596 46824 1674 46880
rect 1730 46824 1735 46880
rect 1596 46822 1735 46824
rect 1596 46820 1602 46822
rect 1669 46819 1735 46822
rect 4208 46816 4528 46817
rect 0 46746 800 46776
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 7472 46816 7792 46817
rect 7472 46752 7480 46816
rect 7544 46752 7560 46816
rect 7624 46752 7640 46816
rect 7704 46752 7720 46816
rect 7784 46752 7792 46816
rect 7472 46751 7792 46752
rect 3969 46746 4035 46749
rect 0 46744 4035 46746
rect 0 46688 3974 46744
rect 4030 46688 4035 46744
rect 0 46686 4035 46688
rect 0 46656 800 46686
rect 3969 46683 4035 46686
rect 1393 46610 1459 46613
rect 1526 46610 1532 46612
rect 1393 46608 1532 46610
rect 105 46578 171 46579
rect 54 46514 60 46578
rect 124 46576 171 46578
rect 124 46574 216 46576
rect 166 46518 216 46574
rect 1393 46552 1398 46608
rect 1454 46552 1532 46608
rect 1393 46550 1532 46552
rect 1393 46547 1459 46550
rect 1526 46548 1532 46550
rect 1596 46548 1602 46612
rect 3693 46610 3759 46613
rect 8334 46610 8340 46612
rect 3693 46608 8340 46610
rect 3693 46552 3698 46608
rect 3754 46552 8340 46608
rect 3693 46550 8340 46552
rect 3693 46547 3759 46550
rect 8334 46548 8340 46550
rect 8404 46548 8410 46612
rect 124 46516 216 46518
rect 124 46514 171 46516
rect 105 46513 171 46514
rect 3877 46474 3943 46477
rect 1350 46472 3943 46474
rect 1350 46416 3882 46472
rect 3938 46416 3943 46472
rect 1350 46414 3943 46416
rect 0 46338 800 46368
rect 1350 46338 1410 46414
rect 3877 46411 3943 46414
rect 5022 46412 5028 46476
rect 5092 46474 5098 46476
rect 6494 46474 6500 46476
rect 5092 46414 6500 46474
rect 5092 46412 5098 46414
rect 6494 46412 6500 46414
rect 6564 46412 6570 46476
rect 10041 46474 10107 46477
rect 11200 46474 12000 46504
rect 10041 46472 12000 46474
rect 10041 46416 10046 46472
rect 10102 46416 12000 46472
rect 10041 46414 12000 46416
rect 10041 46411 10107 46414
rect 11200 46384 12000 46414
rect 0 46278 1410 46338
rect 0 46248 800 46278
rect 2576 46272 2896 46273
rect 2576 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2576 46207 2896 46208
rect 5840 46272 6160 46273
rect 5840 46208 5848 46272
rect 5912 46208 5928 46272
rect 5992 46208 6008 46272
rect 6072 46208 6088 46272
rect 6152 46208 6160 46272
rect 5840 46207 6160 46208
rect 9104 46272 9424 46273
rect 9104 46208 9112 46272
rect 9176 46208 9192 46272
rect 9256 46208 9272 46272
rect 9336 46208 9352 46272
rect 9416 46208 9424 46272
rect 9104 46207 9424 46208
rect 2681 46066 2747 46069
rect 5022 46066 5028 46068
rect 2681 46064 5028 46066
rect 2681 46008 2686 46064
rect 2742 46008 5028 46064
rect 2681 46006 5028 46008
rect 2681 46003 2747 46006
rect 5022 46004 5028 46006
rect 5092 46004 5098 46068
rect 0 45930 800 45960
rect 2865 45930 2931 45933
rect 0 45928 2931 45930
rect 0 45872 2870 45928
rect 2926 45872 2931 45928
rect 0 45870 2931 45872
rect 0 45840 800 45870
rect 2865 45867 2931 45870
rect 2998 45794 3004 45796
rect 2868 45734 3004 45794
rect 2868 45661 2928 45734
rect 2998 45732 3004 45734
rect 3068 45732 3074 45796
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 7472 45728 7792 45729
rect 7472 45664 7480 45728
rect 7544 45664 7560 45728
rect 7624 45664 7640 45728
rect 7704 45664 7720 45728
rect 7784 45664 7792 45728
rect 7472 45663 7792 45664
rect 1393 45658 1459 45661
rect 2400 45658 2406 45660
rect 1393 45656 2406 45658
rect 1393 45600 1398 45656
rect 1454 45600 2406 45656
rect 1393 45598 2406 45600
rect 1393 45595 1459 45598
rect 2400 45596 2406 45598
rect 2470 45596 2476 45660
rect 2865 45656 2931 45661
rect 2865 45600 2870 45656
rect 2926 45600 2931 45656
rect 2865 45595 2931 45600
rect 2998 45596 3004 45660
rect 3068 45658 3074 45660
rect 3785 45658 3851 45661
rect 3068 45656 3851 45658
rect 3068 45600 3790 45656
rect 3846 45600 3851 45656
rect 3068 45598 3851 45600
rect 3068 45596 3074 45598
rect 3785 45595 3851 45598
rect 4654 45596 4660 45660
rect 4724 45658 4730 45660
rect 5533 45658 5599 45661
rect 4724 45656 5599 45658
rect 4724 45600 5538 45656
rect 5594 45600 5599 45656
rect 4724 45598 5599 45600
rect 4724 45596 4730 45598
rect 5533 45595 5599 45598
rect 10041 45658 10107 45661
rect 11200 45658 12000 45688
rect 10041 45656 12000 45658
rect 10041 45600 10046 45656
rect 10102 45600 12000 45656
rect 10041 45598 12000 45600
rect 10041 45595 10107 45598
rect 11200 45568 12000 45598
rect 0 45522 800 45552
rect 3969 45522 4035 45525
rect 0 45520 4035 45522
rect 0 45464 3974 45520
rect 4030 45464 4035 45520
rect 0 45462 4035 45464
rect 0 45432 800 45462
rect 3969 45459 4035 45462
rect 1342 45324 1348 45388
rect 1412 45386 1418 45388
rect 1485 45386 1551 45389
rect 1412 45384 1551 45386
rect 1412 45328 1490 45384
rect 1546 45328 1551 45384
rect 1412 45326 1551 45328
rect 1412 45324 1418 45326
rect 1485 45323 1551 45326
rect 2400 45324 2406 45388
rect 2470 45386 2476 45388
rect 3182 45386 3188 45388
rect 2470 45326 3188 45386
rect 2470 45324 2476 45326
rect 3182 45324 3188 45326
rect 3252 45324 3258 45388
rect 2576 45184 2896 45185
rect 0 45114 800 45144
rect 2576 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2576 45119 2896 45120
rect 5840 45184 6160 45185
rect 5840 45120 5848 45184
rect 5912 45120 5928 45184
rect 5992 45120 6008 45184
rect 6072 45120 6088 45184
rect 6152 45120 6160 45184
rect 5840 45119 6160 45120
rect 9104 45184 9424 45185
rect 9104 45120 9112 45184
rect 9176 45120 9192 45184
rect 9256 45120 9272 45184
rect 9336 45120 9352 45184
rect 9416 45120 9424 45184
rect 9104 45119 9424 45120
rect 1577 45114 1643 45117
rect 0 45112 1643 45114
rect 0 45056 1582 45112
rect 1638 45056 1643 45112
rect 0 45054 1643 45056
rect 0 45024 800 45054
rect 1577 45051 1643 45054
rect 10041 44842 10107 44845
rect 11200 44842 12000 44872
rect 10041 44840 12000 44842
rect 10041 44784 10046 44840
rect 10102 44784 12000 44840
rect 10041 44782 12000 44784
rect 10041 44779 10107 44782
rect 11200 44752 12000 44782
rect 0 44706 800 44736
rect 1577 44706 1643 44709
rect 0 44704 1643 44706
rect 0 44648 1582 44704
rect 1638 44648 1643 44704
rect 0 44646 1643 44648
rect 0 44616 800 44646
rect 1577 44643 1643 44646
rect 3366 44644 3372 44708
rect 3436 44644 3442 44708
rect 289 44434 355 44437
rect 3374 44436 3434 44644
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 7472 44640 7792 44641
rect 7472 44576 7480 44640
rect 7544 44576 7560 44640
rect 7624 44576 7640 44640
rect 7704 44576 7720 44640
rect 7784 44576 7792 44640
rect 7472 44575 7792 44576
rect 422 44434 428 44436
rect 289 44432 428 44434
rect 289 44376 294 44432
rect 350 44376 428 44432
rect 289 44374 428 44376
rect 289 44371 355 44374
rect 422 44372 428 44374
rect 492 44372 498 44436
rect 606 44372 612 44436
rect 676 44434 682 44436
rect 974 44434 980 44436
rect 676 44374 980 44434
rect 676 44372 682 44374
rect 974 44372 980 44374
rect 1044 44372 1050 44436
rect 3366 44372 3372 44436
rect 3436 44372 3442 44436
rect 1158 44236 1164 44300
rect 1228 44298 1234 44300
rect 1393 44298 1459 44301
rect 1228 44296 1459 44298
rect 1228 44240 1398 44296
rect 1454 44240 1459 44296
rect 1228 44238 1459 44240
rect 1228 44236 1234 44238
rect 1393 44235 1459 44238
rect 0 44162 800 44192
rect 1577 44162 1643 44165
rect 0 44160 1643 44162
rect 0 44104 1582 44160
rect 1638 44104 1643 44160
rect 0 44102 1643 44104
rect 0 44072 800 44102
rect 1577 44099 1643 44102
rect 10041 44162 10107 44165
rect 11200 44162 12000 44192
rect 10041 44160 12000 44162
rect 10041 44104 10046 44160
rect 10102 44104 12000 44160
rect 10041 44102 12000 44104
rect 10041 44099 10107 44102
rect 2576 44096 2896 44097
rect 2576 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2576 44031 2896 44032
rect 5840 44096 6160 44097
rect 5840 44032 5848 44096
rect 5912 44032 5928 44096
rect 5992 44032 6008 44096
rect 6072 44032 6088 44096
rect 6152 44032 6160 44096
rect 5840 44031 6160 44032
rect 9104 44096 9424 44097
rect 9104 44032 9112 44096
rect 9176 44032 9192 44096
rect 9256 44032 9272 44096
rect 9336 44032 9352 44096
rect 9416 44032 9424 44096
rect 11200 44072 12000 44102
rect 9104 44031 9424 44032
rect 2078 43828 2084 43892
rect 2148 43890 2154 43892
rect 2681 43890 2747 43893
rect 2148 43888 2747 43890
rect 2148 43832 2686 43888
rect 2742 43832 2747 43888
rect 2148 43830 2747 43832
rect 2148 43828 2154 43830
rect 2681 43827 2747 43830
rect 3877 43890 3943 43893
rect 3877 43888 3986 43890
rect 3877 43832 3882 43888
rect 3938 43832 3986 43888
rect 3877 43827 3986 43832
rect 0 43754 800 43784
rect 0 43694 1456 43754
rect 0 43664 800 43694
rect 1396 43618 1456 43694
rect 1526 43692 1532 43756
rect 1596 43754 1602 43756
rect 2078 43754 2084 43756
rect 1596 43694 2084 43754
rect 1596 43692 1602 43694
rect 2078 43692 2084 43694
rect 2148 43692 2154 43756
rect 3417 43618 3483 43621
rect 1396 43616 3483 43618
rect 1396 43560 3422 43616
rect 3478 43560 3483 43616
rect 1396 43558 3483 43560
rect 3417 43555 3483 43558
rect 1526 43420 1532 43484
rect 1596 43482 1602 43484
rect 3049 43482 3115 43485
rect 1596 43480 3115 43482
rect 1596 43424 3054 43480
rect 3110 43424 3115 43480
rect 1596 43422 3115 43424
rect 1596 43420 1602 43422
rect 3049 43419 3115 43422
rect 0 43346 800 43376
rect 3785 43346 3851 43349
rect 0 43344 3851 43346
rect 0 43288 3790 43344
rect 3846 43288 3851 43344
rect 0 43286 3851 43288
rect 3926 43346 3986 43827
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 7472 43552 7792 43553
rect 7472 43488 7480 43552
rect 7544 43488 7560 43552
rect 7624 43488 7640 43552
rect 7704 43488 7720 43552
rect 7784 43488 7792 43552
rect 7472 43487 7792 43488
rect 4153 43346 4219 43349
rect 3926 43344 4219 43346
rect 3926 43288 4158 43344
rect 4214 43288 4219 43344
rect 3926 43286 4219 43288
rect 0 43256 800 43286
rect 3785 43283 3851 43286
rect 4153 43283 4219 43286
rect 10041 43346 10107 43349
rect 11200 43346 12000 43376
rect 10041 43344 12000 43346
rect 10041 43288 10046 43344
rect 10102 43288 12000 43344
rect 10041 43286 12000 43288
rect 10041 43283 10107 43286
rect 11200 43256 12000 43286
rect 3141 43210 3207 43213
rect 1350 43208 3207 43210
rect 1350 43152 3146 43208
rect 3202 43152 3207 43208
rect 1350 43150 3207 43152
rect 0 42938 800 42968
rect 1350 42938 1410 43150
rect 3141 43147 3207 43150
rect 3550 43148 3556 43212
rect 3620 43210 3626 43212
rect 3969 43210 4035 43213
rect 3620 43208 4035 43210
rect 3620 43152 3974 43208
rect 4030 43152 4035 43208
rect 3620 43150 4035 43152
rect 3620 43148 3626 43150
rect 3969 43147 4035 43150
rect 1485 43074 1551 43077
rect 1894 43074 1900 43076
rect 1485 43072 1900 43074
rect 1485 43016 1490 43072
rect 1546 43016 1900 43072
rect 1485 43014 1900 43016
rect 1485 43011 1551 43014
rect 1894 43012 1900 43014
rect 1964 43012 1970 43076
rect 3182 43074 3188 43076
rect 3052 43014 3188 43074
rect 2576 43008 2896 43009
rect 2576 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2576 42943 2896 42944
rect 1945 42940 2011 42941
rect 0 42878 1410 42938
rect 0 42848 800 42878
rect 1894 42876 1900 42940
rect 1964 42938 2011 42940
rect 1964 42936 2056 42938
rect 2006 42880 2056 42936
rect 1964 42878 2056 42880
rect 1964 42876 2011 42878
rect 1945 42875 2011 42876
rect 1301 42804 1367 42805
rect 1301 42800 1348 42804
rect 1412 42802 1418 42804
rect 1301 42744 1306 42800
rect 1301 42740 1348 42744
rect 1412 42742 1458 42802
rect 1412 42740 1418 42742
rect 1710 42740 1716 42804
rect 1780 42802 1786 42804
rect 1945 42802 2011 42805
rect 1780 42800 2011 42802
rect 1780 42744 1950 42800
rect 2006 42744 2011 42800
rect 1780 42742 2011 42744
rect 1780 42740 1786 42742
rect 1301 42739 1367 42740
rect 1945 42739 2011 42742
rect 2773 42802 2839 42805
rect 3052 42802 3112 43014
rect 3182 43012 3188 43014
rect 3252 43012 3258 43076
rect 5840 43008 6160 43009
rect 5840 42944 5848 43008
rect 5912 42944 5928 43008
rect 5992 42944 6008 43008
rect 6072 42944 6088 43008
rect 6152 42944 6160 43008
rect 5840 42943 6160 42944
rect 9104 43008 9424 43009
rect 9104 42944 9112 43008
rect 9176 42944 9192 43008
rect 9256 42944 9272 43008
rect 9336 42944 9352 43008
rect 9416 42944 9424 43008
rect 9104 42943 9424 42944
rect 3182 42876 3188 42940
rect 3252 42938 3258 42940
rect 3785 42938 3851 42941
rect 3252 42936 3851 42938
rect 3252 42880 3790 42936
rect 3846 42880 3851 42936
rect 3252 42878 3851 42880
rect 3252 42876 3258 42878
rect 3785 42875 3851 42878
rect 2773 42800 3112 42802
rect 2773 42744 2778 42800
rect 2834 42744 3112 42800
rect 2773 42742 3112 42744
rect 3785 42802 3851 42805
rect 3918 42802 3924 42804
rect 3785 42800 3924 42802
rect 3785 42744 3790 42800
rect 3846 42744 3924 42800
rect 3785 42742 3924 42744
rect 2773 42739 2839 42742
rect 3785 42739 3851 42742
rect 3918 42740 3924 42742
rect 3988 42740 3994 42804
rect 1342 42604 1348 42668
rect 1412 42666 1418 42668
rect 2078 42666 2084 42668
rect 1412 42606 2084 42666
rect 1412 42604 1418 42606
rect 2078 42604 2084 42606
rect 2148 42604 2154 42668
rect 0 42530 800 42560
rect 3969 42530 4035 42533
rect 0 42528 4035 42530
rect 0 42472 3974 42528
rect 4030 42472 4035 42528
rect 0 42470 4035 42472
rect 0 42440 800 42470
rect 3969 42467 4035 42470
rect 10041 42530 10107 42533
rect 11200 42530 12000 42560
rect 10041 42528 12000 42530
rect 10041 42472 10046 42528
rect 10102 42472 12000 42528
rect 10041 42470 12000 42472
rect 10041 42467 10107 42470
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 7472 42464 7792 42465
rect 7472 42400 7480 42464
rect 7544 42400 7560 42464
rect 7624 42400 7640 42464
rect 7704 42400 7720 42464
rect 7784 42400 7792 42464
rect 11200 42440 12000 42470
rect 7472 42399 7792 42400
rect 1761 42396 1827 42397
rect 1710 42394 1716 42396
rect 1670 42334 1716 42394
rect 1780 42392 1827 42396
rect 1822 42336 1827 42392
rect 1710 42332 1716 42334
rect 1780 42332 1827 42336
rect 1761 42331 1827 42332
rect 0 42122 800 42152
rect 3785 42122 3851 42125
rect 0 42120 3851 42122
rect 0 42064 3790 42120
rect 3846 42064 3851 42120
rect 0 42062 3851 42064
rect 0 42032 800 42062
rect 3785 42059 3851 42062
rect 4889 42122 4955 42125
rect 5390 42122 5396 42124
rect 4889 42120 5396 42122
rect 4889 42064 4894 42120
rect 4950 42064 5396 42120
rect 4889 42062 5396 42064
rect 4889 42059 4955 42062
rect 5390 42060 5396 42062
rect 5460 42060 5466 42124
rect 3366 41924 3372 41988
rect 3436 41986 3442 41988
rect 3785 41986 3851 41989
rect 3436 41984 3851 41986
rect 3436 41928 3790 41984
rect 3846 41928 3851 41984
rect 3436 41926 3851 41928
rect 3436 41924 3442 41926
rect 3785 41923 3851 41926
rect 4838 41924 4844 41988
rect 4908 41986 4914 41988
rect 5390 41986 5396 41988
rect 4908 41926 5396 41986
rect 4908 41924 4914 41926
rect 5390 41924 5396 41926
rect 5460 41924 5466 41988
rect 2576 41920 2896 41921
rect 2576 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2576 41855 2896 41856
rect 5840 41920 6160 41921
rect 5840 41856 5848 41920
rect 5912 41856 5928 41920
rect 5992 41856 6008 41920
rect 6072 41856 6088 41920
rect 6152 41856 6160 41920
rect 5840 41855 6160 41856
rect 9104 41920 9424 41921
rect 9104 41856 9112 41920
rect 9176 41856 9192 41920
rect 9256 41856 9272 41920
rect 9336 41856 9352 41920
rect 9416 41856 9424 41920
rect 9104 41855 9424 41856
rect 1853 41850 1919 41853
rect 2078 41850 2084 41852
rect 1853 41848 2084 41850
rect 1853 41792 1858 41848
rect 1914 41792 2084 41848
rect 1853 41790 2084 41792
rect 1853 41787 1919 41790
rect 2078 41788 2084 41790
rect 2148 41788 2154 41852
rect 4981 41850 5047 41853
rect 10041 41850 10107 41853
rect 11200 41850 12000 41880
rect 4981 41848 5090 41850
rect 4981 41792 4986 41848
rect 5042 41792 5090 41848
rect 4981 41787 5090 41792
rect 10041 41848 12000 41850
rect 10041 41792 10046 41848
rect 10102 41792 12000 41848
rect 10041 41790 12000 41792
rect 10041 41787 10107 41790
rect 0 41714 800 41744
rect 3417 41714 3483 41717
rect 0 41712 3483 41714
rect 0 41656 3422 41712
rect 3478 41656 3483 41712
rect 0 41654 3483 41656
rect 0 41624 800 41654
rect 3417 41651 3483 41654
rect 1301 41580 1367 41581
rect 1301 41576 1348 41580
rect 1412 41578 1418 41580
rect 3509 41578 3575 41581
rect 5030 41580 5090 41787
rect 11200 41760 12000 41790
rect 3734 41578 3740 41580
rect 1301 41520 1306 41576
rect 1301 41516 1348 41520
rect 1412 41518 1458 41578
rect 3509 41576 3740 41578
rect 3509 41520 3514 41576
rect 3570 41520 3740 41576
rect 3509 41518 3740 41520
rect 1412 41516 1418 41518
rect 1301 41515 1367 41516
rect 3509 41515 3575 41518
rect 3734 41516 3740 41518
rect 3804 41516 3810 41580
rect 5022 41516 5028 41580
rect 5092 41516 5098 41580
rect 54 41380 60 41444
rect 124 41442 130 41444
rect 1025 41442 1091 41445
rect 124 41440 1091 41442
rect 124 41384 1030 41440
rect 1086 41384 1091 41440
rect 124 41382 1091 41384
rect 124 41380 130 41382
rect 1025 41379 1091 41382
rect 1301 41442 1367 41445
rect 1669 41442 1735 41445
rect 1301 41440 1735 41442
rect 1301 41384 1306 41440
rect 1362 41384 1674 41440
rect 1730 41384 1735 41440
rect 1301 41382 1735 41384
rect 1301 41379 1367 41382
rect 1669 41379 1735 41382
rect 3182 41380 3188 41444
rect 3252 41442 3258 41444
rect 3601 41442 3667 41445
rect 3252 41440 3667 41442
rect 3252 41384 3606 41440
rect 3662 41384 3667 41440
rect 3252 41382 3667 41384
rect 3252 41380 3258 41382
rect 3601 41379 3667 41382
rect 3785 41442 3851 41445
rect 3918 41442 3924 41444
rect 3785 41440 3924 41442
rect 3785 41384 3790 41440
rect 3846 41384 3924 41440
rect 3785 41382 3924 41384
rect 3785 41379 3851 41382
rect 3918 41380 3924 41382
rect 3988 41380 3994 41444
rect 4838 41380 4844 41444
rect 4908 41442 4914 41444
rect 5206 41442 5212 41444
rect 4908 41382 5212 41442
rect 4908 41380 4914 41382
rect 5206 41380 5212 41382
rect 5276 41380 5282 41444
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 7472 41376 7792 41377
rect 7472 41312 7480 41376
rect 7544 41312 7560 41376
rect 7624 41312 7640 41376
rect 7704 41312 7720 41376
rect 7784 41312 7792 41376
rect 7472 41311 7792 41312
rect 3601 41308 3667 41309
rect 1342 41244 1348 41308
rect 1412 41306 1418 41308
rect 1710 41306 1716 41308
rect 1412 41246 1716 41306
rect 1412 41244 1418 41246
rect 1710 41244 1716 41246
rect 1780 41244 1786 41308
rect 3550 41306 3556 41308
rect 3510 41246 3556 41306
rect 3620 41304 3667 41308
rect 3877 41306 3943 41309
rect 5257 41308 5323 41309
rect 5206 41306 5212 41308
rect 3662 41248 3667 41304
rect 3550 41244 3556 41246
rect 3620 41244 3667 41248
rect 3601 41243 3667 41244
rect 3742 41304 3943 41306
rect 3742 41248 3882 41304
rect 3938 41248 3943 41304
rect 3742 41246 3943 41248
rect 5166 41246 5212 41306
rect 5276 41304 5323 41308
rect 6729 41306 6795 41309
rect 5318 41248 5323 41304
rect 0 41170 800 41200
rect 2957 41170 3023 41173
rect 0 41168 3023 41170
rect 0 41112 2962 41168
rect 3018 41112 3023 41168
rect 0 41110 3023 41112
rect 0 41080 800 41110
rect 2957 41107 3023 41110
rect 3366 41108 3372 41172
rect 3436 41170 3442 41172
rect 3509 41170 3575 41173
rect 3436 41168 3575 41170
rect 3436 41112 3514 41168
rect 3570 41112 3575 41168
rect 3436 41110 3575 41112
rect 3436 41108 3442 41110
rect 3509 41107 3575 41110
rect 2865 41034 2931 41037
rect 3417 41036 3483 41037
rect 3366 41034 3372 41036
rect 1350 41032 2931 41034
rect 1350 40976 2870 41032
rect 2926 40976 2931 41032
rect 1350 40974 2931 40976
rect 3326 40974 3372 41034
rect 3436 41032 3483 41036
rect 3478 40976 3483 41032
rect 0 40762 800 40792
rect 1350 40762 1410 40974
rect 2865 40971 2931 40974
rect 3366 40972 3372 40974
rect 3436 40972 3483 40976
rect 3550 40972 3556 41036
rect 3620 41034 3626 41036
rect 3742 41034 3802 41246
rect 3877 41243 3943 41246
rect 5206 41244 5212 41246
rect 5276 41244 5323 41248
rect 5257 41243 5323 41244
rect 5398 41304 6795 41306
rect 5398 41248 6734 41304
rect 6790 41248 6795 41304
rect 5398 41246 6795 41248
rect 3620 40974 3802 41034
rect 3620 40972 3626 40974
rect 3417 40971 3483 40972
rect 5257 40898 5323 40901
rect 5398 40898 5458 41246
rect 6729 41243 6795 41246
rect 10041 41034 10107 41037
rect 11200 41034 12000 41064
rect 10041 41032 12000 41034
rect 10041 40976 10046 41032
rect 10102 40976 12000 41032
rect 10041 40974 12000 40976
rect 10041 40971 10107 40974
rect 11200 40944 12000 40974
rect 5257 40896 5458 40898
rect 5257 40840 5262 40896
rect 5318 40840 5458 40896
rect 5257 40838 5458 40840
rect 5257 40835 5323 40838
rect 2576 40832 2896 40833
rect 2576 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2576 40767 2896 40768
rect 5840 40832 6160 40833
rect 5840 40768 5848 40832
rect 5912 40768 5928 40832
rect 5992 40768 6008 40832
rect 6072 40768 6088 40832
rect 6152 40768 6160 40832
rect 5840 40767 6160 40768
rect 9104 40832 9424 40833
rect 9104 40768 9112 40832
rect 9176 40768 9192 40832
rect 9256 40768 9272 40832
rect 9336 40768 9352 40832
rect 9416 40768 9424 40832
rect 9104 40767 9424 40768
rect 0 40702 1410 40762
rect 0 40672 800 40702
rect 4981 40626 5047 40629
rect 4662 40624 5047 40626
rect 4662 40568 4986 40624
rect 5042 40568 5047 40624
rect 4662 40566 5047 40568
rect 2400 40428 2406 40492
rect 2470 40490 2476 40492
rect 2589 40490 2655 40493
rect 3417 40490 3483 40493
rect 2470 40488 2655 40490
rect 2470 40432 2594 40488
rect 2650 40432 2655 40488
rect 2470 40430 2655 40432
rect 2470 40428 2476 40430
rect 2589 40427 2655 40430
rect 2730 40488 3483 40490
rect 2730 40432 3422 40488
rect 3478 40432 3483 40488
rect 2730 40430 3483 40432
rect 0 40354 800 40384
rect 2730 40354 2790 40430
rect 3417 40427 3483 40430
rect 0 40294 2790 40354
rect 0 40264 800 40294
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 4521 40082 4587 40085
rect 4662 40082 4722 40566
rect 4981 40563 5047 40566
rect 10041 40354 10107 40357
rect 11200 40354 12000 40384
rect 10041 40352 12000 40354
rect 10041 40296 10046 40352
rect 10102 40296 12000 40352
rect 10041 40294 12000 40296
rect 10041 40291 10107 40294
rect 7472 40288 7792 40289
rect 7472 40224 7480 40288
rect 7544 40224 7560 40288
rect 7624 40224 7640 40288
rect 7704 40224 7720 40288
rect 7784 40224 7792 40288
rect 11200 40264 12000 40294
rect 7472 40223 7792 40224
rect 4521 40080 4722 40082
rect 4521 40024 4526 40080
rect 4582 40024 4722 40080
rect 4521 40022 4722 40024
rect 4521 40019 4587 40022
rect 0 39946 800 39976
rect 3325 39946 3391 39949
rect 0 39944 3391 39946
rect 0 39888 3330 39944
rect 3386 39888 3391 39944
rect 0 39886 3391 39888
rect 0 39856 800 39886
rect 3325 39883 3391 39886
rect 4705 39946 4771 39949
rect 5390 39946 5396 39948
rect 4705 39944 5396 39946
rect 4705 39888 4710 39944
rect 4766 39888 5396 39944
rect 4705 39886 5396 39888
rect 4705 39883 4771 39886
rect 5390 39884 5396 39886
rect 5460 39884 5466 39948
rect 3969 39810 4035 39813
rect 3374 39808 4035 39810
rect 3374 39752 3974 39808
rect 4030 39752 4035 39808
rect 3374 39750 4035 39752
rect 2576 39744 2896 39745
rect 2576 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2576 39679 2896 39680
rect 0 39538 800 39568
rect 3374 39538 3434 39750
rect 3969 39747 4035 39750
rect 5840 39744 6160 39745
rect 5840 39680 5848 39744
rect 5912 39680 5928 39744
rect 5992 39680 6008 39744
rect 6072 39680 6088 39744
rect 6152 39680 6160 39744
rect 5840 39679 6160 39680
rect 9104 39744 9424 39745
rect 9104 39680 9112 39744
rect 9176 39680 9192 39744
rect 9256 39680 9272 39744
rect 9336 39680 9352 39744
rect 9416 39680 9424 39744
rect 9104 39679 9424 39680
rect 0 39478 3434 39538
rect 0 39448 800 39478
rect 3918 39476 3924 39540
rect 3988 39538 3994 39540
rect 6494 39538 6500 39540
rect 3988 39478 6500 39538
rect 3988 39476 3994 39478
rect 6494 39476 6500 39478
rect 6564 39476 6570 39540
rect 10041 39538 10107 39541
rect 11200 39538 12000 39568
rect 10041 39536 12000 39538
rect 10041 39480 10046 39536
rect 10102 39480 12000 39536
rect 10041 39478 12000 39480
rect 10041 39475 10107 39478
rect 11200 39448 12000 39478
rect 1393 39402 1459 39405
rect 1710 39402 1716 39404
rect 1393 39400 1716 39402
rect 1393 39344 1398 39400
rect 1454 39344 1716 39400
rect 1393 39342 1716 39344
rect 1393 39339 1459 39342
rect 1710 39340 1716 39342
rect 1780 39340 1786 39404
rect 3877 39402 3943 39405
rect 4245 39402 4311 39405
rect 3877 39400 4311 39402
rect 3877 39344 3882 39400
rect 3938 39344 4250 39400
rect 4306 39344 4311 39400
rect 3877 39342 4311 39344
rect 3877 39339 3943 39342
rect 4245 39339 4311 39342
rect 1117 39266 1183 39269
rect 3182 39266 3188 39268
rect 1117 39264 3188 39266
rect 1117 39208 1122 39264
rect 1178 39208 3188 39264
rect 1117 39206 3188 39208
rect 1117 39203 1183 39206
rect 3182 39204 3188 39206
rect 3252 39204 3258 39268
rect 4208 39200 4528 39201
rect 0 39130 800 39160
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 7472 39200 7792 39201
rect 7472 39136 7480 39200
rect 7544 39136 7560 39200
rect 7624 39136 7640 39200
rect 7704 39136 7720 39200
rect 7784 39136 7792 39200
rect 7472 39135 7792 39136
rect 3785 39130 3851 39133
rect 0 39128 3851 39130
rect 0 39072 3790 39128
rect 3846 39072 3851 39128
rect 0 39070 3851 39072
rect 0 39040 800 39070
rect 3785 39067 3851 39070
rect 2078 38932 2084 38996
rect 2148 38994 2154 38996
rect 2221 38994 2287 38997
rect 2148 38992 2287 38994
rect 2148 38936 2226 38992
rect 2282 38936 2287 38992
rect 2148 38934 2287 38936
rect 2148 38932 2154 38934
rect 2221 38931 2287 38934
rect 4337 38994 4403 38997
rect 6310 38994 6316 38996
rect 4337 38992 6316 38994
rect 4337 38936 4342 38992
rect 4398 38936 6316 38992
rect 4337 38934 6316 38936
rect 4337 38931 4403 38934
rect 6310 38932 6316 38934
rect 6380 38932 6386 38996
rect 422 38796 428 38860
rect 492 38858 498 38860
rect 1301 38858 1367 38861
rect 492 38856 1367 38858
rect 492 38800 1306 38856
rect 1362 38800 1367 38856
rect 492 38798 1367 38800
rect 492 38796 498 38798
rect 1301 38795 1367 38798
rect 2078 38796 2084 38860
rect 2148 38858 2154 38860
rect 2589 38858 2655 38861
rect 2148 38856 2655 38858
rect 2148 38800 2594 38856
rect 2650 38800 2655 38856
rect 2148 38798 2655 38800
rect 2148 38796 2154 38798
rect 2589 38795 2655 38798
rect 2773 38858 2839 38861
rect 3550 38858 3556 38860
rect 2773 38856 3556 38858
rect 2773 38800 2778 38856
rect 2834 38800 3556 38856
rect 2773 38798 3556 38800
rect 2773 38795 2839 38798
rect 3550 38796 3556 38798
rect 3620 38796 3626 38860
rect 1117 38722 1183 38725
rect 1117 38720 2514 38722
rect 1117 38664 1122 38720
rect 1178 38664 2514 38720
rect 1117 38662 2514 38664
rect 1117 38659 1183 38662
rect 0 38586 800 38616
rect 933 38586 999 38589
rect 0 38584 999 38586
rect 0 38528 938 38584
rect 994 38528 999 38584
rect 0 38526 999 38528
rect 0 38496 800 38526
rect 933 38523 999 38526
rect 1301 38584 1367 38589
rect 1301 38528 1306 38584
rect 1362 38528 1367 38584
rect 1301 38523 1367 38528
rect 1577 38584 1643 38589
rect 1577 38528 1582 38584
rect 1638 38528 1643 38584
rect 1577 38523 1643 38528
rect 1304 38317 1364 38523
rect 1580 38453 1640 38523
rect 1577 38448 1643 38453
rect 1577 38392 1582 38448
rect 1638 38392 1643 38448
rect 1577 38387 1643 38392
rect 2454 38450 2514 38662
rect 3141 38720 3207 38725
rect 3141 38664 3146 38720
rect 3202 38664 3207 38720
rect 3141 38659 3207 38664
rect 10041 38722 10107 38725
rect 11200 38722 12000 38752
rect 10041 38720 12000 38722
rect 10041 38664 10046 38720
rect 10102 38664 12000 38720
rect 10041 38662 12000 38664
rect 10041 38659 10107 38662
rect 2576 38656 2896 38657
rect 2576 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2576 38591 2896 38592
rect 3144 38589 3204 38659
rect 5840 38656 6160 38657
rect 5840 38592 5848 38656
rect 5912 38592 5928 38656
rect 5992 38592 6008 38656
rect 6072 38592 6088 38656
rect 6152 38592 6160 38656
rect 5840 38591 6160 38592
rect 9104 38656 9424 38657
rect 9104 38592 9112 38656
rect 9176 38592 9192 38656
rect 9256 38592 9272 38656
rect 9336 38592 9352 38656
rect 9416 38592 9424 38656
rect 11200 38632 12000 38662
rect 9104 38591 9424 38592
rect 3141 38584 3207 38589
rect 3141 38528 3146 38584
rect 3202 38528 3207 38584
rect 3141 38523 3207 38528
rect 2773 38450 2839 38453
rect 3877 38450 3943 38453
rect 2454 38448 2839 38450
rect 2454 38392 2778 38448
rect 2834 38392 2839 38448
rect 2454 38390 2839 38392
rect 2773 38387 2839 38390
rect 3006 38448 3943 38450
rect 3006 38392 3882 38448
rect 3938 38392 3943 38448
rect 3006 38390 3943 38392
rect 1301 38312 1367 38317
rect 1301 38256 1306 38312
rect 1362 38256 1367 38312
rect 1301 38251 1367 38256
rect 1485 38314 1551 38317
rect 3006 38314 3066 38390
rect 3877 38387 3943 38390
rect 1485 38312 3066 38314
rect 1485 38256 1490 38312
rect 1546 38256 3066 38312
rect 1485 38254 3066 38256
rect 1485 38251 1551 38254
rect 3182 38252 3188 38316
rect 3252 38314 3258 38316
rect 3325 38314 3391 38317
rect 3252 38312 3391 38314
rect 3252 38256 3330 38312
rect 3386 38256 3391 38312
rect 3252 38254 3391 38256
rect 3252 38252 3258 38254
rect 3325 38251 3391 38254
rect 4337 38314 4403 38317
rect 4337 38312 4722 38314
rect 4337 38256 4342 38312
rect 4398 38256 4722 38312
rect 4337 38254 4722 38256
rect 4337 38251 4403 38254
rect 0 38178 800 38208
rect 0 38118 1778 38178
rect 0 38088 800 38118
rect 1718 37906 1778 38118
rect 2078 38116 2084 38180
rect 2148 38178 2154 38180
rect 2313 38178 2379 38181
rect 2148 38176 2379 38178
rect 2148 38120 2318 38176
rect 2374 38120 2379 38176
rect 2148 38118 2379 38120
rect 2148 38116 2154 38118
rect 2313 38115 2379 38118
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 1853 37906 1919 37909
rect 1718 37904 1919 37906
rect 1718 37848 1858 37904
rect 1914 37848 1919 37904
rect 1718 37846 1919 37848
rect 1853 37843 1919 37846
rect 3141 37906 3207 37909
rect 3366 37906 3372 37908
rect 3141 37904 3372 37906
rect 3141 37848 3146 37904
rect 3202 37848 3372 37904
rect 3141 37846 3372 37848
rect 3141 37843 3207 37846
rect 3366 37844 3372 37846
rect 3436 37844 3442 37908
rect 0 37770 800 37800
rect 3509 37770 3575 37773
rect 0 37768 3575 37770
rect 0 37712 3514 37768
rect 3570 37712 3575 37768
rect 0 37710 3575 37712
rect 0 37680 800 37710
rect 3509 37707 3575 37710
rect 3785 37770 3851 37773
rect 4662 37770 4722 38254
rect 7472 38112 7792 38113
rect 7472 38048 7480 38112
rect 7544 38048 7560 38112
rect 7624 38048 7640 38112
rect 7704 38048 7720 38112
rect 7784 38048 7792 38112
rect 7472 38047 7792 38048
rect 10041 38042 10107 38045
rect 11200 38042 12000 38072
rect 10041 38040 12000 38042
rect 10041 37984 10046 38040
rect 10102 37984 12000 38040
rect 10041 37982 12000 37984
rect 10041 37979 10107 37982
rect 11200 37952 12000 37982
rect 3785 37768 4722 37770
rect 3785 37712 3790 37768
rect 3846 37712 4722 37768
rect 3785 37710 4722 37712
rect 3785 37707 3851 37710
rect 2576 37568 2896 37569
rect 2576 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2576 37503 2896 37504
rect 5840 37568 6160 37569
rect 5840 37504 5848 37568
rect 5912 37504 5928 37568
rect 5992 37504 6008 37568
rect 6072 37504 6088 37568
rect 6152 37504 6160 37568
rect 5840 37503 6160 37504
rect 9104 37568 9424 37569
rect 9104 37504 9112 37568
rect 9176 37504 9192 37568
rect 9256 37504 9272 37568
rect 9336 37504 9352 37568
rect 9416 37504 9424 37568
rect 9104 37503 9424 37504
rect 0 37362 800 37392
rect 3417 37362 3483 37365
rect 0 37360 3483 37362
rect 0 37304 3422 37360
rect 3478 37304 3483 37360
rect 0 37302 3483 37304
rect 0 37272 800 37302
rect 3417 37299 3483 37302
rect 10041 37226 10107 37229
rect 11200 37226 12000 37256
rect 10041 37224 12000 37226
rect 10041 37168 10046 37224
rect 10102 37168 12000 37224
rect 10041 37166 12000 37168
rect 10041 37163 10107 37166
rect 11200 37136 12000 37166
rect 4208 37024 4528 37025
rect 0 36954 800 36984
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 7472 37024 7792 37025
rect 7472 36960 7480 37024
rect 7544 36960 7560 37024
rect 7624 36960 7640 37024
rect 7704 36960 7720 37024
rect 7784 36960 7792 37024
rect 7472 36959 7792 36960
rect 933 36954 999 36957
rect 0 36952 999 36954
rect 0 36896 938 36952
rect 994 36896 999 36952
rect 0 36894 999 36896
rect 0 36864 800 36894
rect 933 36891 999 36894
rect 2262 36756 2268 36820
rect 2332 36818 2338 36820
rect 4521 36818 4587 36821
rect 5022 36818 5028 36820
rect 2332 36758 3618 36818
rect 2332 36756 2338 36758
rect 3417 36682 3483 36685
rect 1350 36680 3483 36682
rect 1350 36624 3422 36680
rect 3478 36624 3483 36680
rect 1350 36622 3483 36624
rect 0 36546 800 36576
rect 1350 36546 1410 36622
rect 3417 36619 3483 36622
rect 2313 36548 2379 36549
rect 0 36486 1410 36546
rect 0 36456 800 36486
rect 2262 36484 2268 36548
rect 2332 36546 2379 36548
rect 3417 36546 3483 36549
rect 3558 36546 3618 36758
rect 4521 36816 5028 36818
rect 4521 36760 4526 36816
rect 4582 36760 5028 36816
rect 4521 36758 5028 36760
rect 4521 36755 4587 36758
rect 5022 36756 5028 36758
rect 5092 36756 5098 36820
rect 2332 36544 2424 36546
rect 2374 36488 2424 36544
rect 2332 36486 2424 36488
rect 3417 36544 3618 36546
rect 3417 36488 3422 36544
rect 3478 36488 3618 36544
rect 3417 36486 3618 36488
rect 2332 36484 2379 36486
rect 2313 36483 2379 36484
rect 3417 36483 3483 36486
rect 2576 36480 2896 36481
rect 2576 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2576 36415 2896 36416
rect 5840 36480 6160 36481
rect 5840 36416 5848 36480
rect 5912 36416 5928 36480
rect 5992 36416 6008 36480
rect 6072 36416 6088 36480
rect 6152 36416 6160 36480
rect 5840 36415 6160 36416
rect 9104 36480 9424 36481
rect 9104 36416 9112 36480
rect 9176 36416 9192 36480
rect 9256 36416 9272 36480
rect 9336 36416 9352 36480
rect 9416 36416 9424 36480
rect 9104 36415 9424 36416
rect 10041 36410 10107 36413
rect 11200 36410 12000 36440
rect 10041 36408 12000 36410
rect 10041 36352 10046 36408
rect 10102 36352 12000 36408
rect 10041 36350 12000 36352
rect 10041 36347 10107 36350
rect 11200 36320 12000 36350
rect 0 36138 800 36168
rect 1577 36138 1643 36141
rect 0 36136 1643 36138
rect 0 36080 1582 36136
rect 1638 36080 1643 36136
rect 0 36078 1643 36080
rect 0 36048 800 36078
rect 1577 36075 1643 36078
rect 1894 36076 1900 36140
rect 1964 36138 1970 36140
rect 2957 36138 3023 36141
rect 1964 36136 3023 36138
rect 1964 36080 2962 36136
rect 3018 36080 3023 36136
rect 1964 36078 3023 36080
rect 1964 36076 1970 36078
rect 2957 36075 3023 36078
rect 4797 36002 4863 36005
rect 5022 36002 5028 36004
rect 4797 36000 5028 36002
rect 4797 35944 4802 36000
rect 4858 35944 5028 36000
rect 4797 35942 5028 35944
rect 4797 35939 4863 35942
rect 5022 35940 5028 35942
rect 5092 35940 5098 36004
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 7472 35936 7792 35937
rect 7472 35872 7480 35936
rect 7544 35872 7560 35936
rect 7624 35872 7640 35936
rect 7704 35872 7720 35936
rect 7784 35872 7792 35936
rect 7472 35871 7792 35872
rect 4613 35730 4679 35733
rect 5390 35730 5396 35732
rect 4613 35728 5396 35730
rect 4613 35672 4618 35728
rect 4674 35672 5396 35728
rect 4613 35670 5396 35672
rect 4613 35667 4679 35670
rect 5390 35668 5396 35670
rect 5460 35668 5466 35732
rect 10041 35730 10107 35733
rect 11200 35730 12000 35760
rect 10041 35728 12000 35730
rect 10041 35672 10046 35728
rect 10102 35672 12000 35728
rect 10041 35670 12000 35672
rect 10041 35667 10107 35670
rect 11200 35640 12000 35670
rect 0 35594 800 35624
rect 2313 35594 2379 35597
rect 0 35592 2379 35594
rect 0 35536 2318 35592
rect 2374 35536 2379 35592
rect 0 35534 2379 35536
rect 0 35504 800 35534
rect 2313 35531 2379 35534
rect 2576 35392 2896 35393
rect 2576 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2576 35327 2896 35328
rect 5840 35392 6160 35393
rect 5840 35328 5848 35392
rect 5912 35328 5928 35392
rect 5992 35328 6008 35392
rect 6072 35328 6088 35392
rect 6152 35328 6160 35392
rect 5840 35327 6160 35328
rect 9104 35392 9424 35393
rect 9104 35328 9112 35392
rect 9176 35328 9192 35392
rect 9256 35328 9272 35392
rect 9336 35328 9352 35392
rect 9416 35328 9424 35392
rect 9104 35327 9424 35328
rect 3785 35324 3851 35325
rect 3734 35260 3740 35324
rect 3804 35322 3851 35324
rect 3804 35320 3896 35322
rect 3846 35264 3896 35320
rect 3804 35262 3896 35264
rect 3804 35260 3851 35262
rect 3785 35259 3851 35260
rect 0 35186 800 35216
rect 1577 35186 1643 35189
rect 3693 35188 3759 35189
rect 3693 35186 3740 35188
rect 0 35184 1643 35186
rect 0 35128 1582 35184
rect 1638 35128 1643 35184
rect 0 35126 1643 35128
rect 3648 35184 3740 35186
rect 3648 35128 3698 35184
rect 3648 35126 3740 35128
rect 0 35096 800 35126
rect 1577 35123 1643 35126
rect 3693 35124 3740 35126
rect 3804 35124 3810 35188
rect 3693 35123 3759 35124
rect 10041 34914 10107 34917
rect 11200 34914 12000 34944
rect 10041 34912 12000 34914
rect 10041 34856 10046 34912
rect 10102 34856 12000 34912
rect 10041 34854 12000 34856
rect 10041 34851 10107 34854
rect 4208 34848 4528 34849
rect 0 34778 800 34808
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 7472 34848 7792 34849
rect 7472 34784 7480 34848
rect 7544 34784 7560 34848
rect 7624 34784 7640 34848
rect 7704 34784 7720 34848
rect 7784 34784 7792 34848
rect 11200 34824 12000 34854
rect 7472 34783 7792 34784
rect 1577 34778 1643 34781
rect 0 34776 1643 34778
rect 0 34720 1582 34776
rect 1638 34720 1643 34776
rect 0 34718 1643 34720
rect 0 34688 800 34718
rect 1577 34715 1643 34718
rect 2773 34506 2839 34509
rect 1350 34504 2839 34506
rect 1350 34448 2778 34504
rect 2834 34448 2839 34504
rect 1350 34446 2839 34448
rect 0 34370 800 34400
rect 1350 34370 1410 34446
rect 2773 34443 2839 34446
rect 0 34310 1410 34370
rect 0 34280 800 34310
rect 2576 34304 2896 34305
rect 2576 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2576 34239 2896 34240
rect 5840 34304 6160 34305
rect 5840 34240 5848 34304
rect 5912 34240 5928 34304
rect 5992 34240 6008 34304
rect 6072 34240 6088 34304
rect 6152 34240 6160 34304
rect 5840 34239 6160 34240
rect 9104 34304 9424 34305
rect 9104 34240 9112 34304
rect 9176 34240 9192 34304
rect 9256 34240 9272 34304
rect 9336 34240 9352 34304
rect 9416 34240 9424 34304
rect 9104 34239 9424 34240
rect 9581 34098 9647 34101
rect 11200 34098 12000 34128
rect 9581 34096 12000 34098
rect 9581 34040 9586 34096
rect 9642 34040 12000 34096
rect 9581 34038 12000 34040
rect 9581 34035 9647 34038
rect 11200 34008 12000 34038
rect 0 33962 800 33992
rect 3049 33962 3115 33965
rect 4153 33962 4219 33965
rect 0 33960 3115 33962
rect 0 33904 3054 33960
rect 3110 33904 3115 33960
rect 0 33902 3115 33904
rect 0 33872 800 33902
rect 3049 33899 3115 33902
rect 3788 33960 4219 33962
rect 3788 33904 4158 33960
rect 4214 33904 4219 33960
rect 3788 33902 4219 33904
rect 3788 33829 3848 33902
rect 4153 33899 4219 33902
rect 3785 33824 3851 33829
rect 3785 33768 3790 33824
rect 3846 33768 3851 33824
rect 3785 33763 3851 33768
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 7472 33760 7792 33761
rect 7472 33696 7480 33760
rect 7544 33696 7560 33760
rect 7624 33696 7640 33760
rect 7704 33696 7720 33760
rect 7784 33696 7792 33760
rect 7472 33695 7792 33696
rect 0 33554 800 33584
rect 1393 33554 1459 33557
rect 0 33552 1459 33554
rect 0 33496 1398 33552
rect 1454 33496 1459 33552
rect 0 33494 1459 33496
rect 0 33464 800 33494
rect 1393 33491 1459 33494
rect 10041 33418 10107 33421
rect 11200 33418 12000 33448
rect 10041 33416 12000 33418
rect 10041 33360 10046 33416
rect 10102 33360 12000 33416
rect 10041 33358 12000 33360
rect 10041 33355 10107 33358
rect 11200 33328 12000 33358
rect 1342 33220 1348 33284
rect 1412 33282 1418 33284
rect 1485 33282 1551 33285
rect 1412 33280 1551 33282
rect 1412 33224 1490 33280
rect 1546 33224 1551 33280
rect 1412 33222 1551 33224
rect 1412 33220 1418 33222
rect 1485 33219 1551 33222
rect 2576 33216 2896 33217
rect 0 33146 800 33176
rect 2576 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2576 33151 2896 33152
rect 5840 33216 6160 33217
rect 5840 33152 5848 33216
rect 5912 33152 5928 33216
rect 5992 33152 6008 33216
rect 6072 33152 6088 33216
rect 6152 33152 6160 33216
rect 5840 33151 6160 33152
rect 9104 33216 9424 33217
rect 9104 33152 9112 33216
rect 9176 33152 9192 33216
rect 9256 33152 9272 33216
rect 9336 33152 9352 33216
rect 9416 33152 9424 33216
rect 9104 33151 9424 33152
rect 0 33086 1410 33146
rect 0 33056 800 33086
rect 1350 33010 1410 33086
rect 1350 32950 2790 33010
rect 2730 32877 2790 32950
rect 749 32876 815 32877
rect 749 32874 796 32876
rect 704 32872 796 32874
rect 704 32816 754 32872
rect 704 32814 796 32816
rect 749 32812 796 32814
rect 860 32812 866 32876
rect 1158 32812 1164 32876
rect 1228 32874 1234 32876
rect 1485 32874 1551 32877
rect 1228 32872 1551 32874
rect 1228 32816 1490 32872
rect 1546 32816 1551 32872
rect 1228 32814 1551 32816
rect 2730 32872 2839 32877
rect 2730 32816 2778 32872
rect 2834 32816 2839 32872
rect 2730 32814 2839 32816
rect 1228 32812 1234 32814
rect 749 32811 815 32812
rect 1485 32811 1551 32814
rect 2773 32811 2839 32814
rect 1526 32676 1532 32740
rect 1596 32738 1602 32740
rect 2129 32738 2195 32741
rect 1596 32736 2195 32738
rect 1596 32680 2134 32736
rect 2190 32680 2195 32736
rect 1596 32678 2195 32680
rect 1596 32676 1602 32678
rect 2129 32675 2195 32678
rect 4208 32672 4528 32673
rect 0 32602 800 32632
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 7472 32672 7792 32673
rect 7472 32608 7480 32672
rect 7544 32608 7560 32672
rect 7624 32608 7640 32672
rect 7704 32608 7720 32672
rect 7784 32608 7792 32672
rect 7472 32607 7792 32608
rect 2313 32602 2379 32605
rect 0 32600 2379 32602
rect 0 32544 2318 32600
rect 2374 32544 2379 32600
rect 0 32542 2379 32544
rect 0 32512 800 32542
rect 2313 32539 2379 32542
rect 10041 32602 10107 32605
rect 11200 32602 12000 32632
rect 10041 32600 12000 32602
rect 10041 32544 10046 32600
rect 10102 32544 12000 32600
rect 10041 32542 12000 32544
rect 10041 32539 10107 32542
rect 11200 32512 12000 32542
rect 3918 32404 3924 32468
rect 3988 32466 3994 32468
rect 4245 32466 4311 32469
rect 3988 32464 4311 32466
rect 3988 32408 4250 32464
rect 4306 32408 4311 32464
rect 3988 32406 4311 32408
rect 3988 32404 3994 32406
rect 4245 32403 4311 32406
rect 3049 32330 3115 32333
rect 1350 32328 3115 32330
rect 1350 32272 3054 32328
rect 3110 32272 3115 32328
rect 1350 32270 3115 32272
rect 0 32194 800 32224
rect 1350 32194 1410 32270
rect 3049 32267 3115 32270
rect 0 32134 1410 32194
rect 1669 32196 1735 32197
rect 1669 32192 1716 32196
rect 1780 32194 1786 32196
rect 5165 32194 5231 32197
rect 5625 32194 5691 32197
rect 1669 32136 1674 32192
rect 0 32104 800 32134
rect 1669 32132 1716 32136
rect 1780 32134 1826 32194
rect 5165 32192 5691 32194
rect 5165 32136 5170 32192
rect 5226 32136 5630 32192
rect 5686 32136 5691 32192
rect 5165 32134 5691 32136
rect 1780 32132 1786 32134
rect 1669 32131 1735 32132
rect 5165 32131 5231 32134
rect 5625 32131 5691 32134
rect 2576 32128 2896 32129
rect 2576 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2576 32063 2896 32064
rect 5840 32128 6160 32129
rect 5840 32064 5848 32128
rect 5912 32064 5928 32128
rect 5992 32064 6008 32128
rect 6072 32064 6088 32128
rect 6152 32064 6160 32128
rect 5840 32063 6160 32064
rect 9104 32128 9424 32129
rect 9104 32064 9112 32128
rect 9176 32064 9192 32128
rect 9256 32064 9272 32128
rect 9336 32064 9352 32128
rect 9416 32064 9424 32128
rect 9104 32063 9424 32064
rect 3417 32058 3483 32061
rect 3969 32060 4035 32061
rect 3550 32058 3556 32060
rect 3417 32056 3556 32058
rect 3417 32000 3422 32056
rect 3478 32000 3556 32056
rect 3417 31998 3556 32000
rect 3417 31995 3483 31998
rect 3550 31996 3556 31998
rect 3620 31996 3626 32060
rect 3918 31996 3924 32060
rect 3988 32058 4035 32060
rect 3988 32056 4080 32058
rect 4030 32000 4080 32056
rect 3988 31998 4080 32000
rect 3988 31996 4035 31998
rect 3969 31995 4035 31996
rect 1393 31922 1459 31925
rect 1526 31922 1532 31924
rect 1393 31920 1532 31922
rect 1393 31864 1398 31920
rect 1454 31864 1532 31920
rect 1393 31862 1532 31864
rect 1393 31859 1459 31862
rect 1526 31860 1532 31862
rect 1596 31860 1602 31924
rect 0 31786 800 31816
rect 3969 31786 4035 31789
rect 0 31784 4035 31786
rect 0 31728 3974 31784
rect 4030 31728 4035 31784
rect 0 31726 4035 31728
rect 0 31696 800 31726
rect 3969 31723 4035 31726
rect 4521 31786 4587 31789
rect 10041 31786 10107 31789
rect 11200 31786 12000 31816
rect 4521 31784 4722 31786
rect 4521 31728 4526 31784
rect 4582 31728 4722 31784
rect 4521 31726 4722 31728
rect 4521 31723 4587 31726
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 1485 31516 1551 31517
rect 1485 31514 1532 31516
rect 1440 31512 1532 31514
rect 1440 31456 1490 31512
rect 1440 31454 1532 31456
rect 1485 31452 1532 31454
rect 1596 31452 1602 31516
rect 1485 31451 1551 31452
rect 0 31378 800 31408
rect 1117 31378 1183 31381
rect 0 31376 1183 31378
rect 0 31320 1122 31376
rect 1178 31320 1183 31376
rect 0 31318 1183 31320
rect 0 31288 800 31318
rect 1117 31315 1183 31318
rect 4521 31378 4587 31381
rect 4662 31378 4722 31726
rect 10041 31784 12000 31786
rect 10041 31728 10046 31784
rect 10102 31728 12000 31784
rect 10041 31726 12000 31728
rect 10041 31723 10107 31726
rect 11200 31696 12000 31726
rect 5533 31650 5599 31653
rect 4521 31376 4722 31378
rect 4521 31320 4526 31376
rect 4582 31320 4722 31376
rect 4521 31318 4722 31320
rect 5398 31648 5599 31650
rect 5398 31592 5538 31648
rect 5594 31592 5599 31648
rect 5398 31590 5599 31592
rect 4521 31315 4587 31318
rect 4981 31242 5047 31245
rect 5398 31242 5458 31590
rect 5533 31587 5599 31590
rect 7472 31584 7792 31585
rect 7472 31520 7480 31584
rect 7544 31520 7560 31584
rect 7624 31520 7640 31584
rect 7704 31520 7720 31584
rect 7784 31520 7792 31584
rect 7472 31519 7792 31520
rect 4981 31240 5458 31242
rect 4981 31184 4986 31240
rect 5042 31184 5458 31240
rect 4981 31182 5458 31184
rect 4981 31179 5047 31182
rect 5390 31044 5396 31108
rect 5460 31106 5466 31108
rect 5533 31106 5599 31109
rect 5460 31104 5599 31106
rect 5460 31048 5538 31104
rect 5594 31048 5599 31104
rect 5460 31046 5599 31048
rect 5460 31044 5466 31046
rect 5533 31043 5599 31046
rect 10041 31106 10107 31109
rect 11200 31106 12000 31136
rect 10041 31104 12000 31106
rect 10041 31048 10046 31104
rect 10102 31048 12000 31104
rect 10041 31046 12000 31048
rect 10041 31043 10107 31046
rect 2576 31040 2896 31041
rect 0 30970 800 31000
rect 2576 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2576 30975 2896 30976
rect 5840 31040 6160 31041
rect 5840 30976 5848 31040
rect 5912 30976 5928 31040
rect 5992 30976 6008 31040
rect 6072 30976 6088 31040
rect 6152 30976 6160 31040
rect 5840 30975 6160 30976
rect 9104 31040 9424 31041
rect 9104 30976 9112 31040
rect 9176 30976 9192 31040
rect 9256 30976 9272 31040
rect 9336 30976 9352 31040
rect 9416 30976 9424 31040
rect 11200 31016 12000 31046
rect 9104 30975 9424 30976
rect 0 30910 1456 30970
rect 0 30880 800 30910
rect 1396 30834 1456 30910
rect 3325 30834 3391 30837
rect 1396 30832 3391 30834
rect 1396 30776 3330 30832
rect 3386 30776 3391 30832
rect 1396 30774 3391 30776
rect 3325 30771 3391 30774
rect 0 30562 800 30592
rect 2773 30562 2839 30565
rect 0 30560 2839 30562
rect 0 30504 2778 30560
rect 2834 30504 2839 30560
rect 0 30502 2839 30504
rect 0 30472 800 30502
rect 2773 30499 2839 30502
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 7472 30496 7792 30497
rect 7472 30432 7480 30496
rect 7544 30432 7560 30496
rect 7624 30432 7640 30496
rect 7704 30432 7720 30496
rect 7784 30432 7792 30496
rect 7472 30431 7792 30432
rect 974 30228 980 30292
rect 1044 30290 1050 30292
rect 1117 30290 1183 30293
rect 2313 30290 2379 30293
rect 1044 30288 1183 30290
rect 1044 30232 1122 30288
rect 1178 30232 1183 30288
rect 1044 30230 1183 30232
rect 1044 30228 1050 30230
rect 1117 30227 1183 30230
rect 2270 30288 2379 30290
rect 2270 30232 2318 30288
rect 2374 30232 2379 30288
rect 2270 30227 2379 30232
rect 10041 30290 10107 30293
rect 11200 30290 12000 30320
rect 10041 30288 12000 30290
rect 10041 30232 10046 30288
rect 10102 30232 12000 30288
rect 10041 30230 12000 30232
rect 10041 30227 10107 30230
rect 0 30154 800 30184
rect 1853 30154 1919 30157
rect 0 30152 1919 30154
rect 0 30096 1858 30152
rect 1914 30096 1919 30152
rect 0 30094 1919 30096
rect 0 30064 800 30094
rect 1853 30091 1919 30094
rect 2037 30154 2103 30157
rect 2270 30154 2330 30227
rect 11200 30200 12000 30230
rect 2037 30152 2330 30154
rect 2037 30096 2042 30152
rect 2098 30096 2330 30152
rect 2037 30094 2330 30096
rect 2037 30091 2103 30094
rect 2576 29952 2896 29953
rect 2576 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2576 29887 2896 29888
rect 5840 29952 6160 29953
rect 5840 29888 5848 29952
rect 5912 29888 5928 29952
rect 5992 29888 6008 29952
rect 6072 29888 6088 29952
rect 6152 29888 6160 29952
rect 5840 29887 6160 29888
rect 9104 29952 9424 29953
rect 9104 29888 9112 29952
rect 9176 29888 9192 29952
rect 9256 29888 9272 29952
rect 9336 29888 9352 29952
rect 9416 29888 9424 29952
rect 9104 29887 9424 29888
rect 0 29610 800 29640
rect 2773 29610 2839 29613
rect 0 29608 2839 29610
rect 0 29552 2778 29608
rect 2834 29552 2839 29608
rect 0 29550 2839 29552
rect 0 29520 800 29550
rect 2773 29547 2839 29550
rect 10133 29474 10199 29477
rect 11200 29474 12000 29504
rect 10133 29472 12000 29474
rect 10133 29416 10138 29472
rect 10194 29416 12000 29472
rect 10133 29414 12000 29416
rect 10133 29411 10199 29414
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 7472 29408 7792 29409
rect 7472 29344 7480 29408
rect 7544 29344 7560 29408
rect 7624 29344 7640 29408
rect 7704 29344 7720 29408
rect 7784 29344 7792 29408
rect 11200 29384 12000 29414
rect 7472 29343 7792 29344
rect 2957 29338 3023 29341
rect 3366 29338 3372 29340
rect 2957 29336 3372 29338
rect 2957 29280 2962 29336
rect 3018 29280 3372 29336
rect 2957 29278 3372 29280
rect 2957 29275 3023 29278
rect 3366 29276 3372 29278
rect 3436 29276 3442 29340
rect 0 29202 800 29232
rect 1669 29202 1735 29205
rect 0 29200 1735 29202
rect 0 29144 1674 29200
rect 1730 29144 1735 29200
rect 0 29142 1735 29144
rect 0 29112 800 29142
rect 1669 29139 1735 29142
rect 2576 28864 2896 28865
rect 0 28794 800 28824
rect 2576 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2576 28799 2896 28800
rect 5840 28864 6160 28865
rect 5840 28800 5848 28864
rect 5912 28800 5928 28864
rect 5992 28800 6008 28864
rect 6072 28800 6088 28864
rect 6152 28800 6160 28864
rect 5840 28799 6160 28800
rect 9104 28864 9424 28865
rect 9104 28800 9112 28864
rect 9176 28800 9192 28864
rect 9256 28800 9272 28864
rect 9336 28800 9352 28864
rect 9416 28800 9424 28864
rect 9104 28799 9424 28800
rect 10133 28794 10199 28797
rect 11200 28794 12000 28824
rect 0 28734 1456 28794
rect 0 28704 800 28734
rect 1396 28658 1456 28734
rect 10133 28792 12000 28794
rect 10133 28736 10138 28792
rect 10194 28736 12000 28792
rect 10133 28734 12000 28736
rect 10133 28731 10199 28734
rect 11200 28704 12000 28734
rect 2957 28658 3023 28661
rect 1396 28656 3023 28658
rect 1396 28600 2962 28656
rect 3018 28600 3023 28656
rect 1396 28598 3023 28600
rect 2957 28595 3023 28598
rect 0 28386 800 28416
rect 3325 28386 3391 28389
rect 0 28384 3391 28386
rect 0 28328 3330 28384
rect 3386 28328 3391 28384
rect 0 28326 3391 28328
rect 0 28296 800 28326
rect 3325 28323 3391 28326
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 7472 28320 7792 28321
rect 7472 28256 7480 28320
rect 7544 28256 7560 28320
rect 7624 28256 7640 28320
rect 7704 28256 7720 28320
rect 7784 28256 7792 28320
rect 7472 28255 7792 28256
rect 2078 28188 2084 28252
rect 2148 28250 2154 28252
rect 3969 28250 4035 28253
rect 5441 28250 5507 28253
rect 2148 28248 4035 28250
rect 2148 28192 3974 28248
rect 4030 28192 4035 28248
rect 2148 28190 4035 28192
rect 2148 28188 2154 28190
rect 3969 28187 4035 28190
rect 5168 28248 5507 28250
rect 5168 28192 5446 28248
rect 5502 28192 5507 28248
rect 5168 28190 5507 28192
rect 4245 28114 4311 28117
rect 5022 28114 5028 28116
rect 4245 28112 5028 28114
rect 4245 28056 4250 28112
rect 4306 28056 5028 28112
rect 4245 28054 5028 28056
rect 4245 28051 4311 28054
rect 5022 28052 5028 28054
rect 5092 28052 5098 28116
rect 0 27978 800 28008
rect 5168 27981 5228 28190
rect 5441 28187 5507 28190
rect 1209 27978 1275 27981
rect 0 27976 1275 27978
rect 0 27920 1214 27976
rect 1270 27920 1275 27976
rect 0 27918 1275 27920
rect 0 27888 800 27918
rect 1209 27915 1275 27918
rect 5165 27976 5231 27981
rect 5165 27920 5170 27976
rect 5226 27920 5231 27976
rect 5165 27915 5231 27920
rect 9949 27978 10015 27981
rect 11200 27978 12000 28008
rect 9949 27976 12000 27978
rect 9949 27920 9954 27976
rect 10010 27920 12000 27976
rect 9949 27918 12000 27920
rect 9949 27915 10015 27918
rect 11200 27888 12000 27918
rect 2576 27776 2896 27777
rect 2576 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2576 27711 2896 27712
rect 5840 27776 6160 27777
rect 5840 27712 5848 27776
rect 5912 27712 5928 27776
rect 5992 27712 6008 27776
rect 6072 27712 6088 27776
rect 6152 27712 6160 27776
rect 5840 27711 6160 27712
rect 9104 27776 9424 27777
rect 9104 27712 9112 27776
rect 9176 27712 9192 27776
rect 9256 27712 9272 27776
rect 9336 27712 9352 27776
rect 9416 27712 9424 27776
rect 9104 27711 9424 27712
rect 3366 27706 3372 27708
rect 3190 27646 3372 27706
rect 2773 27630 2839 27633
rect 3190 27630 3250 27646
rect 3366 27644 3372 27646
rect 3436 27644 3442 27708
rect 2773 27628 3250 27630
rect 0 27570 800 27600
rect 1393 27570 1459 27573
rect 0 27568 1459 27570
rect 0 27512 1398 27568
rect 1454 27512 1459 27568
rect 2773 27572 2778 27628
rect 2834 27572 3250 27628
rect 2773 27570 3250 27572
rect 2773 27567 2839 27570
rect 0 27510 1459 27512
rect 0 27480 800 27510
rect 1393 27507 1459 27510
rect 3550 27508 3556 27572
rect 3620 27570 3626 27572
rect 4245 27570 4311 27573
rect 3620 27568 4311 27570
rect 3620 27512 4250 27568
rect 4306 27512 4311 27568
rect 3620 27510 4311 27512
rect 3620 27508 3626 27510
rect 4245 27507 4311 27510
rect 3366 27372 3372 27436
rect 3436 27434 3442 27436
rect 4429 27434 4495 27437
rect 3436 27432 4495 27434
rect 3436 27376 4434 27432
rect 4490 27376 4495 27432
rect 3436 27374 4495 27376
rect 3436 27372 3442 27374
rect 4429 27371 4495 27374
rect 4208 27232 4528 27233
rect 0 27162 800 27192
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 7472 27232 7792 27233
rect 7472 27168 7480 27232
rect 7544 27168 7560 27232
rect 7624 27168 7640 27232
rect 7704 27168 7720 27232
rect 7784 27168 7792 27232
rect 7472 27167 7792 27168
rect 3601 27162 3667 27165
rect 0 27160 3667 27162
rect 0 27104 3606 27160
rect 3662 27104 3667 27160
rect 0 27102 3667 27104
rect 0 27072 800 27102
rect 3601 27099 3667 27102
rect 9949 27162 10015 27165
rect 11200 27162 12000 27192
rect 9949 27160 12000 27162
rect 9949 27104 9954 27160
rect 10010 27104 12000 27160
rect 9949 27102 12000 27104
rect 9949 27099 10015 27102
rect 11200 27072 12000 27102
rect 1853 26890 1919 26893
rect 1853 26888 1962 26890
rect 1853 26832 1858 26888
rect 1914 26832 1962 26888
rect 1853 26827 1962 26832
rect 1902 26754 1962 26827
rect 2129 26754 2195 26757
rect 1902 26752 2195 26754
rect 1902 26696 2134 26752
rect 2190 26696 2195 26752
rect 1902 26694 2195 26696
rect 2129 26691 2195 26694
rect 2576 26688 2896 26689
rect 0 26618 800 26648
rect 2576 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2576 26623 2896 26624
rect 5840 26688 6160 26689
rect 5840 26624 5848 26688
rect 5912 26624 5928 26688
rect 5992 26624 6008 26688
rect 6072 26624 6088 26688
rect 6152 26624 6160 26688
rect 5840 26623 6160 26624
rect 9104 26688 9424 26689
rect 9104 26624 9112 26688
rect 9176 26624 9192 26688
rect 9256 26624 9272 26688
rect 9336 26624 9352 26688
rect 9416 26624 9424 26688
rect 9104 26623 9424 26624
rect 0 26558 1456 26618
rect 0 26528 800 26558
rect 1396 26482 1456 26558
rect 3601 26482 3667 26485
rect 1396 26480 3667 26482
rect 1396 26424 3606 26480
rect 3662 26424 3667 26480
rect 1396 26422 3667 26424
rect 3601 26419 3667 26422
rect 10133 26482 10199 26485
rect 11200 26482 12000 26512
rect 10133 26480 12000 26482
rect 10133 26424 10138 26480
rect 10194 26424 12000 26480
rect 10133 26422 12000 26424
rect 10133 26419 10199 26422
rect 11200 26392 12000 26422
rect 0 26210 800 26240
rect 3509 26210 3575 26213
rect 0 26208 3575 26210
rect 0 26152 3514 26208
rect 3570 26152 3575 26208
rect 0 26150 3575 26152
rect 0 26120 800 26150
rect 3509 26147 3575 26150
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 7472 26144 7792 26145
rect 7472 26080 7480 26144
rect 7544 26080 7560 26144
rect 7624 26080 7640 26144
rect 7704 26080 7720 26144
rect 7784 26080 7792 26144
rect 7472 26079 7792 26080
rect 4521 25938 4587 25941
rect 5206 25938 5212 25940
rect 4521 25936 5212 25938
rect 4521 25880 4526 25936
rect 4582 25880 5212 25936
rect 4521 25878 5212 25880
rect 4521 25875 4587 25878
rect 5206 25876 5212 25878
rect 5276 25876 5282 25940
rect 0 25802 800 25832
rect 2589 25802 2655 25805
rect 0 25800 2655 25802
rect 0 25744 2594 25800
rect 2650 25744 2655 25800
rect 0 25742 2655 25744
rect 0 25712 800 25742
rect 2589 25739 2655 25742
rect 10133 25666 10199 25669
rect 11200 25666 12000 25696
rect 10133 25664 12000 25666
rect 10133 25608 10138 25664
rect 10194 25608 12000 25664
rect 10133 25606 12000 25608
rect 10133 25603 10199 25606
rect 2576 25600 2896 25601
rect 2576 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2576 25535 2896 25536
rect 5840 25600 6160 25601
rect 5840 25536 5848 25600
rect 5912 25536 5928 25600
rect 5992 25536 6008 25600
rect 6072 25536 6088 25600
rect 6152 25536 6160 25600
rect 5840 25535 6160 25536
rect 9104 25600 9424 25601
rect 9104 25536 9112 25600
rect 9176 25536 9192 25600
rect 9256 25536 9272 25600
rect 9336 25536 9352 25600
rect 9416 25536 9424 25600
rect 11200 25576 12000 25606
rect 9104 25535 9424 25536
rect 0 25394 800 25424
rect 1393 25394 1459 25397
rect 0 25392 1459 25394
rect 0 25336 1398 25392
rect 1454 25336 1459 25392
rect 0 25334 1459 25336
rect 0 25304 800 25334
rect 1393 25331 1459 25334
rect 3601 25258 3667 25261
rect 3734 25258 3740 25260
rect 3601 25256 3740 25258
rect 3601 25200 3606 25256
rect 3662 25200 3740 25256
rect 3601 25198 3740 25200
rect 3601 25195 3667 25198
rect 3734 25196 3740 25198
rect 3804 25196 3810 25260
rect 4208 25056 4528 25057
rect 0 24986 800 25016
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 7472 25056 7792 25057
rect 7472 24992 7480 25056
rect 7544 24992 7560 25056
rect 7624 24992 7640 25056
rect 7704 24992 7720 25056
rect 7784 24992 7792 25056
rect 7472 24991 7792 24992
rect 1393 24986 1459 24989
rect 0 24984 1459 24986
rect 0 24928 1398 24984
rect 1454 24928 1459 24984
rect 0 24926 1459 24928
rect 0 24896 800 24926
rect 1393 24923 1459 24926
rect 2773 24850 2839 24853
rect 3182 24850 3188 24852
rect 2773 24848 3188 24850
rect 2773 24792 2778 24848
rect 2834 24792 3188 24848
rect 2773 24790 3188 24792
rect 2773 24787 2839 24790
rect 3182 24788 3188 24790
rect 3252 24788 3258 24852
rect 10133 24850 10199 24853
rect 11200 24850 12000 24880
rect 10133 24848 12000 24850
rect 10133 24792 10138 24848
rect 10194 24792 12000 24848
rect 10133 24790 12000 24792
rect 10133 24787 10199 24790
rect 11200 24760 12000 24790
rect 3325 24714 3391 24717
rect 1396 24712 3391 24714
rect 1396 24656 3330 24712
rect 3386 24656 3391 24712
rect 1396 24654 3391 24656
rect 0 24578 800 24608
rect 1396 24578 1456 24654
rect 3325 24651 3391 24654
rect 0 24518 1456 24578
rect 3417 24578 3483 24581
rect 3918 24578 3924 24580
rect 3417 24576 3924 24578
rect 3417 24520 3422 24576
rect 3478 24520 3924 24576
rect 3417 24518 3924 24520
rect 0 24488 800 24518
rect 3417 24515 3483 24518
rect 3918 24516 3924 24518
rect 3988 24516 3994 24580
rect 2576 24512 2896 24513
rect 2576 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2576 24447 2896 24448
rect 5840 24512 6160 24513
rect 5840 24448 5848 24512
rect 5912 24448 5928 24512
rect 5992 24448 6008 24512
rect 6072 24448 6088 24512
rect 6152 24448 6160 24512
rect 5840 24447 6160 24448
rect 9104 24512 9424 24513
rect 9104 24448 9112 24512
rect 9176 24448 9192 24512
rect 9256 24448 9272 24512
rect 9336 24448 9352 24512
rect 9416 24448 9424 24512
rect 9104 24447 9424 24448
rect 0 24170 800 24200
rect 2957 24170 3023 24173
rect 0 24168 3023 24170
rect 0 24112 2962 24168
rect 3018 24112 3023 24168
rect 0 24110 3023 24112
rect 0 24080 800 24110
rect 2957 24107 3023 24110
rect 10133 24170 10199 24173
rect 11200 24170 12000 24200
rect 10133 24168 12000 24170
rect 10133 24112 10138 24168
rect 10194 24112 12000 24168
rect 10133 24110 12000 24112
rect 10133 24107 10199 24110
rect 11200 24080 12000 24110
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 7472 23968 7792 23969
rect 7472 23904 7480 23968
rect 7544 23904 7560 23968
rect 7624 23904 7640 23968
rect 7704 23904 7720 23968
rect 7784 23904 7792 23968
rect 7472 23903 7792 23904
rect 1761 23898 1827 23901
rect 2262 23898 2268 23900
rect 1761 23896 2268 23898
rect 1761 23840 1766 23896
rect 1822 23840 2268 23896
rect 1761 23838 2268 23840
rect 1761 23835 1827 23838
rect 2262 23836 2268 23838
rect 2332 23836 2338 23900
rect 0 23626 800 23656
rect 2773 23626 2839 23629
rect 0 23624 2839 23626
rect 0 23568 2778 23624
rect 2834 23568 2839 23624
rect 0 23566 2839 23568
rect 0 23536 800 23566
rect 2773 23563 2839 23566
rect 2576 23424 2896 23425
rect 2576 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2576 23359 2896 23360
rect 5840 23424 6160 23425
rect 5840 23360 5848 23424
rect 5912 23360 5928 23424
rect 5992 23360 6008 23424
rect 6072 23360 6088 23424
rect 6152 23360 6160 23424
rect 5840 23359 6160 23360
rect 9104 23424 9424 23425
rect 9104 23360 9112 23424
rect 9176 23360 9192 23424
rect 9256 23360 9272 23424
rect 9336 23360 9352 23424
rect 9416 23360 9424 23424
rect 9104 23359 9424 23360
rect 10133 23354 10199 23357
rect 11200 23354 12000 23384
rect 10133 23352 12000 23354
rect 10133 23296 10138 23352
rect 10194 23296 12000 23352
rect 10133 23294 12000 23296
rect 10133 23291 10199 23294
rect 11200 23264 12000 23294
rect 0 23218 800 23248
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 800 23158
rect 1393 23155 1459 23158
rect 4208 22880 4528 22881
rect 0 22810 800 22840
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 7472 22880 7792 22881
rect 7472 22816 7480 22880
rect 7544 22816 7560 22880
rect 7624 22816 7640 22880
rect 7704 22816 7720 22880
rect 7784 22816 7792 22880
rect 7472 22815 7792 22816
rect 1209 22810 1275 22813
rect 0 22808 1275 22810
rect 0 22752 1214 22808
rect 1270 22752 1275 22808
rect 0 22750 1275 22752
rect 0 22720 800 22750
rect 1209 22747 1275 22750
rect 3049 22810 3115 22813
rect 3366 22810 3372 22812
rect 3049 22808 3372 22810
rect 3049 22752 3054 22808
rect 3110 22752 3372 22808
rect 3049 22750 3372 22752
rect 3049 22747 3115 22750
rect 3366 22748 3372 22750
rect 3436 22748 3442 22812
rect 3785 22674 3851 22677
rect 3742 22672 3851 22674
rect 3742 22616 3790 22672
rect 3846 22616 3851 22672
rect 3742 22611 3851 22616
rect 0 22402 800 22432
rect 3742 22405 3802 22611
rect 10133 22538 10199 22541
rect 11200 22538 12000 22568
rect 10133 22536 12000 22538
rect 10133 22480 10138 22536
rect 10194 22480 12000 22536
rect 10133 22478 12000 22480
rect 10133 22475 10199 22478
rect 11200 22448 12000 22478
rect 1393 22402 1459 22405
rect 0 22400 1459 22402
rect 0 22344 1398 22400
rect 1454 22344 1459 22400
rect 0 22342 1459 22344
rect 3742 22400 3851 22405
rect 3742 22344 3790 22400
rect 3846 22344 3851 22400
rect 3742 22342 3851 22344
rect 0 22312 800 22342
rect 1393 22339 1459 22342
rect 3785 22339 3851 22342
rect 2576 22336 2896 22337
rect 2576 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2576 22271 2896 22272
rect 5840 22336 6160 22337
rect 5840 22272 5848 22336
rect 5912 22272 5928 22336
rect 5992 22272 6008 22336
rect 6072 22272 6088 22336
rect 6152 22272 6160 22336
rect 5840 22271 6160 22272
rect 9104 22336 9424 22337
rect 9104 22272 9112 22336
rect 9176 22272 9192 22336
rect 9256 22272 9272 22336
rect 9336 22272 9352 22336
rect 9416 22272 9424 22336
rect 9104 22271 9424 22272
rect 2313 22268 2379 22269
rect 2262 22204 2268 22268
rect 2332 22266 2379 22268
rect 2332 22264 2424 22266
rect 2374 22208 2424 22264
rect 2332 22206 2424 22208
rect 2332 22204 2379 22206
rect 3550 22204 3556 22268
rect 3620 22266 3626 22268
rect 3693 22266 3759 22269
rect 3620 22264 3759 22266
rect 3620 22208 3698 22264
rect 3754 22208 3759 22264
rect 3620 22206 3759 22208
rect 3620 22204 3626 22206
rect 2313 22203 2379 22204
rect 3693 22203 3759 22206
rect 2037 22130 2103 22133
rect 2497 22130 2563 22133
rect 2037 22128 2563 22130
rect 2037 22072 2042 22128
rect 2098 22072 2502 22128
rect 2558 22072 2563 22128
rect 2037 22070 2563 22072
rect 2037 22067 2103 22070
rect 2497 22067 2563 22070
rect 0 21994 800 22024
rect 1209 21994 1275 21997
rect 0 21992 1275 21994
rect 0 21936 1214 21992
rect 1270 21936 1275 21992
rect 0 21934 1275 21936
rect 0 21904 800 21934
rect 1209 21931 1275 21934
rect 2221 21996 2287 21997
rect 2221 21992 2268 21996
rect 2332 21994 2338 21996
rect 2221 21936 2226 21992
rect 2221 21932 2268 21936
rect 2332 21934 2378 21994
rect 2332 21932 2338 21934
rect 2221 21931 2287 21932
rect 10133 21858 10199 21861
rect 11200 21858 12000 21888
rect 10133 21856 12000 21858
rect 10133 21800 10138 21856
rect 10194 21800 12000 21856
rect 10133 21798 12000 21800
rect 10133 21795 10199 21798
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 7472 21792 7792 21793
rect 7472 21728 7480 21792
rect 7544 21728 7560 21792
rect 7624 21728 7640 21792
rect 7704 21728 7720 21792
rect 7784 21728 7792 21792
rect 11200 21768 12000 21798
rect 7472 21727 7792 21728
rect 0 21586 800 21616
rect 1393 21586 1459 21589
rect 0 21584 1459 21586
rect 0 21528 1398 21584
rect 1454 21528 1459 21584
rect 0 21526 1459 21528
rect 0 21496 800 21526
rect 1393 21523 1459 21526
rect 2576 21248 2896 21249
rect 0 21178 800 21208
rect 2576 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2576 21183 2896 21184
rect 5840 21248 6160 21249
rect 5840 21184 5848 21248
rect 5912 21184 5928 21248
rect 5992 21184 6008 21248
rect 6072 21184 6088 21248
rect 6152 21184 6160 21248
rect 5840 21183 6160 21184
rect 9104 21248 9424 21249
rect 9104 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9272 21248
rect 9336 21184 9352 21248
rect 9416 21184 9424 21248
rect 9104 21183 9424 21184
rect 1393 21178 1459 21181
rect 0 21176 1459 21178
rect 0 21120 1398 21176
rect 1454 21120 1459 21176
rect 0 21118 1459 21120
rect 0 21088 800 21118
rect 1393 21115 1459 21118
rect 10133 21042 10199 21045
rect 11200 21042 12000 21072
rect 10133 21040 12000 21042
rect 10133 20984 10138 21040
rect 10194 20984 12000 21040
rect 10133 20982 12000 20984
rect 10133 20979 10199 20982
rect 11200 20952 12000 20982
rect 4208 20704 4528 20705
rect 0 20634 800 20664
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 7472 20704 7792 20705
rect 7472 20640 7480 20704
rect 7544 20640 7560 20704
rect 7624 20640 7640 20704
rect 7704 20640 7720 20704
rect 7784 20640 7792 20704
rect 7472 20639 7792 20640
rect 1393 20634 1459 20637
rect 0 20632 1459 20634
rect 0 20576 1398 20632
rect 1454 20576 1459 20632
rect 0 20574 1459 20576
rect 0 20544 800 20574
rect 1393 20571 1459 20574
rect 10041 20362 10107 20365
rect 11200 20362 12000 20392
rect 10041 20360 12000 20362
rect 10041 20304 10046 20360
rect 10102 20304 12000 20360
rect 10041 20302 12000 20304
rect 10041 20299 10107 20302
rect 11200 20272 12000 20302
rect 0 20226 800 20256
rect 1393 20226 1459 20229
rect 0 20224 1459 20226
rect 0 20168 1398 20224
rect 1454 20168 1459 20224
rect 0 20166 1459 20168
rect 0 20136 800 20166
rect 1393 20163 1459 20166
rect 2576 20160 2896 20161
rect 2576 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2576 20095 2896 20096
rect 5840 20160 6160 20161
rect 5840 20096 5848 20160
rect 5912 20096 5928 20160
rect 5992 20096 6008 20160
rect 6072 20096 6088 20160
rect 6152 20096 6160 20160
rect 5840 20095 6160 20096
rect 9104 20160 9424 20161
rect 9104 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9272 20160
rect 9336 20096 9352 20160
rect 9416 20096 9424 20160
rect 9104 20095 9424 20096
rect 0 19818 800 19848
rect 3969 19818 4035 19821
rect 0 19816 4035 19818
rect 0 19760 3974 19816
rect 4030 19760 4035 19816
rect 0 19758 4035 19760
rect 0 19728 800 19758
rect 3969 19755 4035 19758
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 7472 19616 7792 19617
rect 7472 19552 7480 19616
rect 7544 19552 7560 19616
rect 7624 19552 7640 19616
rect 7704 19552 7720 19616
rect 7784 19552 7792 19616
rect 7472 19551 7792 19552
rect 10041 19546 10107 19549
rect 11200 19546 12000 19576
rect 10041 19544 12000 19546
rect 10041 19488 10046 19544
rect 10102 19488 12000 19544
rect 10041 19486 12000 19488
rect 10041 19483 10107 19486
rect 11200 19456 12000 19486
rect 0 19410 800 19440
rect 2865 19410 2931 19413
rect 0 19408 2931 19410
rect 0 19352 2870 19408
rect 2926 19352 2931 19408
rect 0 19350 2931 19352
rect 0 19320 800 19350
rect 2865 19347 2931 19350
rect 2773 19274 2839 19277
rect 1396 19272 2839 19274
rect 1396 19216 2778 19272
rect 2834 19216 2839 19272
rect 1396 19214 2839 19216
rect 0 19002 800 19032
rect 1396 19002 1456 19214
rect 2773 19211 2839 19214
rect 2576 19072 2896 19073
rect 2576 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2576 19007 2896 19008
rect 5840 19072 6160 19073
rect 5840 19008 5848 19072
rect 5912 19008 5928 19072
rect 5992 19008 6008 19072
rect 6072 19008 6088 19072
rect 6152 19008 6160 19072
rect 5840 19007 6160 19008
rect 9104 19072 9424 19073
rect 9104 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9272 19072
rect 9336 19008 9352 19072
rect 9416 19008 9424 19072
rect 9104 19007 9424 19008
rect 0 18942 1456 19002
rect 0 18912 800 18942
rect 10041 18730 10107 18733
rect 11200 18730 12000 18760
rect 10041 18728 12000 18730
rect 10041 18672 10046 18728
rect 10102 18672 12000 18728
rect 10041 18670 12000 18672
rect 10041 18667 10107 18670
rect 11200 18640 12000 18670
rect 0 18594 800 18624
rect 2865 18594 2931 18597
rect 0 18592 2931 18594
rect 0 18536 2870 18592
rect 2926 18536 2931 18592
rect 0 18534 2931 18536
rect 0 18504 800 18534
rect 2865 18531 2931 18534
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 7472 18528 7792 18529
rect 7472 18464 7480 18528
rect 7544 18464 7560 18528
rect 7624 18464 7640 18528
rect 7704 18464 7720 18528
rect 7784 18464 7792 18528
rect 7472 18463 7792 18464
rect 0 18186 800 18216
rect 2221 18186 2287 18189
rect 0 18184 2287 18186
rect 0 18128 2226 18184
rect 2282 18128 2287 18184
rect 0 18126 2287 18128
rect 0 18096 800 18126
rect 2221 18123 2287 18126
rect 10041 18050 10107 18053
rect 11200 18050 12000 18080
rect 10041 18048 12000 18050
rect 10041 17992 10046 18048
rect 10102 17992 12000 18048
rect 10041 17990 12000 17992
rect 10041 17987 10107 17990
rect 2576 17984 2896 17985
rect 2576 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2576 17919 2896 17920
rect 5840 17984 6160 17985
rect 5840 17920 5848 17984
rect 5912 17920 5928 17984
rect 5992 17920 6008 17984
rect 6072 17920 6088 17984
rect 6152 17920 6160 17984
rect 5840 17919 6160 17920
rect 9104 17984 9424 17985
rect 9104 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9272 17984
rect 9336 17920 9352 17984
rect 9416 17920 9424 17984
rect 11200 17960 12000 17990
rect 9104 17919 9424 17920
rect 0 17642 800 17672
rect 1485 17642 1551 17645
rect 0 17640 1551 17642
rect 0 17584 1490 17640
rect 1546 17584 1551 17640
rect 0 17582 1551 17584
rect 0 17552 800 17582
rect 1485 17579 1551 17582
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 7472 17440 7792 17441
rect 7472 17376 7480 17440
rect 7544 17376 7560 17440
rect 7624 17376 7640 17440
rect 7704 17376 7720 17440
rect 7784 17376 7792 17440
rect 7472 17375 7792 17376
rect 0 17234 800 17264
rect 1393 17234 1459 17237
rect 0 17232 1459 17234
rect 0 17176 1398 17232
rect 1454 17176 1459 17232
rect 0 17174 1459 17176
rect 0 17144 800 17174
rect 1393 17171 1459 17174
rect 10041 17234 10107 17237
rect 11200 17234 12000 17264
rect 10041 17232 12000 17234
rect 10041 17176 10046 17232
rect 10102 17176 12000 17232
rect 10041 17174 12000 17176
rect 10041 17171 10107 17174
rect 11200 17144 12000 17174
rect 2576 16896 2896 16897
rect 0 16826 800 16856
rect 2576 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2576 16831 2896 16832
rect 5840 16896 6160 16897
rect 5840 16832 5848 16896
rect 5912 16832 5928 16896
rect 5992 16832 6008 16896
rect 6072 16832 6088 16896
rect 6152 16832 6160 16896
rect 5840 16831 6160 16832
rect 9104 16896 9424 16897
rect 9104 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9272 16896
rect 9336 16832 9352 16896
rect 9416 16832 9424 16896
rect 9104 16831 9424 16832
rect 1577 16826 1643 16829
rect 0 16824 1643 16826
rect 0 16768 1582 16824
rect 1638 16768 1643 16824
rect 0 16766 1643 16768
rect 0 16736 800 16766
rect 1577 16763 1643 16766
rect 0 16418 800 16448
rect 3969 16418 4035 16421
rect 0 16416 4035 16418
rect 0 16360 3974 16416
rect 4030 16360 4035 16416
rect 0 16358 4035 16360
rect 0 16328 800 16358
rect 3969 16355 4035 16358
rect 10041 16418 10107 16421
rect 11200 16418 12000 16448
rect 10041 16416 12000 16418
rect 10041 16360 10046 16416
rect 10102 16360 12000 16416
rect 10041 16358 12000 16360
rect 10041 16355 10107 16358
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 7472 16352 7792 16353
rect 7472 16288 7480 16352
rect 7544 16288 7560 16352
rect 7624 16288 7640 16352
rect 7704 16288 7720 16352
rect 7784 16288 7792 16352
rect 11200 16328 12000 16358
rect 7472 16287 7792 16288
rect 0 16010 800 16040
rect 2773 16010 2839 16013
rect 0 16008 2839 16010
rect 0 15952 2778 16008
rect 2834 15952 2839 16008
rect 0 15950 2839 15952
rect 0 15920 800 15950
rect 2773 15947 2839 15950
rect 2576 15808 2896 15809
rect 2576 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2576 15743 2896 15744
rect 5840 15808 6160 15809
rect 5840 15744 5848 15808
rect 5912 15744 5928 15808
rect 5992 15744 6008 15808
rect 6072 15744 6088 15808
rect 6152 15744 6160 15808
rect 5840 15743 6160 15744
rect 9104 15808 9424 15809
rect 9104 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9272 15808
rect 9336 15744 9352 15808
rect 9416 15744 9424 15808
rect 9104 15743 9424 15744
rect 10041 15738 10107 15741
rect 11200 15738 12000 15768
rect 10041 15736 12000 15738
rect 10041 15680 10046 15736
rect 10102 15680 12000 15736
rect 10041 15678 12000 15680
rect 10041 15675 10107 15678
rect 11200 15648 12000 15678
rect 0 15602 800 15632
rect 1485 15602 1551 15605
rect 0 15600 1551 15602
rect 0 15544 1490 15600
rect 1546 15544 1551 15600
rect 0 15542 1551 15544
rect 0 15512 800 15542
rect 1485 15539 1551 15542
rect 4208 15264 4528 15265
rect 0 15194 800 15224
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 7472 15264 7792 15265
rect 7472 15200 7480 15264
rect 7544 15200 7560 15264
rect 7624 15200 7640 15264
rect 7704 15200 7720 15264
rect 7784 15200 7792 15264
rect 7472 15199 7792 15200
rect 3969 15194 4035 15197
rect 0 15192 4035 15194
rect 0 15136 3974 15192
rect 4030 15136 4035 15192
rect 0 15134 4035 15136
rect 0 15104 800 15134
rect 3969 15131 4035 15134
rect 3141 15058 3207 15061
rect 5574 15058 5580 15060
rect 3141 15056 5580 15058
rect 3141 15000 3146 15056
rect 3202 15000 5580 15056
rect 3141 14998 5580 15000
rect 3141 14995 3207 14998
rect 5574 14996 5580 14998
rect 5644 14996 5650 15060
rect 2865 14922 2931 14925
rect 1396 14920 2931 14922
rect 1396 14864 2870 14920
rect 2926 14864 2931 14920
rect 1396 14862 2931 14864
rect 0 14650 800 14680
rect 1396 14650 1456 14862
rect 2865 14859 2931 14862
rect 10041 14922 10107 14925
rect 11200 14922 12000 14952
rect 10041 14920 12000 14922
rect 10041 14864 10046 14920
rect 10102 14864 12000 14920
rect 10041 14862 12000 14864
rect 10041 14859 10107 14862
rect 11200 14832 12000 14862
rect 1669 14786 1735 14789
rect 1669 14784 1778 14786
rect 1669 14728 1674 14784
rect 1730 14728 1778 14784
rect 1669 14723 1778 14728
rect 0 14590 1456 14650
rect 0 14560 800 14590
rect 1718 14378 1778 14723
rect 2576 14720 2896 14721
rect 2576 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2576 14655 2896 14656
rect 5840 14720 6160 14721
rect 5840 14656 5848 14720
rect 5912 14656 5928 14720
rect 5992 14656 6008 14720
rect 6072 14656 6088 14720
rect 6152 14656 6160 14720
rect 5840 14655 6160 14656
rect 9104 14720 9424 14721
rect 9104 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9272 14720
rect 9336 14656 9352 14720
rect 9416 14656 9424 14720
rect 9104 14655 9424 14656
rect 1945 14378 2011 14381
rect 1718 14376 2011 14378
rect 1718 14320 1950 14376
rect 2006 14320 2011 14376
rect 1718 14318 2011 14320
rect 1945 14315 2011 14318
rect 0 14242 800 14272
rect 3969 14242 4035 14245
rect 0 14240 4035 14242
rect 0 14184 3974 14240
rect 4030 14184 4035 14240
rect 0 14182 4035 14184
rect 0 14152 800 14182
rect 3969 14179 4035 14182
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 7472 14176 7792 14177
rect 7472 14112 7480 14176
rect 7544 14112 7560 14176
rect 7624 14112 7640 14176
rect 7704 14112 7720 14176
rect 7784 14112 7792 14176
rect 7472 14111 7792 14112
rect 10041 14106 10107 14109
rect 11200 14106 12000 14136
rect 10041 14104 12000 14106
rect 10041 14048 10046 14104
rect 10102 14048 12000 14104
rect 10041 14046 12000 14048
rect 10041 14043 10107 14046
rect 11200 14016 12000 14046
rect 0 13834 800 13864
rect 3969 13834 4035 13837
rect 0 13832 4035 13834
rect 0 13776 3974 13832
rect 4030 13776 4035 13832
rect 0 13774 4035 13776
rect 0 13744 800 13774
rect 3969 13771 4035 13774
rect 2576 13632 2896 13633
rect 2576 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2576 13567 2896 13568
rect 5840 13632 6160 13633
rect 5840 13568 5848 13632
rect 5912 13568 5928 13632
rect 5992 13568 6008 13632
rect 6072 13568 6088 13632
rect 6152 13568 6160 13632
rect 5840 13567 6160 13568
rect 9104 13632 9424 13633
rect 9104 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9272 13632
rect 9336 13568 9352 13632
rect 9416 13568 9424 13632
rect 9104 13567 9424 13568
rect 0 13426 800 13456
rect 3877 13426 3943 13429
rect 0 13424 3943 13426
rect 0 13368 3882 13424
rect 3938 13368 3943 13424
rect 0 13366 3943 13368
rect 0 13336 800 13366
rect 3877 13363 3943 13366
rect 9581 13426 9647 13429
rect 11200 13426 12000 13456
rect 9581 13424 12000 13426
rect 9581 13368 9586 13424
rect 9642 13368 12000 13424
rect 9581 13366 12000 13368
rect 9581 13363 9647 13366
rect 11200 13336 12000 13366
rect 1894 13092 1900 13156
rect 1964 13154 1970 13156
rect 2037 13154 2103 13157
rect 1964 13152 2103 13154
rect 1964 13096 2042 13152
rect 2098 13096 2103 13152
rect 1964 13094 2103 13096
rect 1964 13092 1970 13094
rect 2037 13091 2103 13094
rect 4208 13088 4528 13089
rect 0 13018 800 13048
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 7472 13088 7792 13089
rect 7472 13024 7480 13088
rect 7544 13024 7560 13088
rect 7624 13024 7640 13088
rect 7704 13024 7720 13088
rect 7784 13024 7792 13088
rect 7472 13023 7792 13024
rect 3233 13018 3299 13021
rect 0 13016 3299 13018
rect 0 12960 3238 13016
rect 3294 12960 3299 13016
rect 0 12958 3299 12960
rect 0 12928 800 12958
rect 3233 12955 3299 12958
rect 0 12610 800 12640
rect 1577 12610 1643 12613
rect 0 12608 1643 12610
rect 0 12552 1582 12608
rect 1638 12552 1643 12608
rect 0 12550 1643 12552
rect 0 12520 800 12550
rect 1577 12547 1643 12550
rect 10041 12610 10107 12613
rect 11200 12610 12000 12640
rect 10041 12608 12000 12610
rect 10041 12552 10046 12608
rect 10102 12552 12000 12608
rect 10041 12550 12000 12552
rect 10041 12547 10107 12550
rect 2576 12544 2896 12545
rect 2576 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2576 12479 2896 12480
rect 5840 12544 6160 12545
rect 5840 12480 5848 12544
rect 5912 12480 5928 12544
rect 5992 12480 6008 12544
rect 6072 12480 6088 12544
rect 6152 12480 6160 12544
rect 5840 12479 6160 12480
rect 9104 12544 9424 12545
rect 9104 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9272 12544
rect 9336 12480 9352 12544
rect 9416 12480 9424 12544
rect 11200 12520 12000 12550
rect 9104 12479 9424 12480
rect 1894 12412 1900 12476
rect 1964 12412 1970 12476
rect 1577 12338 1643 12341
rect 1902 12338 1962 12412
rect 1577 12336 1962 12338
rect 1577 12280 1582 12336
rect 1638 12280 1962 12336
rect 1577 12278 1962 12280
rect 1577 12275 1643 12278
rect 0 12202 800 12232
rect 3233 12202 3299 12205
rect 0 12200 3299 12202
rect 0 12144 3238 12200
rect 3294 12144 3299 12200
rect 0 12142 3299 12144
rect 0 12112 800 12142
rect 3233 12139 3299 12142
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 7472 12000 7792 12001
rect 7472 11936 7480 12000
rect 7544 11936 7560 12000
rect 7624 11936 7640 12000
rect 7704 11936 7720 12000
rect 7784 11936 7792 12000
rect 7472 11935 7792 11936
rect 1301 11794 1367 11797
rect 798 11792 1367 11794
rect 798 11736 1306 11792
rect 1362 11736 1367 11792
rect 798 11734 1367 11736
rect 798 11688 858 11734
rect 1301 11731 1367 11734
rect 10041 11794 10107 11797
rect 11200 11794 12000 11824
rect 10041 11792 12000 11794
rect 10041 11736 10046 11792
rect 10102 11736 12000 11792
rect 10041 11734 12000 11736
rect 10041 11731 10107 11734
rect 11200 11704 12000 11734
rect 0 11598 858 11688
rect 0 11568 800 11598
rect 2576 11456 2896 11457
rect 2576 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2576 11391 2896 11392
rect 5840 11456 6160 11457
rect 5840 11392 5848 11456
rect 5912 11392 5928 11456
rect 5992 11392 6008 11456
rect 6072 11392 6088 11456
rect 6152 11392 6160 11456
rect 5840 11391 6160 11392
rect 9104 11456 9424 11457
rect 9104 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9272 11456
rect 9336 11392 9352 11456
rect 9416 11392 9424 11456
rect 9104 11391 9424 11392
rect 0 11250 800 11280
rect 1209 11250 1275 11253
rect 0 11248 1275 11250
rect 0 11192 1214 11248
rect 1270 11192 1275 11248
rect 0 11190 1275 11192
rect 0 11160 800 11190
rect 1209 11187 1275 11190
rect 10041 11114 10107 11117
rect 11200 11114 12000 11144
rect 10041 11112 12000 11114
rect 10041 11056 10046 11112
rect 10102 11056 12000 11112
rect 10041 11054 12000 11056
rect 10041 11051 10107 11054
rect 11200 11024 12000 11054
rect 4208 10912 4528 10913
rect 0 10842 800 10872
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 7472 10912 7792 10913
rect 7472 10848 7480 10912
rect 7544 10848 7560 10912
rect 7624 10848 7640 10912
rect 7704 10848 7720 10912
rect 7784 10848 7792 10912
rect 7472 10847 7792 10848
rect 1301 10842 1367 10845
rect 0 10840 1367 10842
rect 0 10784 1306 10840
rect 1362 10784 1367 10840
rect 0 10782 1367 10784
rect 0 10752 800 10782
rect 1301 10779 1367 10782
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 2576 10368 2896 10369
rect 2576 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2576 10303 2896 10304
rect 5840 10368 6160 10369
rect 5840 10304 5848 10368
rect 5912 10304 5928 10368
rect 5992 10304 6008 10368
rect 6072 10304 6088 10368
rect 6152 10304 6160 10368
rect 5840 10303 6160 10304
rect 9104 10368 9424 10369
rect 9104 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9272 10368
rect 9336 10304 9352 10368
rect 9416 10304 9424 10368
rect 9104 10303 9424 10304
rect 10041 10298 10107 10301
rect 11200 10298 12000 10328
rect 10041 10296 12000 10298
rect 10041 10240 10046 10296
rect 10102 10240 12000 10296
rect 10041 10238 12000 10240
rect 10041 10235 10107 10238
rect 11200 10208 12000 10238
rect 0 10026 800 10056
rect 1301 10026 1367 10029
rect 0 10024 1367 10026
rect 0 9968 1306 10024
rect 1362 9968 1367 10024
rect 0 9966 1367 9968
rect 0 9936 800 9966
rect 1301 9963 1367 9966
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 7472 9824 7792 9825
rect 7472 9760 7480 9824
rect 7544 9760 7560 9824
rect 7624 9760 7640 9824
rect 7704 9760 7720 9824
rect 7784 9760 7792 9824
rect 7472 9759 7792 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 2865 9482 2931 9485
rect 4838 9482 4844 9484
rect 2865 9480 4844 9482
rect 2865 9424 2870 9480
rect 2926 9424 4844 9480
rect 2865 9422 4844 9424
rect 2865 9419 2931 9422
rect 4838 9420 4844 9422
rect 4908 9420 4914 9484
rect 10041 9482 10107 9485
rect 11200 9482 12000 9512
rect 10041 9480 12000 9482
rect 10041 9424 10046 9480
rect 10102 9424 12000 9480
rect 10041 9422 12000 9424
rect 10041 9419 10107 9422
rect 11200 9392 12000 9422
rect 2576 9280 2896 9281
rect 0 9210 800 9240
rect 2576 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2576 9215 2896 9216
rect 5840 9280 6160 9281
rect 5840 9216 5848 9280
rect 5912 9216 5928 9280
rect 5992 9216 6008 9280
rect 6072 9216 6088 9280
rect 6152 9216 6160 9280
rect 5840 9215 6160 9216
rect 9104 9280 9424 9281
rect 9104 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9272 9280
rect 9336 9216 9352 9280
rect 9416 9216 9424 9280
rect 9104 9215 9424 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 2957 9212 3023 9213
rect 2957 9208 3004 9212
rect 3068 9210 3074 9212
rect 2957 9152 2962 9208
rect 2957 9148 3004 9152
rect 3068 9150 3114 9210
rect 3068 9148 3074 9150
rect 2957 9147 3023 9148
rect 3969 9074 4035 9077
rect 3742 9072 4035 9074
rect 3742 9016 3974 9072
rect 4030 9016 4035 9072
rect 3742 9014 4035 9016
rect 0 8666 800 8696
rect 1393 8666 1459 8669
rect 0 8664 1459 8666
rect 0 8608 1398 8664
rect 1454 8608 1459 8664
rect 0 8606 1459 8608
rect 0 8576 800 8606
rect 1393 8603 1459 8606
rect 3742 8533 3802 9014
rect 3969 9011 4035 9014
rect 10041 8802 10107 8805
rect 11200 8802 12000 8832
rect 10041 8800 12000 8802
rect 10041 8744 10046 8800
rect 10102 8744 12000 8800
rect 10041 8742 12000 8744
rect 10041 8739 10107 8742
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 7472 8736 7792 8737
rect 7472 8672 7480 8736
rect 7544 8672 7560 8736
rect 7624 8672 7640 8736
rect 7704 8672 7720 8736
rect 7784 8672 7792 8736
rect 11200 8712 12000 8742
rect 7472 8671 7792 8672
rect 3693 8528 3802 8533
rect 3693 8472 3698 8528
rect 3754 8472 3802 8528
rect 3693 8470 3802 8472
rect 3693 8467 3759 8470
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 2576 8192 2896 8193
rect 2576 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2576 8127 2896 8128
rect 5840 8192 6160 8193
rect 5840 8128 5848 8192
rect 5912 8128 5928 8192
rect 5992 8128 6008 8192
rect 6072 8128 6088 8192
rect 6152 8128 6160 8192
rect 5840 8127 6160 8128
rect 9104 8192 9424 8193
rect 9104 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9272 8192
rect 9336 8128 9352 8192
rect 9416 8128 9424 8192
rect 9104 8127 9424 8128
rect 10041 7986 10107 7989
rect 11200 7986 12000 8016
rect 10041 7984 12000 7986
rect 10041 7928 10046 7984
rect 10102 7928 12000 7984
rect 10041 7926 12000 7928
rect 10041 7923 10107 7926
rect 11200 7896 12000 7926
rect 0 7850 800 7880
rect 1393 7850 1459 7853
rect 0 7848 1459 7850
rect 0 7792 1398 7848
rect 1454 7792 1459 7848
rect 0 7790 1459 7792
rect 0 7760 800 7790
rect 1393 7787 1459 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 7472 7648 7792 7649
rect 7472 7584 7480 7648
rect 7544 7584 7560 7648
rect 7624 7584 7640 7648
rect 7704 7584 7720 7648
rect 7784 7584 7792 7648
rect 7472 7583 7792 7584
rect 0 7442 800 7472
rect 1393 7442 1459 7445
rect 0 7440 1459 7442
rect 0 7384 1398 7440
rect 1454 7384 1459 7440
rect 0 7382 1459 7384
rect 0 7352 800 7382
rect 1393 7379 1459 7382
rect 10041 7170 10107 7173
rect 11200 7170 12000 7200
rect 10041 7168 12000 7170
rect 10041 7112 10046 7168
rect 10102 7112 12000 7168
rect 10041 7110 12000 7112
rect 10041 7107 10107 7110
rect 2576 7104 2896 7105
rect 0 7034 800 7064
rect 2576 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2576 7039 2896 7040
rect 5840 7104 6160 7105
rect 5840 7040 5848 7104
rect 5912 7040 5928 7104
rect 5992 7040 6008 7104
rect 6072 7040 6088 7104
rect 6152 7040 6160 7104
rect 5840 7039 6160 7040
rect 9104 7104 9424 7105
rect 9104 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9272 7104
rect 9336 7040 9352 7104
rect 9416 7040 9424 7104
rect 11200 7080 12000 7110
rect 9104 7039 9424 7040
rect 2221 7034 2287 7037
rect 0 7032 2287 7034
rect 0 6976 2226 7032
rect 2282 6976 2287 7032
rect 0 6974 2287 6976
rect 0 6944 800 6974
rect 2221 6971 2287 6974
rect 974 6700 980 6764
rect 1044 6762 1050 6764
rect 1577 6762 1643 6765
rect 1044 6760 1643 6762
rect 1044 6704 1582 6760
rect 1638 6704 1643 6760
rect 1044 6702 1643 6704
rect 1044 6700 1050 6702
rect 1577 6699 1643 6702
rect 0 6626 800 6656
rect 2221 6626 2287 6629
rect 0 6624 2287 6626
rect 0 6568 2226 6624
rect 2282 6568 2287 6624
rect 0 6566 2287 6568
rect 0 6536 800 6566
rect 2221 6563 2287 6566
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 7472 6560 7792 6561
rect 7472 6496 7480 6560
rect 7544 6496 7560 6560
rect 7624 6496 7640 6560
rect 7704 6496 7720 6560
rect 7784 6496 7792 6560
rect 7472 6495 7792 6496
rect 10041 6490 10107 6493
rect 11200 6490 12000 6520
rect 10041 6488 12000 6490
rect 10041 6432 10046 6488
rect 10102 6432 12000 6488
rect 10041 6430 12000 6432
rect 10041 6427 10107 6430
rect 11200 6400 12000 6430
rect 0 6218 800 6248
rect 1853 6218 1919 6221
rect 0 6216 1919 6218
rect 0 6160 1858 6216
rect 1914 6160 1919 6216
rect 0 6158 1919 6160
rect 0 6128 800 6158
rect 1853 6155 1919 6158
rect 2576 6016 2896 6017
rect 2576 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2576 5951 2896 5952
rect 5840 6016 6160 6017
rect 5840 5952 5848 6016
rect 5912 5952 5928 6016
rect 5992 5952 6008 6016
rect 6072 5952 6088 6016
rect 6152 5952 6160 6016
rect 5840 5951 6160 5952
rect 9104 6016 9424 6017
rect 9104 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9272 6016
rect 9336 5952 9352 6016
rect 9416 5952 9424 6016
rect 9104 5951 9424 5952
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 10041 5674 10107 5677
rect 11200 5674 12000 5704
rect 10041 5672 12000 5674
rect 10041 5616 10046 5672
rect 10102 5616 12000 5672
rect 10041 5614 12000 5616
rect 10041 5611 10107 5614
rect 11200 5584 12000 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 7472 5472 7792 5473
rect 7472 5408 7480 5472
rect 7544 5408 7560 5472
rect 7624 5408 7640 5472
rect 7704 5408 7720 5472
rect 7784 5408 7792 5472
rect 7472 5407 7792 5408
rect 0 5266 800 5296
rect 1393 5266 1459 5269
rect 0 5264 1459 5266
rect 0 5208 1398 5264
rect 1454 5208 1459 5264
rect 0 5206 1459 5208
rect 0 5176 800 5206
rect 1393 5203 1459 5206
rect 3693 5266 3759 5269
rect 8334 5266 8340 5268
rect 3693 5264 8340 5266
rect 3693 5208 3698 5264
rect 3754 5208 8340 5264
rect 3693 5206 8340 5208
rect 3693 5203 3759 5206
rect 8334 5204 8340 5206
rect 8404 5204 8410 5268
rect 2576 4928 2896 4929
rect 0 4858 800 4888
rect 2576 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2576 4863 2896 4864
rect 5840 4928 6160 4929
rect 5840 4864 5848 4928
rect 5912 4864 5928 4928
rect 5992 4864 6008 4928
rect 6072 4864 6088 4928
rect 6152 4864 6160 4928
rect 5840 4863 6160 4864
rect 9104 4928 9424 4929
rect 9104 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9272 4928
rect 9336 4864 9352 4928
rect 9416 4864 9424 4928
rect 9104 4863 9424 4864
rect 3969 4858 4035 4861
rect 4654 4858 4660 4860
rect 0 4798 1410 4858
rect 0 4768 800 4798
rect 1350 4722 1410 4798
rect 3969 4856 4660 4858
rect 3969 4800 3974 4856
rect 4030 4800 4660 4856
rect 3969 4798 4660 4800
rect 3969 4795 4035 4798
rect 4654 4796 4660 4798
rect 4724 4796 4730 4860
rect 10041 4858 10107 4861
rect 11200 4858 12000 4888
rect 10041 4856 12000 4858
rect 10041 4800 10046 4856
rect 10102 4800 12000 4856
rect 10041 4798 12000 4800
rect 10041 4795 10107 4798
rect 11200 4768 12000 4798
rect 3325 4722 3391 4725
rect 1350 4720 3391 4722
rect 1350 4664 3330 4720
rect 3386 4664 3391 4720
rect 1350 4662 3391 4664
rect 3325 4659 3391 4662
rect 0 4450 800 4480
rect 2957 4450 3023 4453
rect 0 4448 3023 4450
rect 0 4392 2962 4448
rect 3018 4392 3023 4448
rect 0 4390 3023 4392
rect 0 4360 800 4390
rect 2957 4387 3023 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 7472 4384 7792 4385
rect 7472 4320 7480 4384
rect 7544 4320 7560 4384
rect 7624 4320 7640 4384
rect 7704 4320 7720 4384
rect 7784 4320 7792 4384
rect 7472 4319 7792 4320
rect 10041 4178 10107 4181
rect 11200 4178 12000 4208
rect 10041 4176 12000 4178
rect 10041 4120 10046 4176
rect 10102 4120 12000 4176
rect 10041 4118 12000 4120
rect 10041 4115 10107 4118
rect 11200 4088 12000 4118
rect 0 4042 800 4072
rect 1393 4042 1459 4045
rect 0 4040 1459 4042
rect 0 3984 1398 4040
rect 1454 3984 1459 4040
rect 0 3982 1459 3984
rect 0 3952 800 3982
rect 1393 3979 1459 3982
rect 2576 3840 2896 3841
rect 2576 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2576 3775 2896 3776
rect 5840 3840 6160 3841
rect 5840 3776 5848 3840
rect 5912 3776 5928 3840
rect 5992 3776 6008 3840
rect 6072 3776 6088 3840
rect 6152 3776 6160 3840
rect 5840 3775 6160 3776
rect 9104 3840 9424 3841
rect 9104 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9272 3840
rect 9336 3776 9352 3840
rect 9416 3776 9424 3840
rect 9104 3775 9424 3776
rect 0 3634 800 3664
rect 2957 3634 3023 3637
rect 0 3632 3023 3634
rect 0 3576 2962 3632
rect 3018 3576 3023 3632
rect 0 3574 3023 3576
rect 0 3544 800 3574
rect 2957 3571 3023 3574
rect 10041 3362 10107 3365
rect 11200 3362 12000 3392
rect 10041 3360 12000 3362
rect 10041 3304 10046 3360
rect 10102 3304 12000 3360
rect 10041 3302 12000 3304
rect 10041 3299 10107 3302
rect 4208 3296 4528 3297
rect 0 3226 800 3256
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 7472 3296 7792 3297
rect 7472 3232 7480 3296
rect 7544 3232 7560 3296
rect 7624 3232 7640 3296
rect 7704 3232 7720 3296
rect 7784 3232 7792 3296
rect 11200 3272 12000 3302
rect 7472 3231 7792 3232
rect 2313 3226 2379 3229
rect 0 3224 2379 3226
rect 0 3168 2318 3224
rect 2374 3168 2379 3224
rect 0 3166 2379 3168
rect 0 3136 800 3166
rect 2313 3163 2379 3166
rect 2576 2752 2896 2753
rect 0 2682 800 2712
rect 2576 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2576 2687 2896 2688
rect 5840 2752 6160 2753
rect 5840 2688 5848 2752
rect 5912 2688 5928 2752
rect 5992 2688 6008 2752
rect 6072 2688 6088 2752
rect 6152 2688 6160 2752
rect 5840 2687 6160 2688
rect 9104 2752 9424 2753
rect 9104 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9272 2752
rect 9336 2688 9352 2752
rect 9416 2688 9424 2752
rect 9104 2687 9424 2688
rect 0 2622 2514 2682
rect 0 2592 800 2622
rect 2454 2546 2514 2622
rect 4061 2546 4127 2549
rect 2454 2544 4127 2546
rect 2454 2488 4066 2544
rect 4122 2488 4127 2544
rect 2454 2486 4127 2488
rect 4061 2483 4127 2486
rect 10041 2546 10107 2549
rect 11200 2546 12000 2576
rect 10041 2544 12000 2546
rect 10041 2488 10046 2544
rect 10102 2488 12000 2544
rect 10041 2486 12000 2488
rect 10041 2483 10107 2486
rect 11200 2456 12000 2486
rect 0 2274 800 2304
rect 2773 2274 2839 2277
rect 0 2272 2839 2274
rect 0 2216 2778 2272
rect 2834 2216 2839 2272
rect 0 2214 2839 2216
rect 0 2184 800 2214
rect 2773 2211 2839 2214
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 7472 2208 7792 2209
rect 7472 2144 7480 2208
rect 7544 2144 7560 2208
rect 7624 2144 7640 2208
rect 7704 2144 7720 2208
rect 7784 2144 7792 2208
rect 7472 2143 7792 2144
rect 0 1866 800 1896
rect 4061 1866 4127 1869
rect 0 1864 4127 1866
rect 0 1808 4066 1864
rect 4122 1808 4127 1864
rect 0 1806 4127 1808
rect 0 1776 800 1806
rect 4061 1803 4127 1806
rect 9489 1866 9555 1869
rect 11200 1866 12000 1896
rect 9489 1864 12000 1866
rect 9489 1808 9494 1864
rect 9550 1808 12000 1864
rect 9489 1806 12000 1808
rect 9489 1803 9555 1806
rect 11200 1776 12000 1806
rect 0 1458 800 1488
rect 3969 1458 4035 1461
rect 0 1456 4035 1458
rect 0 1400 3974 1456
rect 4030 1400 4035 1456
rect 0 1398 4035 1400
rect 0 1368 800 1398
rect 3969 1395 4035 1398
rect 0 1050 800 1080
rect 2773 1050 2839 1053
rect 0 1048 2839 1050
rect 0 992 2778 1048
rect 2834 992 2839 1048
rect 0 990 2839 992
rect 0 960 800 990
rect 2773 987 2839 990
rect 9581 1050 9647 1053
rect 11200 1050 12000 1080
rect 9581 1048 12000 1050
rect 9581 992 9586 1048
rect 9642 992 12000 1048
rect 9581 990 12000 992
rect 9581 987 9647 990
rect 11200 960 12000 990
rect 0 642 800 672
rect 2865 642 2931 645
rect 0 640 2931 642
rect 0 584 2870 640
rect 2926 584 2931 640
rect 0 582 2931 584
rect 0 552 800 582
rect 2865 579 2931 582
rect 9305 370 9371 373
rect 11200 370 12000 400
rect 9305 368 12000 370
rect 9305 312 9310 368
rect 9366 312 12000 368
rect 9305 310 12000 312
rect 9305 307 9371 310
rect 11200 280 12000 310
rect 0 234 800 264
rect 1393 234 1459 237
rect 0 232 1459 234
rect 0 176 1398 232
rect 1454 176 1459 232
rect 0 174 1459 176
rect 0 144 800 174
rect 1393 171 1459 174
<< via3 >>
rect 2584 77820 2648 77824
rect 2584 77764 2588 77820
rect 2588 77764 2644 77820
rect 2644 77764 2648 77820
rect 2584 77760 2648 77764
rect 2664 77820 2728 77824
rect 2664 77764 2668 77820
rect 2668 77764 2724 77820
rect 2724 77764 2728 77820
rect 2664 77760 2728 77764
rect 2744 77820 2808 77824
rect 2744 77764 2748 77820
rect 2748 77764 2804 77820
rect 2804 77764 2808 77820
rect 2744 77760 2808 77764
rect 2824 77820 2888 77824
rect 2824 77764 2828 77820
rect 2828 77764 2884 77820
rect 2884 77764 2888 77820
rect 2824 77760 2888 77764
rect 5848 77820 5912 77824
rect 5848 77764 5852 77820
rect 5852 77764 5908 77820
rect 5908 77764 5912 77820
rect 5848 77760 5912 77764
rect 5928 77820 5992 77824
rect 5928 77764 5932 77820
rect 5932 77764 5988 77820
rect 5988 77764 5992 77820
rect 5928 77760 5992 77764
rect 6008 77820 6072 77824
rect 6008 77764 6012 77820
rect 6012 77764 6068 77820
rect 6068 77764 6072 77820
rect 6008 77760 6072 77764
rect 6088 77820 6152 77824
rect 6088 77764 6092 77820
rect 6092 77764 6148 77820
rect 6148 77764 6152 77820
rect 6088 77760 6152 77764
rect 9112 77820 9176 77824
rect 9112 77764 9116 77820
rect 9116 77764 9172 77820
rect 9172 77764 9176 77820
rect 9112 77760 9176 77764
rect 9192 77820 9256 77824
rect 9192 77764 9196 77820
rect 9196 77764 9252 77820
rect 9252 77764 9256 77820
rect 9192 77760 9256 77764
rect 9272 77820 9336 77824
rect 9272 77764 9276 77820
rect 9276 77764 9332 77820
rect 9332 77764 9336 77820
rect 9272 77760 9336 77764
rect 9352 77820 9416 77824
rect 9352 77764 9356 77820
rect 9356 77764 9412 77820
rect 9412 77764 9416 77820
rect 9352 77760 9416 77764
rect 4216 77276 4280 77280
rect 4216 77220 4220 77276
rect 4220 77220 4276 77276
rect 4276 77220 4280 77276
rect 4216 77216 4280 77220
rect 4296 77276 4360 77280
rect 4296 77220 4300 77276
rect 4300 77220 4356 77276
rect 4356 77220 4360 77276
rect 4296 77216 4360 77220
rect 4376 77276 4440 77280
rect 4376 77220 4380 77276
rect 4380 77220 4436 77276
rect 4436 77220 4440 77276
rect 4376 77216 4440 77220
rect 4456 77276 4520 77280
rect 4456 77220 4460 77276
rect 4460 77220 4516 77276
rect 4516 77220 4520 77276
rect 4456 77216 4520 77220
rect 7480 77276 7544 77280
rect 7480 77220 7484 77276
rect 7484 77220 7540 77276
rect 7540 77220 7544 77276
rect 7480 77216 7544 77220
rect 7560 77276 7624 77280
rect 7560 77220 7564 77276
rect 7564 77220 7620 77276
rect 7620 77220 7624 77276
rect 7560 77216 7624 77220
rect 7640 77276 7704 77280
rect 7640 77220 7644 77276
rect 7644 77220 7700 77276
rect 7700 77220 7704 77276
rect 7640 77216 7704 77220
rect 7720 77276 7784 77280
rect 7720 77220 7724 77276
rect 7724 77220 7780 77276
rect 7780 77220 7784 77276
rect 7720 77216 7784 77220
rect 2584 76732 2648 76736
rect 2584 76676 2588 76732
rect 2588 76676 2644 76732
rect 2644 76676 2648 76732
rect 2584 76672 2648 76676
rect 2664 76732 2728 76736
rect 2664 76676 2668 76732
rect 2668 76676 2724 76732
rect 2724 76676 2728 76732
rect 2664 76672 2728 76676
rect 2744 76732 2808 76736
rect 2744 76676 2748 76732
rect 2748 76676 2804 76732
rect 2804 76676 2808 76732
rect 2744 76672 2808 76676
rect 2824 76732 2888 76736
rect 2824 76676 2828 76732
rect 2828 76676 2884 76732
rect 2884 76676 2888 76732
rect 2824 76672 2888 76676
rect 5848 76732 5912 76736
rect 5848 76676 5852 76732
rect 5852 76676 5908 76732
rect 5908 76676 5912 76732
rect 5848 76672 5912 76676
rect 5928 76732 5992 76736
rect 5928 76676 5932 76732
rect 5932 76676 5988 76732
rect 5988 76676 5992 76732
rect 5928 76672 5992 76676
rect 6008 76732 6072 76736
rect 6008 76676 6012 76732
rect 6012 76676 6068 76732
rect 6068 76676 6072 76732
rect 6008 76672 6072 76676
rect 6088 76732 6152 76736
rect 6088 76676 6092 76732
rect 6092 76676 6148 76732
rect 6148 76676 6152 76732
rect 6088 76672 6152 76676
rect 9112 76732 9176 76736
rect 9112 76676 9116 76732
rect 9116 76676 9172 76732
rect 9172 76676 9176 76732
rect 9112 76672 9176 76676
rect 9192 76732 9256 76736
rect 9192 76676 9196 76732
rect 9196 76676 9252 76732
rect 9252 76676 9256 76732
rect 9192 76672 9256 76676
rect 9272 76732 9336 76736
rect 9272 76676 9276 76732
rect 9276 76676 9332 76732
rect 9332 76676 9336 76732
rect 9272 76672 9336 76676
rect 9352 76732 9416 76736
rect 9352 76676 9356 76732
rect 9356 76676 9412 76732
rect 9412 76676 9416 76732
rect 9352 76672 9416 76676
rect 4216 76188 4280 76192
rect 4216 76132 4220 76188
rect 4220 76132 4276 76188
rect 4276 76132 4280 76188
rect 4216 76128 4280 76132
rect 4296 76188 4360 76192
rect 4296 76132 4300 76188
rect 4300 76132 4356 76188
rect 4356 76132 4360 76188
rect 4296 76128 4360 76132
rect 4376 76188 4440 76192
rect 4376 76132 4380 76188
rect 4380 76132 4436 76188
rect 4436 76132 4440 76188
rect 4376 76128 4440 76132
rect 4456 76188 4520 76192
rect 4456 76132 4460 76188
rect 4460 76132 4516 76188
rect 4516 76132 4520 76188
rect 4456 76128 4520 76132
rect 7480 76188 7544 76192
rect 7480 76132 7484 76188
rect 7484 76132 7540 76188
rect 7540 76132 7544 76188
rect 7480 76128 7544 76132
rect 7560 76188 7624 76192
rect 7560 76132 7564 76188
rect 7564 76132 7620 76188
rect 7620 76132 7624 76188
rect 7560 76128 7624 76132
rect 7640 76188 7704 76192
rect 7640 76132 7644 76188
rect 7644 76132 7700 76188
rect 7700 76132 7704 76188
rect 7640 76128 7704 76132
rect 7720 76188 7784 76192
rect 7720 76132 7724 76188
rect 7724 76132 7780 76188
rect 7780 76132 7784 76188
rect 7720 76128 7784 76132
rect 2584 75644 2648 75648
rect 2584 75588 2588 75644
rect 2588 75588 2644 75644
rect 2644 75588 2648 75644
rect 2584 75584 2648 75588
rect 2664 75644 2728 75648
rect 2664 75588 2668 75644
rect 2668 75588 2724 75644
rect 2724 75588 2728 75644
rect 2664 75584 2728 75588
rect 2744 75644 2808 75648
rect 2744 75588 2748 75644
rect 2748 75588 2804 75644
rect 2804 75588 2808 75644
rect 2744 75584 2808 75588
rect 2824 75644 2888 75648
rect 2824 75588 2828 75644
rect 2828 75588 2884 75644
rect 2884 75588 2888 75644
rect 2824 75584 2888 75588
rect 5848 75644 5912 75648
rect 5848 75588 5852 75644
rect 5852 75588 5908 75644
rect 5908 75588 5912 75644
rect 5848 75584 5912 75588
rect 5928 75644 5992 75648
rect 5928 75588 5932 75644
rect 5932 75588 5988 75644
rect 5988 75588 5992 75644
rect 5928 75584 5992 75588
rect 6008 75644 6072 75648
rect 6008 75588 6012 75644
rect 6012 75588 6068 75644
rect 6068 75588 6072 75644
rect 6008 75584 6072 75588
rect 6088 75644 6152 75648
rect 6088 75588 6092 75644
rect 6092 75588 6148 75644
rect 6148 75588 6152 75644
rect 6088 75584 6152 75588
rect 9112 75644 9176 75648
rect 9112 75588 9116 75644
rect 9116 75588 9172 75644
rect 9172 75588 9176 75644
rect 9112 75584 9176 75588
rect 9192 75644 9256 75648
rect 9192 75588 9196 75644
rect 9196 75588 9252 75644
rect 9252 75588 9256 75644
rect 9192 75584 9256 75588
rect 9272 75644 9336 75648
rect 9272 75588 9276 75644
rect 9276 75588 9332 75644
rect 9332 75588 9336 75644
rect 9272 75584 9336 75588
rect 9352 75644 9416 75648
rect 9352 75588 9356 75644
rect 9356 75588 9412 75644
rect 9412 75588 9416 75644
rect 9352 75584 9416 75588
rect 4216 75100 4280 75104
rect 4216 75044 4220 75100
rect 4220 75044 4276 75100
rect 4276 75044 4280 75100
rect 4216 75040 4280 75044
rect 4296 75100 4360 75104
rect 4296 75044 4300 75100
rect 4300 75044 4356 75100
rect 4356 75044 4360 75100
rect 4296 75040 4360 75044
rect 4376 75100 4440 75104
rect 4376 75044 4380 75100
rect 4380 75044 4436 75100
rect 4436 75044 4440 75100
rect 4376 75040 4440 75044
rect 4456 75100 4520 75104
rect 4456 75044 4460 75100
rect 4460 75044 4516 75100
rect 4516 75044 4520 75100
rect 4456 75040 4520 75044
rect 7480 75100 7544 75104
rect 7480 75044 7484 75100
rect 7484 75044 7540 75100
rect 7540 75044 7544 75100
rect 7480 75040 7544 75044
rect 7560 75100 7624 75104
rect 7560 75044 7564 75100
rect 7564 75044 7620 75100
rect 7620 75044 7624 75100
rect 7560 75040 7624 75044
rect 7640 75100 7704 75104
rect 7640 75044 7644 75100
rect 7644 75044 7700 75100
rect 7700 75044 7704 75100
rect 7640 75040 7704 75044
rect 7720 75100 7784 75104
rect 7720 75044 7724 75100
rect 7724 75044 7780 75100
rect 7780 75044 7784 75100
rect 7720 75040 7784 75044
rect 3924 74972 3988 75036
rect 2584 74556 2648 74560
rect 2584 74500 2588 74556
rect 2588 74500 2644 74556
rect 2644 74500 2648 74556
rect 2584 74496 2648 74500
rect 2664 74556 2728 74560
rect 2664 74500 2668 74556
rect 2668 74500 2724 74556
rect 2724 74500 2728 74556
rect 2664 74496 2728 74500
rect 2744 74556 2808 74560
rect 2744 74500 2748 74556
rect 2748 74500 2804 74556
rect 2804 74500 2808 74556
rect 2744 74496 2808 74500
rect 2824 74556 2888 74560
rect 2824 74500 2828 74556
rect 2828 74500 2884 74556
rect 2884 74500 2888 74556
rect 2824 74496 2888 74500
rect 5848 74556 5912 74560
rect 5848 74500 5852 74556
rect 5852 74500 5908 74556
rect 5908 74500 5912 74556
rect 5848 74496 5912 74500
rect 5928 74556 5992 74560
rect 5928 74500 5932 74556
rect 5932 74500 5988 74556
rect 5988 74500 5992 74556
rect 5928 74496 5992 74500
rect 6008 74556 6072 74560
rect 6008 74500 6012 74556
rect 6012 74500 6068 74556
rect 6068 74500 6072 74556
rect 6008 74496 6072 74500
rect 6088 74556 6152 74560
rect 6088 74500 6092 74556
rect 6092 74500 6148 74556
rect 6148 74500 6152 74556
rect 6088 74496 6152 74500
rect 9112 74556 9176 74560
rect 9112 74500 9116 74556
rect 9116 74500 9172 74556
rect 9172 74500 9176 74556
rect 9112 74496 9176 74500
rect 9192 74556 9256 74560
rect 9192 74500 9196 74556
rect 9196 74500 9252 74556
rect 9252 74500 9256 74556
rect 9192 74496 9256 74500
rect 9272 74556 9336 74560
rect 9272 74500 9276 74556
rect 9276 74500 9332 74556
rect 9332 74500 9336 74556
rect 9272 74496 9336 74500
rect 9352 74556 9416 74560
rect 9352 74500 9356 74556
rect 9356 74500 9412 74556
rect 9412 74500 9416 74556
rect 9352 74496 9416 74500
rect 4216 74012 4280 74016
rect 4216 73956 4220 74012
rect 4220 73956 4276 74012
rect 4276 73956 4280 74012
rect 4216 73952 4280 73956
rect 4296 74012 4360 74016
rect 4296 73956 4300 74012
rect 4300 73956 4356 74012
rect 4356 73956 4360 74012
rect 4296 73952 4360 73956
rect 4376 74012 4440 74016
rect 4376 73956 4380 74012
rect 4380 73956 4436 74012
rect 4436 73956 4440 74012
rect 4376 73952 4440 73956
rect 4456 74012 4520 74016
rect 4456 73956 4460 74012
rect 4460 73956 4516 74012
rect 4516 73956 4520 74012
rect 4456 73952 4520 73956
rect 7480 74012 7544 74016
rect 7480 73956 7484 74012
rect 7484 73956 7540 74012
rect 7540 73956 7544 74012
rect 7480 73952 7544 73956
rect 7560 74012 7624 74016
rect 7560 73956 7564 74012
rect 7564 73956 7620 74012
rect 7620 73956 7624 74012
rect 7560 73952 7624 73956
rect 7640 74012 7704 74016
rect 7640 73956 7644 74012
rect 7644 73956 7700 74012
rect 7700 73956 7704 74012
rect 7640 73952 7704 73956
rect 7720 74012 7784 74016
rect 7720 73956 7724 74012
rect 7724 73956 7780 74012
rect 7780 73956 7784 74012
rect 7720 73952 7784 73956
rect 2584 73468 2648 73472
rect 2584 73412 2588 73468
rect 2588 73412 2644 73468
rect 2644 73412 2648 73468
rect 2584 73408 2648 73412
rect 2664 73468 2728 73472
rect 2664 73412 2668 73468
rect 2668 73412 2724 73468
rect 2724 73412 2728 73468
rect 2664 73408 2728 73412
rect 2744 73468 2808 73472
rect 2744 73412 2748 73468
rect 2748 73412 2804 73468
rect 2804 73412 2808 73468
rect 2744 73408 2808 73412
rect 2824 73468 2888 73472
rect 2824 73412 2828 73468
rect 2828 73412 2884 73468
rect 2884 73412 2888 73468
rect 2824 73408 2888 73412
rect 5848 73468 5912 73472
rect 5848 73412 5852 73468
rect 5852 73412 5908 73468
rect 5908 73412 5912 73468
rect 5848 73408 5912 73412
rect 5928 73468 5992 73472
rect 5928 73412 5932 73468
rect 5932 73412 5988 73468
rect 5988 73412 5992 73468
rect 5928 73408 5992 73412
rect 6008 73468 6072 73472
rect 6008 73412 6012 73468
rect 6012 73412 6068 73468
rect 6068 73412 6072 73468
rect 6008 73408 6072 73412
rect 6088 73468 6152 73472
rect 6088 73412 6092 73468
rect 6092 73412 6148 73468
rect 6148 73412 6152 73468
rect 6088 73408 6152 73412
rect 9112 73468 9176 73472
rect 9112 73412 9116 73468
rect 9116 73412 9172 73468
rect 9172 73412 9176 73468
rect 9112 73408 9176 73412
rect 9192 73468 9256 73472
rect 9192 73412 9196 73468
rect 9196 73412 9252 73468
rect 9252 73412 9256 73468
rect 9192 73408 9256 73412
rect 9272 73468 9336 73472
rect 9272 73412 9276 73468
rect 9276 73412 9332 73468
rect 9332 73412 9336 73468
rect 9272 73408 9336 73412
rect 9352 73468 9416 73472
rect 9352 73412 9356 73468
rect 9356 73412 9412 73468
rect 9412 73412 9416 73468
rect 9352 73408 9416 73412
rect 4216 72924 4280 72928
rect 4216 72868 4220 72924
rect 4220 72868 4276 72924
rect 4276 72868 4280 72924
rect 4216 72864 4280 72868
rect 4296 72924 4360 72928
rect 4296 72868 4300 72924
rect 4300 72868 4356 72924
rect 4356 72868 4360 72924
rect 4296 72864 4360 72868
rect 4376 72924 4440 72928
rect 4376 72868 4380 72924
rect 4380 72868 4436 72924
rect 4436 72868 4440 72924
rect 4376 72864 4440 72868
rect 4456 72924 4520 72928
rect 4456 72868 4460 72924
rect 4460 72868 4516 72924
rect 4516 72868 4520 72924
rect 4456 72864 4520 72868
rect 7480 72924 7544 72928
rect 7480 72868 7484 72924
rect 7484 72868 7540 72924
rect 7540 72868 7544 72924
rect 7480 72864 7544 72868
rect 7560 72924 7624 72928
rect 7560 72868 7564 72924
rect 7564 72868 7620 72924
rect 7620 72868 7624 72924
rect 7560 72864 7624 72868
rect 7640 72924 7704 72928
rect 7640 72868 7644 72924
rect 7644 72868 7700 72924
rect 7700 72868 7704 72924
rect 7640 72864 7704 72868
rect 7720 72924 7784 72928
rect 7720 72868 7724 72924
rect 7724 72868 7780 72924
rect 7780 72868 7784 72924
rect 7720 72864 7784 72868
rect 2584 72380 2648 72384
rect 2584 72324 2588 72380
rect 2588 72324 2644 72380
rect 2644 72324 2648 72380
rect 2584 72320 2648 72324
rect 2664 72380 2728 72384
rect 2664 72324 2668 72380
rect 2668 72324 2724 72380
rect 2724 72324 2728 72380
rect 2664 72320 2728 72324
rect 2744 72380 2808 72384
rect 2744 72324 2748 72380
rect 2748 72324 2804 72380
rect 2804 72324 2808 72380
rect 2744 72320 2808 72324
rect 2824 72380 2888 72384
rect 2824 72324 2828 72380
rect 2828 72324 2884 72380
rect 2884 72324 2888 72380
rect 2824 72320 2888 72324
rect 5848 72380 5912 72384
rect 5848 72324 5852 72380
rect 5852 72324 5908 72380
rect 5908 72324 5912 72380
rect 5848 72320 5912 72324
rect 5928 72380 5992 72384
rect 5928 72324 5932 72380
rect 5932 72324 5988 72380
rect 5988 72324 5992 72380
rect 5928 72320 5992 72324
rect 6008 72380 6072 72384
rect 6008 72324 6012 72380
rect 6012 72324 6068 72380
rect 6068 72324 6072 72380
rect 6008 72320 6072 72324
rect 6088 72380 6152 72384
rect 6088 72324 6092 72380
rect 6092 72324 6148 72380
rect 6148 72324 6152 72380
rect 6088 72320 6152 72324
rect 9112 72380 9176 72384
rect 9112 72324 9116 72380
rect 9116 72324 9172 72380
rect 9172 72324 9176 72380
rect 9112 72320 9176 72324
rect 9192 72380 9256 72384
rect 9192 72324 9196 72380
rect 9196 72324 9252 72380
rect 9252 72324 9256 72380
rect 9192 72320 9256 72324
rect 9272 72380 9336 72384
rect 9272 72324 9276 72380
rect 9276 72324 9332 72380
rect 9332 72324 9336 72380
rect 9272 72320 9336 72324
rect 9352 72380 9416 72384
rect 9352 72324 9356 72380
rect 9356 72324 9412 72380
rect 9412 72324 9416 72380
rect 9352 72320 9416 72324
rect 4216 71836 4280 71840
rect 4216 71780 4220 71836
rect 4220 71780 4276 71836
rect 4276 71780 4280 71836
rect 4216 71776 4280 71780
rect 4296 71836 4360 71840
rect 4296 71780 4300 71836
rect 4300 71780 4356 71836
rect 4356 71780 4360 71836
rect 4296 71776 4360 71780
rect 4376 71836 4440 71840
rect 4376 71780 4380 71836
rect 4380 71780 4436 71836
rect 4436 71780 4440 71836
rect 4376 71776 4440 71780
rect 4456 71836 4520 71840
rect 4456 71780 4460 71836
rect 4460 71780 4516 71836
rect 4516 71780 4520 71836
rect 4456 71776 4520 71780
rect 7480 71836 7544 71840
rect 7480 71780 7484 71836
rect 7484 71780 7540 71836
rect 7540 71780 7544 71836
rect 7480 71776 7544 71780
rect 7560 71836 7624 71840
rect 7560 71780 7564 71836
rect 7564 71780 7620 71836
rect 7620 71780 7624 71836
rect 7560 71776 7624 71780
rect 7640 71836 7704 71840
rect 7640 71780 7644 71836
rect 7644 71780 7700 71836
rect 7700 71780 7704 71836
rect 7640 71776 7704 71780
rect 7720 71836 7784 71840
rect 7720 71780 7724 71836
rect 7724 71780 7780 71836
rect 7780 71780 7784 71836
rect 7720 71776 7784 71780
rect 2584 71292 2648 71296
rect 2584 71236 2588 71292
rect 2588 71236 2644 71292
rect 2644 71236 2648 71292
rect 2584 71232 2648 71236
rect 2664 71292 2728 71296
rect 2664 71236 2668 71292
rect 2668 71236 2724 71292
rect 2724 71236 2728 71292
rect 2664 71232 2728 71236
rect 2744 71292 2808 71296
rect 2744 71236 2748 71292
rect 2748 71236 2804 71292
rect 2804 71236 2808 71292
rect 2744 71232 2808 71236
rect 2824 71292 2888 71296
rect 2824 71236 2828 71292
rect 2828 71236 2884 71292
rect 2884 71236 2888 71292
rect 2824 71232 2888 71236
rect 5848 71292 5912 71296
rect 5848 71236 5852 71292
rect 5852 71236 5908 71292
rect 5908 71236 5912 71292
rect 5848 71232 5912 71236
rect 5928 71292 5992 71296
rect 5928 71236 5932 71292
rect 5932 71236 5988 71292
rect 5988 71236 5992 71292
rect 5928 71232 5992 71236
rect 6008 71292 6072 71296
rect 6008 71236 6012 71292
rect 6012 71236 6068 71292
rect 6068 71236 6072 71292
rect 6008 71232 6072 71236
rect 6088 71292 6152 71296
rect 6088 71236 6092 71292
rect 6092 71236 6148 71292
rect 6148 71236 6152 71292
rect 6088 71232 6152 71236
rect 9112 71292 9176 71296
rect 9112 71236 9116 71292
rect 9116 71236 9172 71292
rect 9172 71236 9176 71292
rect 9112 71232 9176 71236
rect 9192 71292 9256 71296
rect 9192 71236 9196 71292
rect 9196 71236 9252 71292
rect 9252 71236 9256 71292
rect 9192 71232 9256 71236
rect 9272 71292 9336 71296
rect 9272 71236 9276 71292
rect 9276 71236 9332 71292
rect 9332 71236 9336 71292
rect 9272 71232 9336 71236
rect 9352 71292 9416 71296
rect 9352 71236 9356 71292
rect 9356 71236 9412 71292
rect 9412 71236 9416 71292
rect 9352 71232 9416 71236
rect 4216 70748 4280 70752
rect 4216 70692 4220 70748
rect 4220 70692 4276 70748
rect 4276 70692 4280 70748
rect 4216 70688 4280 70692
rect 4296 70748 4360 70752
rect 4296 70692 4300 70748
rect 4300 70692 4356 70748
rect 4356 70692 4360 70748
rect 4296 70688 4360 70692
rect 4376 70748 4440 70752
rect 4376 70692 4380 70748
rect 4380 70692 4436 70748
rect 4436 70692 4440 70748
rect 4376 70688 4440 70692
rect 4456 70748 4520 70752
rect 4456 70692 4460 70748
rect 4460 70692 4516 70748
rect 4516 70692 4520 70748
rect 4456 70688 4520 70692
rect 7480 70748 7544 70752
rect 7480 70692 7484 70748
rect 7484 70692 7540 70748
rect 7540 70692 7544 70748
rect 7480 70688 7544 70692
rect 7560 70748 7624 70752
rect 7560 70692 7564 70748
rect 7564 70692 7620 70748
rect 7620 70692 7624 70748
rect 7560 70688 7624 70692
rect 7640 70748 7704 70752
rect 7640 70692 7644 70748
rect 7644 70692 7700 70748
rect 7700 70692 7704 70748
rect 7640 70688 7704 70692
rect 7720 70748 7784 70752
rect 7720 70692 7724 70748
rect 7724 70692 7780 70748
rect 7780 70692 7784 70748
rect 7720 70688 7784 70692
rect 2584 70204 2648 70208
rect 2584 70148 2588 70204
rect 2588 70148 2644 70204
rect 2644 70148 2648 70204
rect 2584 70144 2648 70148
rect 2664 70204 2728 70208
rect 2664 70148 2668 70204
rect 2668 70148 2724 70204
rect 2724 70148 2728 70204
rect 2664 70144 2728 70148
rect 2744 70204 2808 70208
rect 2744 70148 2748 70204
rect 2748 70148 2804 70204
rect 2804 70148 2808 70204
rect 2744 70144 2808 70148
rect 2824 70204 2888 70208
rect 2824 70148 2828 70204
rect 2828 70148 2884 70204
rect 2884 70148 2888 70204
rect 2824 70144 2888 70148
rect 5848 70204 5912 70208
rect 5848 70148 5852 70204
rect 5852 70148 5908 70204
rect 5908 70148 5912 70204
rect 5848 70144 5912 70148
rect 5928 70204 5992 70208
rect 5928 70148 5932 70204
rect 5932 70148 5988 70204
rect 5988 70148 5992 70204
rect 5928 70144 5992 70148
rect 6008 70204 6072 70208
rect 6008 70148 6012 70204
rect 6012 70148 6068 70204
rect 6068 70148 6072 70204
rect 6008 70144 6072 70148
rect 6088 70204 6152 70208
rect 6088 70148 6092 70204
rect 6092 70148 6148 70204
rect 6148 70148 6152 70204
rect 6088 70144 6152 70148
rect 9112 70204 9176 70208
rect 9112 70148 9116 70204
rect 9116 70148 9172 70204
rect 9172 70148 9176 70204
rect 9112 70144 9176 70148
rect 9192 70204 9256 70208
rect 9192 70148 9196 70204
rect 9196 70148 9252 70204
rect 9252 70148 9256 70204
rect 9192 70144 9256 70148
rect 9272 70204 9336 70208
rect 9272 70148 9276 70204
rect 9276 70148 9332 70204
rect 9332 70148 9336 70204
rect 9272 70144 9336 70148
rect 9352 70204 9416 70208
rect 9352 70148 9356 70204
rect 9356 70148 9412 70204
rect 9412 70148 9416 70204
rect 9352 70144 9416 70148
rect 4216 69660 4280 69664
rect 4216 69604 4220 69660
rect 4220 69604 4276 69660
rect 4276 69604 4280 69660
rect 4216 69600 4280 69604
rect 4296 69660 4360 69664
rect 4296 69604 4300 69660
rect 4300 69604 4356 69660
rect 4356 69604 4360 69660
rect 4296 69600 4360 69604
rect 4376 69660 4440 69664
rect 4376 69604 4380 69660
rect 4380 69604 4436 69660
rect 4436 69604 4440 69660
rect 4376 69600 4440 69604
rect 4456 69660 4520 69664
rect 4456 69604 4460 69660
rect 4460 69604 4516 69660
rect 4516 69604 4520 69660
rect 4456 69600 4520 69604
rect 7480 69660 7544 69664
rect 7480 69604 7484 69660
rect 7484 69604 7540 69660
rect 7540 69604 7544 69660
rect 7480 69600 7544 69604
rect 7560 69660 7624 69664
rect 7560 69604 7564 69660
rect 7564 69604 7620 69660
rect 7620 69604 7624 69660
rect 7560 69600 7624 69604
rect 7640 69660 7704 69664
rect 7640 69604 7644 69660
rect 7644 69604 7700 69660
rect 7700 69604 7704 69660
rect 7640 69600 7704 69604
rect 7720 69660 7784 69664
rect 7720 69604 7724 69660
rect 7724 69604 7780 69660
rect 7780 69604 7784 69660
rect 7720 69600 7784 69604
rect 2268 69260 2332 69324
rect 2584 69116 2648 69120
rect 2584 69060 2588 69116
rect 2588 69060 2644 69116
rect 2644 69060 2648 69116
rect 2584 69056 2648 69060
rect 2664 69116 2728 69120
rect 2664 69060 2668 69116
rect 2668 69060 2724 69116
rect 2724 69060 2728 69116
rect 2664 69056 2728 69060
rect 2744 69116 2808 69120
rect 2744 69060 2748 69116
rect 2748 69060 2804 69116
rect 2804 69060 2808 69116
rect 2744 69056 2808 69060
rect 2824 69116 2888 69120
rect 2824 69060 2828 69116
rect 2828 69060 2884 69116
rect 2884 69060 2888 69116
rect 2824 69056 2888 69060
rect 5848 69116 5912 69120
rect 5848 69060 5852 69116
rect 5852 69060 5908 69116
rect 5908 69060 5912 69116
rect 5848 69056 5912 69060
rect 5928 69116 5992 69120
rect 5928 69060 5932 69116
rect 5932 69060 5988 69116
rect 5988 69060 5992 69116
rect 5928 69056 5992 69060
rect 6008 69116 6072 69120
rect 6008 69060 6012 69116
rect 6012 69060 6068 69116
rect 6068 69060 6072 69116
rect 6008 69056 6072 69060
rect 6088 69116 6152 69120
rect 6088 69060 6092 69116
rect 6092 69060 6148 69116
rect 6148 69060 6152 69116
rect 6088 69056 6152 69060
rect 9112 69116 9176 69120
rect 9112 69060 9116 69116
rect 9116 69060 9172 69116
rect 9172 69060 9176 69116
rect 9112 69056 9176 69060
rect 9192 69116 9256 69120
rect 9192 69060 9196 69116
rect 9196 69060 9252 69116
rect 9252 69060 9256 69116
rect 9192 69056 9256 69060
rect 9272 69116 9336 69120
rect 9272 69060 9276 69116
rect 9276 69060 9332 69116
rect 9332 69060 9336 69116
rect 9272 69056 9336 69060
rect 9352 69116 9416 69120
rect 9352 69060 9356 69116
rect 9356 69060 9412 69116
rect 9412 69060 9416 69116
rect 9352 69056 9416 69060
rect 4216 68572 4280 68576
rect 4216 68516 4220 68572
rect 4220 68516 4276 68572
rect 4276 68516 4280 68572
rect 4216 68512 4280 68516
rect 4296 68572 4360 68576
rect 4296 68516 4300 68572
rect 4300 68516 4356 68572
rect 4356 68516 4360 68572
rect 4296 68512 4360 68516
rect 4376 68572 4440 68576
rect 4376 68516 4380 68572
rect 4380 68516 4436 68572
rect 4436 68516 4440 68572
rect 4376 68512 4440 68516
rect 4456 68572 4520 68576
rect 4456 68516 4460 68572
rect 4460 68516 4516 68572
rect 4516 68516 4520 68572
rect 4456 68512 4520 68516
rect 7480 68572 7544 68576
rect 7480 68516 7484 68572
rect 7484 68516 7540 68572
rect 7540 68516 7544 68572
rect 7480 68512 7544 68516
rect 7560 68572 7624 68576
rect 7560 68516 7564 68572
rect 7564 68516 7620 68572
rect 7620 68516 7624 68572
rect 7560 68512 7624 68516
rect 7640 68572 7704 68576
rect 7640 68516 7644 68572
rect 7644 68516 7700 68572
rect 7700 68516 7704 68572
rect 7640 68512 7704 68516
rect 7720 68572 7784 68576
rect 7720 68516 7724 68572
rect 7724 68516 7780 68572
rect 7780 68516 7784 68572
rect 7720 68512 7784 68516
rect 2584 68028 2648 68032
rect 2584 67972 2588 68028
rect 2588 67972 2644 68028
rect 2644 67972 2648 68028
rect 2584 67968 2648 67972
rect 2664 68028 2728 68032
rect 2664 67972 2668 68028
rect 2668 67972 2724 68028
rect 2724 67972 2728 68028
rect 2664 67968 2728 67972
rect 2744 68028 2808 68032
rect 2744 67972 2748 68028
rect 2748 67972 2804 68028
rect 2804 67972 2808 68028
rect 2744 67968 2808 67972
rect 2824 68028 2888 68032
rect 2824 67972 2828 68028
rect 2828 67972 2884 68028
rect 2884 67972 2888 68028
rect 2824 67968 2888 67972
rect 5848 68028 5912 68032
rect 5848 67972 5852 68028
rect 5852 67972 5908 68028
rect 5908 67972 5912 68028
rect 5848 67968 5912 67972
rect 5928 68028 5992 68032
rect 5928 67972 5932 68028
rect 5932 67972 5988 68028
rect 5988 67972 5992 68028
rect 5928 67968 5992 67972
rect 6008 68028 6072 68032
rect 6008 67972 6012 68028
rect 6012 67972 6068 68028
rect 6068 67972 6072 68028
rect 6008 67968 6072 67972
rect 6088 68028 6152 68032
rect 6088 67972 6092 68028
rect 6092 67972 6148 68028
rect 6148 67972 6152 68028
rect 6088 67968 6152 67972
rect 9112 68028 9176 68032
rect 9112 67972 9116 68028
rect 9116 67972 9172 68028
rect 9172 67972 9176 68028
rect 9112 67968 9176 67972
rect 9192 68028 9256 68032
rect 9192 67972 9196 68028
rect 9196 67972 9252 68028
rect 9252 67972 9256 68028
rect 9192 67968 9256 67972
rect 9272 68028 9336 68032
rect 9272 67972 9276 68028
rect 9276 67972 9332 68028
rect 9332 67972 9336 68028
rect 9272 67968 9336 67972
rect 9352 68028 9416 68032
rect 9352 67972 9356 68028
rect 9356 67972 9412 68028
rect 9412 67972 9416 68028
rect 9352 67968 9416 67972
rect 1716 67688 1780 67692
rect 1716 67632 1730 67688
rect 1730 67632 1780 67688
rect 1716 67628 1780 67632
rect 4216 67484 4280 67488
rect 4216 67428 4220 67484
rect 4220 67428 4276 67484
rect 4276 67428 4280 67484
rect 4216 67424 4280 67428
rect 4296 67484 4360 67488
rect 4296 67428 4300 67484
rect 4300 67428 4356 67484
rect 4356 67428 4360 67484
rect 4296 67424 4360 67428
rect 4376 67484 4440 67488
rect 4376 67428 4380 67484
rect 4380 67428 4436 67484
rect 4436 67428 4440 67484
rect 4376 67424 4440 67428
rect 4456 67484 4520 67488
rect 4456 67428 4460 67484
rect 4460 67428 4516 67484
rect 4516 67428 4520 67484
rect 4456 67424 4520 67428
rect 7480 67484 7544 67488
rect 7480 67428 7484 67484
rect 7484 67428 7540 67484
rect 7540 67428 7544 67484
rect 7480 67424 7544 67428
rect 7560 67484 7624 67488
rect 7560 67428 7564 67484
rect 7564 67428 7620 67484
rect 7620 67428 7624 67484
rect 7560 67424 7624 67428
rect 7640 67484 7704 67488
rect 7640 67428 7644 67484
rect 7644 67428 7700 67484
rect 7700 67428 7704 67484
rect 7640 67424 7704 67428
rect 7720 67484 7784 67488
rect 7720 67428 7724 67484
rect 7724 67428 7780 67484
rect 7780 67428 7784 67484
rect 7720 67424 7784 67428
rect 2084 67356 2148 67420
rect 2584 66940 2648 66944
rect 2584 66884 2588 66940
rect 2588 66884 2644 66940
rect 2644 66884 2648 66940
rect 2584 66880 2648 66884
rect 2664 66940 2728 66944
rect 2664 66884 2668 66940
rect 2668 66884 2724 66940
rect 2724 66884 2728 66940
rect 2664 66880 2728 66884
rect 2744 66940 2808 66944
rect 2744 66884 2748 66940
rect 2748 66884 2804 66940
rect 2804 66884 2808 66940
rect 2744 66880 2808 66884
rect 2824 66940 2888 66944
rect 2824 66884 2828 66940
rect 2828 66884 2884 66940
rect 2884 66884 2888 66940
rect 2824 66880 2888 66884
rect 5848 66940 5912 66944
rect 5848 66884 5852 66940
rect 5852 66884 5908 66940
rect 5908 66884 5912 66940
rect 5848 66880 5912 66884
rect 5928 66940 5992 66944
rect 5928 66884 5932 66940
rect 5932 66884 5988 66940
rect 5988 66884 5992 66940
rect 5928 66880 5992 66884
rect 6008 66940 6072 66944
rect 6008 66884 6012 66940
rect 6012 66884 6068 66940
rect 6068 66884 6072 66940
rect 6008 66880 6072 66884
rect 6088 66940 6152 66944
rect 6088 66884 6092 66940
rect 6092 66884 6148 66940
rect 6148 66884 6152 66940
rect 6088 66880 6152 66884
rect 9112 66940 9176 66944
rect 9112 66884 9116 66940
rect 9116 66884 9172 66940
rect 9172 66884 9176 66940
rect 9112 66880 9176 66884
rect 9192 66940 9256 66944
rect 9192 66884 9196 66940
rect 9196 66884 9252 66940
rect 9252 66884 9256 66940
rect 9192 66880 9256 66884
rect 9272 66940 9336 66944
rect 9272 66884 9276 66940
rect 9276 66884 9332 66940
rect 9332 66884 9336 66940
rect 9272 66880 9336 66884
rect 9352 66940 9416 66944
rect 9352 66884 9356 66940
rect 9356 66884 9412 66940
rect 9412 66884 9416 66940
rect 9352 66880 9416 66884
rect 4216 66396 4280 66400
rect 4216 66340 4220 66396
rect 4220 66340 4276 66396
rect 4276 66340 4280 66396
rect 4216 66336 4280 66340
rect 4296 66396 4360 66400
rect 4296 66340 4300 66396
rect 4300 66340 4356 66396
rect 4356 66340 4360 66396
rect 4296 66336 4360 66340
rect 4376 66396 4440 66400
rect 4376 66340 4380 66396
rect 4380 66340 4436 66396
rect 4436 66340 4440 66396
rect 4376 66336 4440 66340
rect 4456 66396 4520 66400
rect 4456 66340 4460 66396
rect 4460 66340 4516 66396
rect 4516 66340 4520 66396
rect 4456 66336 4520 66340
rect 7480 66396 7544 66400
rect 7480 66340 7484 66396
rect 7484 66340 7540 66396
rect 7540 66340 7544 66396
rect 7480 66336 7544 66340
rect 7560 66396 7624 66400
rect 7560 66340 7564 66396
rect 7564 66340 7620 66396
rect 7620 66340 7624 66396
rect 7560 66336 7624 66340
rect 7640 66396 7704 66400
rect 7640 66340 7644 66396
rect 7644 66340 7700 66396
rect 7700 66340 7704 66396
rect 7640 66336 7704 66340
rect 7720 66396 7784 66400
rect 7720 66340 7724 66396
rect 7724 66340 7780 66396
rect 7780 66340 7784 66396
rect 7720 66336 7784 66340
rect 2584 65852 2648 65856
rect 2584 65796 2588 65852
rect 2588 65796 2644 65852
rect 2644 65796 2648 65852
rect 2584 65792 2648 65796
rect 2664 65852 2728 65856
rect 2664 65796 2668 65852
rect 2668 65796 2724 65852
rect 2724 65796 2728 65852
rect 2664 65792 2728 65796
rect 2744 65852 2808 65856
rect 2744 65796 2748 65852
rect 2748 65796 2804 65852
rect 2804 65796 2808 65852
rect 2744 65792 2808 65796
rect 2824 65852 2888 65856
rect 2824 65796 2828 65852
rect 2828 65796 2884 65852
rect 2884 65796 2888 65852
rect 2824 65792 2888 65796
rect 5848 65852 5912 65856
rect 5848 65796 5852 65852
rect 5852 65796 5908 65852
rect 5908 65796 5912 65852
rect 5848 65792 5912 65796
rect 5928 65852 5992 65856
rect 5928 65796 5932 65852
rect 5932 65796 5988 65852
rect 5988 65796 5992 65852
rect 5928 65792 5992 65796
rect 6008 65852 6072 65856
rect 6008 65796 6012 65852
rect 6012 65796 6068 65852
rect 6068 65796 6072 65852
rect 6008 65792 6072 65796
rect 6088 65852 6152 65856
rect 6088 65796 6092 65852
rect 6092 65796 6148 65852
rect 6148 65796 6152 65852
rect 6088 65792 6152 65796
rect 9112 65852 9176 65856
rect 9112 65796 9116 65852
rect 9116 65796 9172 65852
rect 9172 65796 9176 65852
rect 9112 65792 9176 65796
rect 9192 65852 9256 65856
rect 9192 65796 9196 65852
rect 9196 65796 9252 65852
rect 9252 65796 9256 65852
rect 9192 65792 9256 65796
rect 9272 65852 9336 65856
rect 9272 65796 9276 65852
rect 9276 65796 9332 65852
rect 9332 65796 9336 65852
rect 9272 65792 9336 65796
rect 9352 65852 9416 65856
rect 9352 65796 9356 65852
rect 9356 65796 9412 65852
rect 9412 65796 9416 65852
rect 9352 65792 9416 65796
rect 4216 65308 4280 65312
rect 4216 65252 4220 65308
rect 4220 65252 4276 65308
rect 4276 65252 4280 65308
rect 4216 65248 4280 65252
rect 4296 65308 4360 65312
rect 4296 65252 4300 65308
rect 4300 65252 4356 65308
rect 4356 65252 4360 65308
rect 4296 65248 4360 65252
rect 4376 65308 4440 65312
rect 4376 65252 4380 65308
rect 4380 65252 4436 65308
rect 4436 65252 4440 65308
rect 4376 65248 4440 65252
rect 4456 65308 4520 65312
rect 4456 65252 4460 65308
rect 4460 65252 4516 65308
rect 4516 65252 4520 65308
rect 4456 65248 4520 65252
rect 7480 65308 7544 65312
rect 7480 65252 7484 65308
rect 7484 65252 7540 65308
rect 7540 65252 7544 65308
rect 7480 65248 7544 65252
rect 7560 65308 7624 65312
rect 7560 65252 7564 65308
rect 7564 65252 7620 65308
rect 7620 65252 7624 65308
rect 7560 65248 7624 65252
rect 7640 65308 7704 65312
rect 7640 65252 7644 65308
rect 7644 65252 7700 65308
rect 7700 65252 7704 65308
rect 7640 65248 7704 65252
rect 7720 65308 7784 65312
rect 7720 65252 7724 65308
rect 7724 65252 7780 65308
rect 7780 65252 7784 65308
rect 7720 65248 7784 65252
rect 1348 64908 1412 64972
rect 2584 64764 2648 64768
rect 2584 64708 2588 64764
rect 2588 64708 2644 64764
rect 2644 64708 2648 64764
rect 2584 64704 2648 64708
rect 2664 64764 2728 64768
rect 2664 64708 2668 64764
rect 2668 64708 2724 64764
rect 2724 64708 2728 64764
rect 2664 64704 2728 64708
rect 2744 64764 2808 64768
rect 2744 64708 2748 64764
rect 2748 64708 2804 64764
rect 2804 64708 2808 64764
rect 2744 64704 2808 64708
rect 2824 64764 2888 64768
rect 2824 64708 2828 64764
rect 2828 64708 2884 64764
rect 2884 64708 2888 64764
rect 2824 64704 2888 64708
rect 5848 64764 5912 64768
rect 5848 64708 5852 64764
rect 5852 64708 5908 64764
rect 5908 64708 5912 64764
rect 5848 64704 5912 64708
rect 5928 64764 5992 64768
rect 5928 64708 5932 64764
rect 5932 64708 5988 64764
rect 5988 64708 5992 64764
rect 5928 64704 5992 64708
rect 6008 64764 6072 64768
rect 6008 64708 6012 64764
rect 6012 64708 6068 64764
rect 6068 64708 6072 64764
rect 6008 64704 6072 64708
rect 6088 64764 6152 64768
rect 6088 64708 6092 64764
rect 6092 64708 6148 64764
rect 6148 64708 6152 64764
rect 6088 64704 6152 64708
rect 9112 64764 9176 64768
rect 9112 64708 9116 64764
rect 9116 64708 9172 64764
rect 9172 64708 9176 64764
rect 9112 64704 9176 64708
rect 9192 64764 9256 64768
rect 9192 64708 9196 64764
rect 9196 64708 9252 64764
rect 9252 64708 9256 64764
rect 9192 64704 9256 64708
rect 9272 64764 9336 64768
rect 9272 64708 9276 64764
rect 9276 64708 9332 64764
rect 9332 64708 9336 64764
rect 9272 64704 9336 64708
rect 9352 64764 9416 64768
rect 9352 64708 9356 64764
rect 9356 64708 9412 64764
rect 9412 64708 9416 64764
rect 9352 64704 9416 64708
rect 4216 64220 4280 64224
rect 4216 64164 4220 64220
rect 4220 64164 4276 64220
rect 4276 64164 4280 64220
rect 4216 64160 4280 64164
rect 4296 64220 4360 64224
rect 4296 64164 4300 64220
rect 4300 64164 4356 64220
rect 4356 64164 4360 64220
rect 4296 64160 4360 64164
rect 4376 64220 4440 64224
rect 4376 64164 4380 64220
rect 4380 64164 4436 64220
rect 4436 64164 4440 64220
rect 4376 64160 4440 64164
rect 4456 64220 4520 64224
rect 4456 64164 4460 64220
rect 4460 64164 4516 64220
rect 4516 64164 4520 64220
rect 4456 64160 4520 64164
rect 7480 64220 7544 64224
rect 7480 64164 7484 64220
rect 7484 64164 7540 64220
rect 7540 64164 7544 64220
rect 7480 64160 7544 64164
rect 7560 64220 7624 64224
rect 7560 64164 7564 64220
rect 7564 64164 7620 64220
rect 7620 64164 7624 64220
rect 7560 64160 7624 64164
rect 7640 64220 7704 64224
rect 7640 64164 7644 64220
rect 7644 64164 7700 64220
rect 7700 64164 7704 64220
rect 7640 64160 7704 64164
rect 7720 64220 7784 64224
rect 7720 64164 7724 64220
rect 7724 64164 7780 64220
rect 7780 64164 7784 64220
rect 7720 64160 7784 64164
rect 2268 64152 2332 64156
rect 2268 64096 2282 64152
rect 2282 64096 2332 64152
rect 2268 64092 2332 64096
rect 2584 63676 2648 63680
rect 2584 63620 2588 63676
rect 2588 63620 2644 63676
rect 2644 63620 2648 63676
rect 2584 63616 2648 63620
rect 2664 63676 2728 63680
rect 2664 63620 2668 63676
rect 2668 63620 2724 63676
rect 2724 63620 2728 63676
rect 2664 63616 2728 63620
rect 2744 63676 2808 63680
rect 2744 63620 2748 63676
rect 2748 63620 2804 63676
rect 2804 63620 2808 63676
rect 2744 63616 2808 63620
rect 2824 63676 2888 63680
rect 2824 63620 2828 63676
rect 2828 63620 2884 63676
rect 2884 63620 2888 63676
rect 2824 63616 2888 63620
rect 5848 63676 5912 63680
rect 5848 63620 5852 63676
rect 5852 63620 5908 63676
rect 5908 63620 5912 63676
rect 5848 63616 5912 63620
rect 5928 63676 5992 63680
rect 5928 63620 5932 63676
rect 5932 63620 5988 63676
rect 5988 63620 5992 63676
rect 5928 63616 5992 63620
rect 6008 63676 6072 63680
rect 6008 63620 6012 63676
rect 6012 63620 6068 63676
rect 6068 63620 6072 63676
rect 6008 63616 6072 63620
rect 6088 63676 6152 63680
rect 6088 63620 6092 63676
rect 6092 63620 6148 63676
rect 6148 63620 6152 63676
rect 6088 63616 6152 63620
rect 9112 63676 9176 63680
rect 9112 63620 9116 63676
rect 9116 63620 9172 63676
rect 9172 63620 9176 63676
rect 9112 63616 9176 63620
rect 9192 63676 9256 63680
rect 9192 63620 9196 63676
rect 9196 63620 9252 63676
rect 9252 63620 9256 63676
rect 9192 63616 9256 63620
rect 9272 63676 9336 63680
rect 9272 63620 9276 63676
rect 9276 63620 9332 63676
rect 9332 63620 9336 63676
rect 9272 63616 9336 63620
rect 9352 63676 9416 63680
rect 9352 63620 9356 63676
rect 9356 63620 9412 63676
rect 9412 63620 9416 63676
rect 9352 63616 9416 63620
rect 3556 63412 3620 63476
rect 4216 63132 4280 63136
rect 4216 63076 4220 63132
rect 4220 63076 4276 63132
rect 4276 63076 4280 63132
rect 4216 63072 4280 63076
rect 4296 63132 4360 63136
rect 4296 63076 4300 63132
rect 4300 63076 4356 63132
rect 4356 63076 4360 63132
rect 4296 63072 4360 63076
rect 4376 63132 4440 63136
rect 4376 63076 4380 63132
rect 4380 63076 4436 63132
rect 4436 63076 4440 63132
rect 4376 63072 4440 63076
rect 4456 63132 4520 63136
rect 4456 63076 4460 63132
rect 4460 63076 4516 63132
rect 4516 63076 4520 63132
rect 4456 63072 4520 63076
rect 7480 63132 7544 63136
rect 7480 63076 7484 63132
rect 7484 63076 7540 63132
rect 7540 63076 7544 63132
rect 7480 63072 7544 63076
rect 7560 63132 7624 63136
rect 7560 63076 7564 63132
rect 7564 63076 7620 63132
rect 7620 63076 7624 63132
rect 7560 63072 7624 63076
rect 7640 63132 7704 63136
rect 7640 63076 7644 63132
rect 7644 63076 7700 63132
rect 7700 63076 7704 63132
rect 7640 63072 7704 63076
rect 7720 63132 7784 63136
rect 7720 63076 7724 63132
rect 7724 63076 7780 63132
rect 7780 63076 7784 63132
rect 7720 63072 7784 63076
rect 1900 62868 1964 62932
rect 2584 62588 2648 62592
rect 2584 62532 2588 62588
rect 2588 62532 2644 62588
rect 2644 62532 2648 62588
rect 2584 62528 2648 62532
rect 2664 62588 2728 62592
rect 2664 62532 2668 62588
rect 2668 62532 2724 62588
rect 2724 62532 2728 62588
rect 2664 62528 2728 62532
rect 2744 62588 2808 62592
rect 2744 62532 2748 62588
rect 2748 62532 2804 62588
rect 2804 62532 2808 62588
rect 2744 62528 2808 62532
rect 2824 62588 2888 62592
rect 2824 62532 2828 62588
rect 2828 62532 2884 62588
rect 2884 62532 2888 62588
rect 2824 62528 2888 62532
rect 5848 62588 5912 62592
rect 5848 62532 5852 62588
rect 5852 62532 5908 62588
rect 5908 62532 5912 62588
rect 5848 62528 5912 62532
rect 5928 62588 5992 62592
rect 5928 62532 5932 62588
rect 5932 62532 5988 62588
rect 5988 62532 5992 62588
rect 5928 62528 5992 62532
rect 6008 62588 6072 62592
rect 6008 62532 6012 62588
rect 6012 62532 6068 62588
rect 6068 62532 6072 62588
rect 6008 62528 6072 62532
rect 6088 62588 6152 62592
rect 6088 62532 6092 62588
rect 6092 62532 6148 62588
rect 6148 62532 6152 62588
rect 6088 62528 6152 62532
rect 9112 62588 9176 62592
rect 9112 62532 9116 62588
rect 9116 62532 9172 62588
rect 9172 62532 9176 62588
rect 9112 62528 9176 62532
rect 9192 62588 9256 62592
rect 9192 62532 9196 62588
rect 9196 62532 9252 62588
rect 9252 62532 9256 62588
rect 9192 62528 9256 62532
rect 9272 62588 9336 62592
rect 9272 62532 9276 62588
rect 9276 62532 9332 62588
rect 9332 62532 9336 62588
rect 9272 62528 9336 62532
rect 9352 62588 9416 62592
rect 9352 62532 9356 62588
rect 9356 62532 9412 62588
rect 9412 62532 9416 62588
rect 9352 62528 9416 62532
rect 1532 62188 1596 62252
rect 4216 62044 4280 62048
rect 4216 61988 4220 62044
rect 4220 61988 4276 62044
rect 4276 61988 4280 62044
rect 4216 61984 4280 61988
rect 4296 62044 4360 62048
rect 4296 61988 4300 62044
rect 4300 61988 4356 62044
rect 4356 61988 4360 62044
rect 4296 61984 4360 61988
rect 4376 62044 4440 62048
rect 4376 61988 4380 62044
rect 4380 61988 4436 62044
rect 4436 61988 4440 62044
rect 4376 61984 4440 61988
rect 4456 62044 4520 62048
rect 4456 61988 4460 62044
rect 4460 61988 4516 62044
rect 4516 61988 4520 62044
rect 4456 61984 4520 61988
rect 7480 62044 7544 62048
rect 7480 61988 7484 62044
rect 7484 61988 7540 62044
rect 7540 61988 7544 62044
rect 7480 61984 7544 61988
rect 7560 62044 7624 62048
rect 7560 61988 7564 62044
rect 7564 61988 7620 62044
rect 7620 61988 7624 62044
rect 7560 61984 7624 61988
rect 7640 62044 7704 62048
rect 7640 61988 7644 62044
rect 7644 61988 7700 62044
rect 7700 61988 7704 62044
rect 7640 61984 7704 61988
rect 7720 62044 7784 62048
rect 7720 61988 7724 62044
rect 7724 61988 7780 62044
rect 7780 61988 7784 62044
rect 7720 61984 7784 61988
rect 3372 61780 3436 61844
rect 2584 61500 2648 61504
rect 2584 61444 2588 61500
rect 2588 61444 2644 61500
rect 2644 61444 2648 61500
rect 2584 61440 2648 61444
rect 2664 61500 2728 61504
rect 2664 61444 2668 61500
rect 2668 61444 2724 61500
rect 2724 61444 2728 61500
rect 2664 61440 2728 61444
rect 2744 61500 2808 61504
rect 2744 61444 2748 61500
rect 2748 61444 2804 61500
rect 2804 61444 2808 61500
rect 2744 61440 2808 61444
rect 2824 61500 2888 61504
rect 2824 61444 2828 61500
rect 2828 61444 2884 61500
rect 2884 61444 2888 61500
rect 2824 61440 2888 61444
rect 5848 61500 5912 61504
rect 5848 61444 5852 61500
rect 5852 61444 5908 61500
rect 5908 61444 5912 61500
rect 5848 61440 5912 61444
rect 5928 61500 5992 61504
rect 5928 61444 5932 61500
rect 5932 61444 5988 61500
rect 5988 61444 5992 61500
rect 5928 61440 5992 61444
rect 6008 61500 6072 61504
rect 6008 61444 6012 61500
rect 6012 61444 6068 61500
rect 6068 61444 6072 61500
rect 6008 61440 6072 61444
rect 6088 61500 6152 61504
rect 6088 61444 6092 61500
rect 6092 61444 6148 61500
rect 6148 61444 6152 61500
rect 6088 61440 6152 61444
rect 9112 61500 9176 61504
rect 9112 61444 9116 61500
rect 9116 61444 9172 61500
rect 9172 61444 9176 61500
rect 9112 61440 9176 61444
rect 9192 61500 9256 61504
rect 9192 61444 9196 61500
rect 9196 61444 9252 61500
rect 9252 61444 9256 61500
rect 9192 61440 9256 61444
rect 9272 61500 9336 61504
rect 9272 61444 9276 61500
rect 9276 61444 9332 61500
rect 9332 61444 9336 61500
rect 9272 61440 9336 61444
rect 9352 61500 9416 61504
rect 9352 61444 9356 61500
rect 9356 61444 9412 61500
rect 9412 61444 9416 61500
rect 9352 61440 9416 61444
rect 2268 61236 2332 61300
rect 2084 61100 2148 61164
rect 2084 60964 2148 61028
rect 3188 60964 3252 61028
rect 4216 60956 4280 60960
rect 4216 60900 4220 60956
rect 4220 60900 4276 60956
rect 4276 60900 4280 60956
rect 4216 60896 4280 60900
rect 4296 60956 4360 60960
rect 4296 60900 4300 60956
rect 4300 60900 4356 60956
rect 4356 60900 4360 60956
rect 4296 60896 4360 60900
rect 4376 60956 4440 60960
rect 4376 60900 4380 60956
rect 4380 60900 4436 60956
rect 4436 60900 4440 60956
rect 4376 60896 4440 60900
rect 4456 60956 4520 60960
rect 4456 60900 4460 60956
rect 4460 60900 4516 60956
rect 4516 60900 4520 60956
rect 4456 60896 4520 60900
rect 7480 60956 7544 60960
rect 7480 60900 7484 60956
rect 7484 60900 7540 60956
rect 7540 60900 7544 60956
rect 7480 60896 7544 60900
rect 7560 60956 7624 60960
rect 7560 60900 7564 60956
rect 7564 60900 7620 60956
rect 7620 60900 7624 60956
rect 7560 60896 7624 60900
rect 7640 60956 7704 60960
rect 7640 60900 7644 60956
rect 7644 60900 7700 60956
rect 7700 60900 7704 60956
rect 7640 60896 7704 60900
rect 7720 60956 7784 60960
rect 7720 60900 7724 60956
rect 7724 60900 7780 60956
rect 7780 60900 7784 60956
rect 7720 60896 7784 60900
rect 3004 60828 3068 60892
rect 3740 60556 3804 60620
rect 3004 60420 3068 60484
rect 2584 60412 2648 60416
rect 2584 60356 2588 60412
rect 2588 60356 2644 60412
rect 2644 60356 2648 60412
rect 2584 60352 2648 60356
rect 2664 60412 2728 60416
rect 2664 60356 2668 60412
rect 2668 60356 2724 60412
rect 2724 60356 2728 60412
rect 2664 60352 2728 60356
rect 2744 60412 2808 60416
rect 2744 60356 2748 60412
rect 2748 60356 2804 60412
rect 2804 60356 2808 60412
rect 2744 60352 2808 60356
rect 2824 60412 2888 60416
rect 2824 60356 2828 60412
rect 2828 60356 2884 60412
rect 2884 60356 2888 60412
rect 2824 60352 2888 60356
rect 5848 60412 5912 60416
rect 5848 60356 5852 60412
rect 5852 60356 5908 60412
rect 5908 60356 5912 60412
rect 5848 60352 5912 60356
rect 5928 60412 5992 60416
rect 5928 60356 5932 60412
rect 5932 60356 5988 60412
rect 5988 60356 5992 60412
rect 5928 60352 5992 60356
rect 6008 60412 6072 60416
rect 6008 60356 6012 60412
rect 6012 60356 6068 60412
rect 6068 60356 6072 60412
rect 6008 60352 6072 60356
rect 6088 60412 6152 60416
rect 6088 60356 6092 60412
rect 6092 60356 6148 60412
rect 6148 60356 6152 60412
rect 6088 60352 6152 60356
rect 9112 60412 9176 60416
rect 9112 60356 9116 60412
rect 9116 60356 9172 60412
rect 9172 60356 9176 60412
rect 9112 60352 9176 60356
rect 9192 60412 9256 60416
rect 9192 60356 9196 60412
rect 9196 60356 9252 60412
rect 9252 60356 9256 60412
rect 9192 60352 9256 60356
rect 9272 60412 9336 60416
rect 9272 60356 9276 60412
rect 9276 60356 9332 60412
rect 9332 60356 9336 60412
rect 9272 60352 9336 60356
rect 9352 60412 9416 60416
rect 9352 60356 9356 60412
rect 9356 60356 9412 60412
rect 9412 60356 9416 60412
rect 9352 60352 9416 60356
rect 3372 60284 3436 60348
rect 4216 59868 4280 59872
rect 4216 59812 4220 59868
rect 4220 59812 4276 59868
rect 4276 59812 4280 59868
rect 4216 59808 4280 59812
rect 4296 59868 4360 59872
rect 4296 59812 4300 59868
rect 4300 59812 4356 59868
rect 4356 59812 4360 59868
rect 4296 59808 4360 59812
rect 4376 59868 4440 59872
rect 4376 59812 4380 59868
rect 4380 59812 4436 59868
rect 4436 59812 4440 59868
rect 4376 59808 4440 59812
rect 4456 59868 4520 59872
rect 4456 59812 4460 59868
rect 4460 59812 4516 59868
rect 4516 59812 4520 59868
rect 4456 59808 4520 59812
rect 7480 59868 7544 59872
rect 7480 59812 7484 59868
rect 7484 59812 7540 59868
rect 7540 59812 7544 59868
rect 7480 59808 7544 59812
rect 7560 59868 7624 59872
rect 7560 59812 7564 59868
rect 7564 59812 7620 59868
rect 7620 59812 7624 59868
rect 7560 59808 7624 59812
rect 7640 59868 7704 59872
rect 7640 59812 7644 59868
rect 7644 59812 7700 59868
rect 7700 59812 7704 59868
rect 7640 59808 7704 59812
rect 7720 59868 7784 59872
rect 7720 59812 7724 59868
rect 7724 59812 7780 59868
rect 7780 59812 7784 59868
rect 7720 59808 7784 59812
rect 2268 59468 2332 59532
rect 2584 59324 2648 59328
rect 2584 59268 2588 59324
rect 2588 59268 2644 59324
rect 2644 59268 2648 59324
rect 2584 59264 2648 59268
rect 2664 59324 2728 59328
rect 2664 59268 2668 59324
rect 2668 59268 2724 59324
rect 2724 59268 2728 59324
rect 2664 59264 2728 59268
rect 2744 59324 2808 59328
rect 2744 59268 2748 59324
rect 2748 59268 2804 59324
rect 2804 59268 2808 59324
rect 2744 59264 2808 59268
rect 2824 59324 2888 59328
rect 2824 59268 2828 59324
rect 2828 59268 2884 59324
rect 2884 59268 2888 59324
rect 2824 59264 2888 59268
rect 5848 59324 5912 59328
rect 5848 59268 5852 59324
rect 5852 59268 5908 59324
rect 5908 59268 5912 59324
rect 5848 59264 5912 59268
rect 5928 59324 5992 59328
rect 5928 59268 5932 59324
rect 5932 59268 5988 59324
rect 5988 59268 5992 59324
rect 5928 59264 5992 59268
rect 6008 59324 6072 59328
rect 6008 59268 6012 59324
rect 6012 59268 6068 59324
rect 6068 59268 6072 59324
rect 6008 59264 6072 59268
rect 6088 59324 6152 59328
rect 6088 59268 6092 59324
rect 6092 59268 6148 59324
rect 6148 59268 6152 59324
rect 6088 59264 6152 59268
rect 9112 59324 9176 59328
rect 9112 59268 9116 59324
rect 9116 59268 9172 59324
rect 9172 59268 9176 59324
rect 9112 59264 9176 59268
rect 9192 59324 9256 59328
rect 9192 59268 9196 59324
rect 9196 59268 9252 59324
rect 9252 59268 9256 59324
rect 9192 59264 9256 59268
rect 9272 59324 9336 59328
rect 9272 59268 9276 59324
rect 9276 59268 9332 59324
rect 9332 59268 9336 59324
rect 9272 59264 9336 59268
rect 9352 59324 9416 59328
rect 9352 59268 9356 59324
rect 9356 59268 9412 59324
rect 9412 59268 9416 59324
rect 9352 59264 9416 59268
rect 4216 58780 4280 58784
rect 4216 58724 4220 58780
rect 4220 58724 4276 58780
rect 4276 58724 4280 58780
rect 4216 58720 4280 58724
rect 4296 58780 4360 58784
rect 4296 58724 4300 58780
rect 4300 58724 4356 58780
rect 4356 58724 4360 58780
rect 4296 58720 4360 58724
rect 4376 58780 4440 58784
rect 4376 58724 4380 58780
rect 4380 58724 4436 58780
rect 4436 58724 4440 58780
rect 4376 58720 4440 58724
rect 4456 58780 4520 58784
rect 4456 58724 4460 58780
rect 4460 58724 4516 58780
rect 4516 58724 4520 58780
rect 4456 58720 4520 58724
rect 7480 58780 7544 58784
rect 7480 58724 7484 58780
rect 7484 58724 7540 58780
rect 7540 58724 7544 58780
rect 7480 58720 7544 58724
rect 7560 58780 7624 58784
rect 7560 58724 7564 58780
rect 7564 58724 7620 58780
rect 7620 58724 7624 58780
rect 7560 58720 7624 58724
rect 7640 58780 7704 58784
rect 7640 58724 7644 58780
rect 7644 58724 7700 58780
rect 7700 58724 7704 58780
rect 7640 58720 7704 58724
rect 7720 58780 7784 58784
rect 7720 58724 7724 58780
rect 7724 58724 7780 58780
rect 7780 58724 7784 58780
rect 7720 58720 7784 58724
rect 3556 58516 3620 58580
rect 2584 58236 2648 58240
rect 2584 58180 2588 58236
rect 2588 58180 2644 58236
rect 2644 58180 2648 58236
rect 2584 58176 2648 58180
rect 2664 58236 2728 58240
rect 2664 58180 2668 58236
rect 2668 58180 2724 58236
rect 2724 58180 2728 58236
rect 2664 58176 2728 58180
rect 2744 58236 2808 58240
rect 2744 58180 2748 58236
rect 2748 58180 2804 58236
rect 2804 58180 2808 58236
rect 2744 58176 2808 58180
rect 2824 58236 2888 58240
rect 2824 58180 2828 58236
rect 2828 58180 2884 58236
rect 2884 58180 2888 58236
rect 2824 58176 2888 58180
rect 5848 58236 5912 58240
rect 5848 58180 5852 58236
rect 5852 58180 5908 58236
rect 5908 58180 5912 58236
rect 5848 58176 5912 58180
rect 5928 58236 5992 58240
rect 5928 58180 5932 58236
rect 5932 58180 5988 58236
rect 5988 58180 5992 58236
rect 5928 58176 5992 58180
rect 6008 58236 6072 58240
rect 6008 58180 6012 58236
rect 6012 58180 6068 58236
rect 6068 58180 6072 58236
rect 6008 58176 6072 58180
rect 6088 58236 6152 58240
rect 6088 58180 6092 58236
rect 6092 58180 6148 58236
rect 6148 58180 6152 58236
rect 6088 58176 6152 58180
rect 9112 58236 9176 58240
rect 9112 58180 9116 58236
rect 9116 58180 9172 58236
rect 9172 58180 9176 58236
rect 9112 58176 9176 58180
rect 9192 58236 9256 58240
rect 9192 58180 9196 58236
rect 9196 58180 9252 58236
rect 9252 58180 9256 58236
rect 9192 58176 9256 58180
rect 9272 58236 9336 58240
rect 9272 58180 9276 58236
rect 9276 58180 9332 58236
rect 9332 58180 9336 58236
rect 9272 58176 9336 58180
rect 9352 58236 9416 58240
rect 9352 58180 9356 58236
rect 9356 58180 9412 58236
rect 9412 58180 9416 58236
rect 9352 58176 9416 58180
rect 4216 57692 4280 57696
rect 4216 57636 4220 57692
rect 4220 57636 4276 57692
rect 4276 57636 4280 57692
rect 4216 57632 4280 57636
rect 4296 57692 4360 57696
rect 4296 57636 4300 57692
rect 4300 57636 4356 57692
rect 4356 57636 4360 57692
rect 4296 57632 4360 57636
rect 4376 57692 4440 57696
rect 4376 57636 4380 57692
rect 4380 57636 4436 57692
rect 4436 57636 4440 57692
rect 4376 57632 4440 57636
rect 4456 57692 4520 57696
rect 4456 57636 4460 57692
rect 4460 57636 4516 57692
rect 4516 57636 4520 57692
rect 4456 57632 4520 57636
rect 7480 57692 7544 57696
rect 7480 57636 7484 57692
rect 7484 57636 7540 57692
rect 7540 57636 7544 57692
rect 7480 57632 7544 57636
rect 7560 57692 7624 57696
rect 7560 57636 7564 57692
rect 7564 57636 7620 57692
rect 7620 57636 7624 57692
rect 7560 57632 7624 57636
rect 7640 57692 7704 57696
rect 7640 57636 7644 57692
rect 7644 57636 7700 57692
rect 7700 57636 7704 57692
rect 7640 57632 7704 57636
rect 7720 57692 7784 57696
rect 7720 57636 7724 57692
rect 7724 57636 7780 57692
rect 7780 57636 7784 57692
rect 7720 57632 7784 57636
rect 2268 57564 2332 57628
rect 5580 57428 5644 57492
rect 2268 57292 2332 57356
rect 2584 57148 2648 57152
rect 2584 57092 2588 57148
rect 2588 57092 2644 57148
rect 2644 57092 2648 57148
rect 2584 57088 2648 57092
rect 2664 57148 2728 57152
rect 2664 57092 2668 57148
rect 2668 57092 2724 57148
rect 2724 57092 2728 57148
rect 2664 57088 2728 57092
rect 2744 57148 2808 57152
rect 2744 57092 2748 57148
rect 2748 57092 2804 57148
rect 2804 57092 2808 57148
rect 2744 57088 2808 57092
rect 2824 57148 2888 57152
rect 2824 57092 2828 57148
rect 2828 57092 2884 57148
rect 2884 57092 2888 57148
rect 2824 57088 2888 57092
rect 5848 57148 5912 57152
rect 5848 57092 5852 57148
rect 5852 57092 5908 57148
rect 5908 57092 5912 57148
rect 5848 57088 5912 57092
rect 5928 57148 5992 57152
rect 5928 57092 5932 57148
rect 5932 57092 5988 57148
rect 5988 57092 5992 57148
rect 5928 57088 5992 57092
rect 6008 57148 6072 57152
rect 6008 57092 6012 57148
rect 6012 57092 6068 57148
rect 6068 57092 6072 57148
rect 6008 57088 6072 57092
rect 6088 57148 6152 57152
rect 6088 57092 6092 57148
rect 6092 57092 6148 57148
rect 6148 57092 6152 57148
rect 6088 57088 6152 57092
rect 9112 57148 9176 57152
rect 9112 57092 9116 57148
rect 9116 57092 9172 57148
rect 9172 57092 9176 57148
rect 9112 57088 9176 57092
rect 9192 57148 9256 57152
rect 9192 57092 9196 57148
rect 9196 57092 9252 57148
rect 9252 57092 9256 57148
rect 9192 57088 9256 57092
rect 9272 57148 9336 57152
rect 9272 57092 9276 57148
rect 9276 57092 9332 57148
rect 9332 57092 9336 57148
rect 9272 57088 9336 57092
rect 9352 57148 9416 57152
rect 9352 57092 9356 57148
rect 9356 57092 9412 57148
rect 9412 57092 9416 57148
rect 9352 57088 9416 57092
rect 4216 56604 4280 56608
rect 4216 56548 4220 56604
rect 4220 56548 4276 56604
rect 4276 56548 4280 56604
rect 4216 56544 4280 56548
rect 4296 56604 4360 56608
rect 4296 56548 4300 56604
rect 4300 56548 4356 56604
rect 4356 56548 4360 56604
rect 4296 56544 4360 56548
rect 4376 56604 4440 56608
rect 4376 56548 4380 56604
rect 4380 56548 4436 56604
rect 4436 56548 4440 56604
rect 4376 56544 4440 56548
rect 4456 56604 4520 56608
rect 4456 56548 4460 56604
rect 4460 56548 4516 56604
rect 4516 56548 4520 56604
rect 4456 56544 4520 56548
rect 7480 56604 7544 56608
rect 7480 56548 7484 56604
rect 7484 56548 7540 56604
rect 7540 56548 7544 56604
rect 7480 56544 7544 56548
rect 7560 56604 7624 56608
rect 7560 56548 7564 56604
rect 7564 56548 7620 56604
rect 7620 56548 7624 56604
rect 7560 56544 7624 56548
rect 7640 56604 7704 56608
rect 7640 56548 7644 56604
rect 7644 56548 7700 56604
rect 7700 56548 7704 56604
rect 7640 56544 7704 56548
rect 7720 56604 7784 56608
rect 7720 56548 7724 56604
rect 7724 56548 7780 56604
rect 7780 56548 7784 56604
rect 7720 56544 7784 56548
rect 60 56340 124 56404
rect 2584 56060 2648 56064
rect 2584 56004 2588 56060
rect 2588 56004 2644 56060
rect 2644 56004 2648 56060
rect 2584 56000 2648 56004
rect 2664 56060 2728 56064
rect 2664 56004 2668 56060
rect 2668 56004 2724 56060
rect 2724 56004 2728 56060
rect 2664 56000 2728 56004
rect 2744 56060 2808 56064
rect 2744 56004 2748 56060
rect 2748 56004 2804 56060
rect 2804 56004 2808 56060
rect 2744 56000 2808 56004
rect 2824 56060 2888 56064
rect 2824 56004 2828 56060
rect 2828 56004 2884 56060
rect 2884 56004 2888 56060
rect 2824 56000 2888 56004
rect 5848 56060 5912 56064
rect 5848 56004 5852 56060
rect 5852 56004 5908 56060
rect 5908 56004 5912 56060
rect 5848 56000 5912 56004
rect 5928 56060 5992 56064
rect 5928 56004 5932 56060
rect 5932 56004 5988 56060
rect 5988 56004 5992 56060
rect 5928 56000 5992 56004
rect 6008 56060 6072 56064
rect 6008 56004 6012 56060
rect 6012 56004 6068 56060
rect 6068 56004 6072 56060
rect 6008 56000 6072 56004
rect 6088 56060 6152 56064
rect 6088 56004 6092 56060
rect 6092 56004 6148 56060
rect 6148 56004 6152 56060
rect 6088 56000 6152 56004
rect 9112 56060 9176 56064
rect 9112 56004 9116 56060
rect 9116 56004 9172 56060
rect 9172 56004 9176 56060
rect 9112 56000 9176 56004
rect 9192 56060 9256 56064
rect 9192 56004 9196 56060
rect 9196 56004 9252 56060
rect 9252 56004 9256 56060
rect 9192 56000 9256 56004
rect 9272 56060 9336 56064
rect 9272 56004 9276 56060
rect 9276 56004 9332 56060
rect 9332 56004 9336 56060
rect 9272 56000 9336 56004
rect 9352 56060 9416 56064
rect 9352 56004 9356 56060
rect 9356 56004 9412 56060
rect 9412 56004 9416 56060
rect 9352 56000 9416 56004
rect 3372 55660 3436 55724
rect 4660 55660 4724 55724
rect 4216 55516 4280 55520
rect 4216 55460 4220 55516
rect 4220 55460 4276 55516
rect 4276 55460 4280 55516
rect 4216 55456 4280 55460
rect 4296 55516 4360 55520
rect 4296 55460 4300 55516
rect 4300 55460 4356 55516
rect 4356 55460 4360 55516
rect 4296 55456 4360 55460
rect 4376 55516 4440 55520
rect 4376 55460 4380 55516
rect 4380 55460 4436 55516
rect 4436 55460 4440 55516
rect 4376 55456 4440 55460
rect 4456 55516 4520 55520
rect 4456 55460 4460 55516
rect 4460 55460 4516 55516
rect 4516 55460 4520 55516
rect 4456 55456 4520 55460
rect 7480 55516 7544 55520
rect 7480 55460 7484 55516
rect 7484 55460 7540 55516
rect 7540 55460 7544 55516
rect 7480 55456 7544 55460
rect 7560 55516 7624 55520
rect 7560 55460 7564 55516
rect 7564 55460 7620 55516
rect 7620 55460 7624 55516
rect 7560 55456 7624 55460
rect 7640 55516 7704 55520
rect 7640 55460 7644 55516
rect 7644 55460 7700 55516
rect 7700 55460 7704 55516
rect 7640 55456 7704 55460
rect 7720 55516 7784 55520
rect 7720 55460 7724 55516
rect 7724 55460 7780 55516
rect 7780 55460 7784 55516
rect 7720 55456 7784 55460
rect 1164 55388 1228 55452
rect 980 55116 1044 55180
rect 2084 55116 2148 55180
rect 3004 55116 3068 55180
rect 4660 55116 4724 55180
rect 2584 54972 2648 54976
rect 2584 54916 2588 54972
rect 2588 54916 2644 54972
rect 2644 54916 2648 54972
rect 2584 54912 2648 54916
rect 2664 54972 2728 54976
rect 2664 54916 2668 54972
rect 2668 54916 2724 54972
rect 2724 54916 2728 54972
rect 2664 54912 2728 54916
rect 2744 54972 2808 54976
rect 2744 54916 2748 54972
rect 2748 54916 2804 54972
rect 2804 54916 2808 54972
rect 2744 54912 2808 54916
rect 2824 54972 2888 54976
rect 2824 54916 2828 54972
rect 2828 54916 2884 54972
rect 2884 54916 2888 54972
rect 2824 54912 2888 54916
rect 1164 54844 1228 54908
rect 980 54708 1044 54772
rect 5848 54972 5912 54976
rect 5848 54916 5852 54972
rect 5852 54916 5908 54972
rect 5908 54916 5912 54972
rect 5848 54912 5912 54916
rect 5928 54972 5992 54976
rect 5928 54916 5932 54972
rect 5932 54916 5988 54972
rect 5988 54916 5992 54972
rect 5928 54912 5992 54916
rect 6008 54972 6072 54976
rect 6008 54916 6012 54972
rect 6012 54916 6068 54972
rect 6068 54916 6072 54972
rect 6008 54912 6072 54916
rect 6088 54972 6152 54976
rect 6088 54916 6092 54972
rect 6092 54916 6148 54972
rect 6148 54916 6152 54972
rect 6088 54912 6152 54916
rect 9112 54972 9176 54976
rect 9112 54916 9116 54972
rect 9116 54916 9172 54972
rect 9172 54916 9176 54972
rect 9112 54912 9176 54916
rect 9192 54972 9256 54976
rect 9192 54916 9196 54972
rect 9196 54916 9252 54972
rect 9252 54916 9256 54972
rect 9192 54912 9256 54916
rect 9272 54972 9336 54976
rect 9272 54916 9276 54972
rect 9276 54916 9332 54972
rect 9332 54916 9336 54972
rect 9272 54912 9336 54916
rect 9352 54972 9416 54976
rect 9352 54916 9356 54972
rect 9356 54916 9412 54972
rect 9412 54916 9416 54972
rect 9352 54912 9416 54916
rect 4216 54428 4280 54432
rect 4216 54372 4220 54428
rect 4220 54372 4276 54428
rect 4276 54372 4280 54428
rect 4216 54368 4280 54372
rect 4296 54428 4360 54432
rect 4296 54372 4300 54428
rect 4300 54372 4356 54428
rect 4356 54372 4360 54428
rect 4296 54368 4360 54372
rect 4376 54428 4440 54432
rect 4376 54372 4380 54428
rect 4380 54372 4436 54428
rect 4436 54372 4440 54428
rect 4376 54368 4440 54372
rect 4456 54428 4520 54432
rect 4456 54372 4460 54428
rect 4460 54372 4516 54428
rect 4516 54372 4520 54428
rect 4456 54368 4520 54372
rect 7480 54428 7544 54432
rect 7480 54372 7484 54428
rect 7484 54372 7540 54428
rect 7540 54372 7544 54428
rect 7480 54368 7544 54372
rect 7560 54428 7624 54432
rect 7560 54372 7564 54428
rect 7564 54372 7620 54428
rect 7620 54372 7624 54428
rect 7560 54368 7624 54372
rect 7640 54428 7704 54432
rect 7640 54372 7644 54428
rect 7644 54372 7700 54428
rect 7700 54372 7704 54428
rect 7640 54368 7704 54372
rect 7720 54428 7784 54432
rect 7720 54372 7724 54428
rect 7724 54372 7780 54428
rect 7780 54372 7784 54428
rect 7720 54368 7784 54372
rect 2084 54300 2148 54364
rect 2584 53884 2648 53888
rect 2584 53828 2588 53884
rect 2588 53828 2644 53884
rect 2644 53828 2648 53884
rect 2584 53824 2648 53828
rect 2664 53884 2728 53888
rect 2664 53828 2668 53884
rect 2668 53828 2724 53884
rect 2724 53828 2728 53884
rect 2664 53824 2728 53828
rect 2744 53884 2808 53888
rect 2744 53828 2748 53884
rect 2748 53828 2804 53884
rect 2804 53828 2808 53884
rect 2744 53824 2808 53828
rect 2824 53884 2888 53888
rect 2824 53828 2828 53884
rect 2828 53828 2884 53884
rect 2884 53828 2888 53884
rect 2824 53824 2888 53828
rect 5848 53884 5912 53888
rect 5848 53828 5852 53884
rect 5852 53828 5908 53884
rect 5908 53828 5912 53884
rect 5848 53824 5912 53828
rect 5928 53884 5992 53888
rect 5928 53828 5932 53884
rect 5932 53828 5988 53884
rect 5988 53828 5992 53884
rect 5928 53824 5992 53828
rect 6008 53884 6072 53888
rect 6008 53828 6012 53884
rect 6012 53828 6068 53884
rect 6068 53828 6072 53884
rect 6008 53824 6072 53828
rect 6088 53884 6152 53888
rect 6088 53828 6092 53884
rect 6092 53828 6148 53884
rect 6148 53828 6152 53884
rect 6088 53824 6152 53828
rect 9112 53884 9176 53888
rect 9112 53828 9116 53884
rect 9116 53828 9172 53884
rect 9172 53828 9176 53884
rect 9112 53824 9176 53828
rect 9192 53884 9256 53888
rect 9192 53828 9196 53884
rect 9196 53828 9252 53884
rect 9252 53828 9256 53884
rect 9192 53824 9256 53828
rect 9272 53884 9336 53888
rect 9272 53828 9276 53884
rect 9276 53828 9332 53884
rect 9332 53828 9336 53884
rect 9272 53824 9336 53828
rect 9352 53884 9416 53888
rect 9352 53828 9356 53884
rect 9356 53828 9412 53884
rect 9412 53828 9416 53884
rect 9352 53824 9416 53828
rect 3188 53484 3252 53548
rect 4844 53484 4908 53548
rect 3188 53348 3252 53412
rect 4216 53340 4280 53344
rect 4216 53284 4220 53340
rect 4220 53284 4276 53340
rect 4276 53284 4280 53340
rect 4216 53280 4280 53284
rect 4296 53340 4360 53344
rect 4296 53284 4300 53340
rect 4300 53284 4356 53340
rect 4356 53284 4360 53340
rect 4296 53280 4360 53284
rect 4376 53340 4440 53344
rect 4376 53284 4380 53340
rect 4380 53284 4436 53340
rect 4436 53284 4440 53340
rect 4376 53280 4440 53284
rect 4456 53340 4520 53344
rect 4456 53284 4460 53340
rect 4460 53284 4516 53340
rect 4516 53284 4520 53340
rect 4456 53280 4520 53284
rect 7480 53340 7544 53344
rect 7480 53284 7484 53340
rect 7484 53284 7540 53340
rect 7540 53284 7544 53340
rect 7480 53280 7544 53284
rect 7560 53340 7624 53344
rect 7560 53284 7564 53340
rect 7564 53284 7620 53340
rect 7620 53284 7624 53340
rect 7560 53280 7624 53284
rect 7640 53340 7704 53344
rect 7640 53284 7644 53340
rect 7644 53284 7700 53340
rect 7700 53284 7704 53340
rect 7640 53280 7704 53284
rect 7720 53340 7784 53344
rect 7720 53284 7724 53340
rect 7724 53284 7780 53340
rect 7780 53284 7784 53340
rect 7720 53280 7784 53284
rect 4660 52804 4724 52868
rect 2584 52796 2648 52800
rect 2584 52740 2588 52796
rect 2588 52740 2644 52796
rect 2644 52740 2648 52796
rect 2584 52736 2648 52740
rect 2664 52796 2728 52800
rect 2664 52740 2668 52796
rect 2668 52740 2724 52796
rect 2724 52740 2728 52796
rect 2664 52736 2728 52740
rect 2744 52796 2808 52800
rect 2744 52740 2748 52796
rect 2748 52740 2804 52796
rect 2804 52740 2808 52796
rect 2744 52736 2808 52740
rect 2824 52796 2888 52800
rect 2824 52740 2828 52796
rect 2828 52740 2884 52796
rect 2884 52740 2888 52796
rect 2824 52736 2888 52740
rect 5848 52796 5912 52800
rect 5848 52740 5852 52796
rect 5852 52740 5908 52796
rect 5908 52740 5912 52796
rect 5848 52736 5912 52740
rect 5928 52796 5992 52800
rect 5928 52740 5932 52796
rect 5932 52740 5988 52796
rect 5988 52740 5992 52796
rect 5928 52736 5992 52740
rect 6008 52796 6072 52800
rect 6008 52740 6012 52796
rect 6012 52740 6068 52796
rect 6068 52740 6072 52796
rect 6008 52736 6072 52740
rect 6088 52796 6152 52800
rect 6088 52740 6092 52796
rect 6092 52740 6148 52796
rect 6148 52740 6152 52796
rect 6088 52736 6152 52740
rect 9112 52796 9176 52800
rect 9112 52740 9116 52796
rect 9116 52740 9172 52796
rect 9172 52740 9176 52796
rect 9112 52736 9176 52740
rect 9192 52796 9256 52800
rect 9192 52740 9196 52796
rect 9196 52740 9252 52796
rect 9252 52740 9256 52796
rect 9192 52736 9256 52740
rect 9272 52796 9336 52800
rect 9272 52740 9276 52796
rect 9276 52740 9332 52796
rect 9332 52740 9336 52796
rect 9272 52736 9336 52740
rect 9352 52796 9416 52800
rect 9352 52740 9356 52796
rect 9356 52740 9412 52796
rect 9412 52740 9416 52796
rect 9352 52736 9416 52740
rect 3740 52668 3804 52732
rect 5396 52728 5460 52732
rect 5396 52672 5410 52728
rect 5410 52672 5460 52728
rect 5396 52668 5460 52672
rect 4216 52252 4280 52256
rect 4216 52196 4220 52252
rect 4220 52196 4276 52252
rect 4276 52196 4280 52252
rect 4216 52192 4280 52196
rect 4296 52252 4360 52256
rect 4296 52196 4300 52252
rect 4300 52196 4356 52252
rect 4356 52196 4360 52252
rect 4296 52192 4360 52196
rect 4376 52252 4440 52256
rect 4376 52196 4380 52252
rect 4380 52196 4436 52252
rect 4436 52196 4440 52252
rect 4376 52192 4440 52196
rect 4456 52252 4520 52256
rect 4456 52196 4460 52252
rect 4460 52196 4516 52252
rect 4516 52196 4520 52252
rect 4456 52192 4520 52196
rect 7480 52252 7544 52256
rect 7480 52196 7484 52252
rect 7484 52196 7540 52252
rect 7540 52196 7544 52252
rect 7480 52192 7544 52196
rect 7560 52252 7624 52256
rect 7560 52196 7564 52252
rect 7564 52196 7620 52252
rect 7620 52196 7624 52252
rect 7560 52192 7624 52196
rect 7640 52252 7704 52256
rect 7640 52196 7644 52252
rect 7644 52196 7700 52252
rect 7700 52196 7704 52252
rect 7640 52192 7704 52196
rect 7720 52252 7784 52256
rect 7720 52196 7724 52252
rect 7724 52196 7780 52252
rect 7780 52196 7784 52252
rect 7720 52192 7784 52196
rect 5212 52124 5276 52188
rect 2584 51708 2648 51712
rect 2584 51652 2588 51708
rect 2588 51652 2644 51708
rect 2644 51652 2648 51708
rect 2584 51648 2648 51652
rect 2664 51708 2728 51712
rect 2664 51652 2668 51708
rect 2668 51652 2724 51708
rect 2724 51652 2728 51708
rect 2664 51648 2728 51652
rect 2744 51708 2808 51712
rect 2744 51652 2748 51708
rect 2748 51652 2804 51708
rect 2804 51652 2808 51708
rect 2744 51648 2808 51652
rect 2824 51708 2888 51712
rect 2824 51652 2828 51708
rect 2828 51652 2884 51708
rect 2884 51652 2888 51708
rect 2824 51648 2888 51652
rect 980 51580 1044 51644
rect 5848 51708 5912 51712
rect 5848 51652 5852 51708
rect 5852 51652 5908 51708
rect 5908 51652 5912 51708
rect 5848 51648 5912 51652
rect 5928 51708 5992 51712
rect 5928 51652 5932 51708
rect 5932 51652 5988 51708
rect 5988 51652 5992 51708
rect 5928 51648 5992 51652
rect 6008 51708 6072 51712
rect 6008 51652 6012 51708
rect 6012 51652 6068 51708
rect 6068 51652 6072 51708
rect 6008 51648 6072 51652
rect 6088 51708 6152 51712
rect 6088 51652 6092 51708
rect 6092 51652 6148 51708
rect 6148 51652 6152 51708
rect 6088 51648 6152 51652
rect 9112 51708 9176 51712
rect 9112 51652 9116 51708
rect 9116 51652 9172 51708
rect 9172 51652 9176 51708
rect 9112 51648 9176 51652
rect 9192 51708 9256 51712
rect 9192 51652 9196 51708
rect 9196 51652 9252 51708
rect 9252 51652 9256 51708
rect 9192 51648 9256 51652
rect 9272 51708 9336 51712
rect 9272 51652 9276 51708
rect 9276 51652 9332 51708
rect 9332 51652 9336 51708
rect 9272 51648 9336 51652
rect 9352 51708 9416 51712
rect 9352 51652 9356 51708
rect 9356 51652 9412 51708
rect 9412 51652 9416 51708
rect 9352 51648 9416 51652
rect 1164 51308 1228 51372
rect 2084 51308 2148 51372
rect 980 50900 1044 50964
rect 980 50764 1044 50828
rect 60 50416 124 50420
rect 60 50360 110 50416
rect 110 50360 124 50416
rect 60 50356 124 50360
rect 1716 50416 1780 50420
rect 4660 51504 4724 51508
rect 4660 51448 4674 51504
rect 4674 51448 4724 51504
rect 4660 51444 4724 51448
rect 3372 51308 3436 51372
rect 3372 51172 3436 51236
rect 4216 51164 4280 51168
rect 4216 51108 4220 51164
rect 4220 51108 4276 51164
rect 4276 51108 4280 51164
rect 4216 51104 4280 51108
rect 4296 51164 4360 51168
rect 4296 51108 4300 51164
rect 4300 51108 4356 51164
rect 4356 51108 4360 51164
rect 4296 51104 4360 51108
rect 4376 51164 4440 51168
rect 4376 51108 4380 51164
rect 4380 51108 4436 51164
rect 4436 51108 4440 51164
rect 4376 51104 4440 51108
rect 4456 51164 4520 51168
rect 4456 51108 4460 51164
rect 4460 51108 4516 51164
rect 4516 51108 4520 51164
rect 4456 51104 4520 51108
rect 7480 51164 7544 51168
rect 7480 51108 7484 51164
rect 7484 51108 7540 51164
rect 7540 51108 7544 51164
rect 7480 51104 7544 51108
rect 7560 51164 7624 51168
rect 7560 51108 7564 51164
rect 7564 51108 7620 51164
rect 7620 51108 7624 51164
rect 7560 51104 7624 51108
rect 7640 51164 7704 51168
rect 7640 51108 7644 51164
rect 7644 51108 7700 51164
rect 7700 51108 7704 51164
rect 7640 51104 7704 51108
rect 7720 51164 7784 51168
rect 7720 51108 7724 51164
rect 7724 51108 7780 51164
rect 7780 51108 7784 51164
rect 7720 51104 7784 51108
rect 5028 51028 5092 51092
rect 3372 50900 3436 50964
rect 3556 50900 3620 50964
rect 5212 50764 5276 50828
rect 4660 50628 4724 50692
rect 5396 50628 5460 50692
rect 2584 50620 2648 50624
rect 2584 50564 2588 50620
rect 2588 50564 2644 50620
rect 2644 50564 2648 50620
rect 2584 50560 2648 50564
rect 2664 50620 2728 50624
rect 2664 50564 2668 50620
rect 2668 50564 2724 50620
rect 2724 50564 2728 50620
rect 2664 50560 2728 50564
rect 2744 50620 2808 50624
rect 2744 50564 2748 50620
rect 2748 50564 2804 50620
rect 2804 50564 2808 50620
rect 2744 50560 2808 50564
rect 2824 50620 2888 50624
rect 2824 50564 2828 50620
rect 2828 50564 2884 50620
rect 2884 50564 2888 50620
rect 2824 50560 2888 50564
rect 5848 50620 5912 50624
rect 5848 50564 5852 50620
rect 5852 50564 5908 50620
rect 5908 50564 5912 50620
rect 5848 50560 5912 50564
rect 5928 50620 5992 50624
rect 5928 50564 5932 50620
rect 5932 50564 5988 50620
rect 5988 50564 5992 50620
rect 5928 50560 5992 50564
rect 6008 50620 6072 50624
rect 6008 50564 6012 50620
rect 6012 50564 6068 50620
rect 6068 50564 6072 50620
rect 6008 50560 6072 50564
rect 6088 50620 6152 50624
rect 6088 50564 6092 50620
rect 6092 50564 6148 50620
rect 6148 50564 6152 50620
rect 6088 50560 6152 50564
rect 9112 50620 9176 50624
rect 9112 50564 9116 50620
rect 9116 50564 9172 50620
rect 9172 50564 9176 50620
rect 9112 50560 9176 50564
rect 9192 50620 9256 50624
rect 9192 50564 9196 50620
rect 9196 50564 9252 50620
rect 9252 50564 9256 50620
rect 9192 50560 9256 50564
rect 9272 50620 9336 50624
rect 9272 50564 9276 50620
rect 9276 50564 9332 50620
rect 9332 50564 9336 50620
rect 9272 50560 9336 50564
rect 9352 50620 9416 50624
rect 9352 50564 9356 50620
rect 9356 50564 9412 50620
rect 9412 50564 9416 50620
rect 9352 50560 9416 50564
rect 1716 50360 1730 50416
rect 1730 50360 1780 50416
rect 1716 50356 1780 50360
rect 4660 50356 4724 50420
rect 1716 50220 1780 50284
rect 4844 50220 4908 50284
rect 3372 50084 3436 50148
rect 4216 50076 4280 50080
rect 4216 50020 4220 50076
rect 4220 50020 4276 50076
rect 4276 50020 4280 50076
rect 4216 50016 4280 50020
rect 4296 50076 4360 50080
rect 4296 50020 4300 50076
rect 4300 50020 4356 50076
rect 4356 50020 4360 50076
rect 4296 50016 4360 50020
rect 4376 50076 4440 50080
rect 4376 50020 4380 50076
rect 4380 50020 4436 50076
rect 4436 50020 4440 50076
rect 4376 50016 4440 50020
rect 4456 50076 4520 50080
rect 4456 50020 4460 50076
rect 4460 50020 4516 50076
rect 4516 50020 4520 50076
rect 4456 50016 4520 50020
rect 7480 50076 7544 50080
rect 7480 50020 7484 50076
rect 7484 50020 7540 50076
rect 7540 50020 7544 50076
rect 7480 50016 7544 50020
rect 7560 50076 7624 50080
rect 7560 50020 7564 50076
rect 7564 50020 7620 50076
rect 7620 50020 7624 50076
rect 7560 50016 7624 50020
rect 7640 50076 7704 50080
rect 7640 50020 7644 50076
rect 7644 50020 7700 50076
rect 7700 50020 7704 50076
rect 7640 50016 7704 50020
rect 7720 50076 7784 50080
rect 7720 50020 7724 50076
rect 7724 50020 7780 50076
rect 7780 50020 7784 50076
rect 7720 50016 7784 50020
rect 3740 50008 3804 50012
rect 3740 49952 3790 50008
rect 3790 49952 3804 50008
rect 3740 49948 3804 49952
rect 2584 49532 2648 49536
rect 2584 49476 2588 49532
rect 2588 49476 2644 49532
rect 2644 49476 2648 49532
rect 2584 49472 2648 49476
rect 2664 49532 2728 49536
rect 2664 49476 2668 49532
rect 2668 49476 2724 49532
rect 2724 49476 2728 49532
rect 2664 49472 2728 49476
rect 2744 49532 2808 49536
rect 2744 49476 2748 49532
rect 2748 49476 2804 49532
rect 2804 49476 2808 49532
rect 2744 49472 2808 49476
rect 2824 49532 2888 49536
rect 2824 49476 2828 49532
rect 2828 49476 2884 49532
rect 2884 49476 2888 49532
rect 2824 49472 2888 49476
rect 5848 49532 5912 49536
rect 5848 49476 5852 49532
rect 5852 49476 5908 49532
rect 5908 49476 5912 49532
rect 5848 49472 5912 49476
rect 5928 49532 5992 49536
rect 5928 49476 5932 49532
rect 5932 49476 5988 49532
rect 5988 49476 5992 49532
rect 5928 49472 5992 49476
rect 6008 49532 6072 49536
rect 6008 49476 6012 49532
rect 6012 49476 6068 49532
rect 6068 49476 6072 49532
rect 6008 49472 6072 49476
rect 6088 49532 6152 49536
rect 6088 49476 6092 49532
rect 6092 49476 6148 49532
rect 6148 49476 6152 49532
rect 6088 49472 6152 49476
rect 9112 49532 9176 49536
rect 9112 49476 9116 49532
rect 9116 49476 9172 49532
rect 9172 49476 9176 49532
rect 9112 49472 9176 49476
rect 9192 49532 9256 49536
rect 9192 49476 9196 49532
rect 9196 49476 9252 49532
rect 9252 49476 9256 49532
rect 9192 49472 9256 49476
rect 9272 49532 9336 49536
rect 9272 49476 9276 49532
rect 9276 49476 9332 49532
rect 9332 49476 9336 49532
rect 9272 49472 9336 49476
rect 9352 49532 9416 49536
rect 9352 49476 9356 49532
rect 9356 49476 9412 49532
rect 9412 49476 9416 49532
rect 9352 49472 9416 49476
rect 5212 49268 5276 49332
rect 2268 49132 2332 49196
rect 5396 49132 5460 49196
rect 4216 48988 4280 48992
rect 4216 48932 4220 48988
rect 4220 48932 4276 48988
rect 4276 48932 4280 48988
rect 4216 48928 4280 48932
rect 4296 48988 4360 48992
rect 4296 48932 4300 48988
rect 4300 48932 4356 48988
rect 4356 48932 4360 48988
rect 4296 48928 4360 48932
rect 4376 48988 4440 48992
rect 4376 48932 4380 48988
rect 4380 48932 4436 48988
rect 4436 48932 4440 48988
rect 4376 48928 4440 48932
rect 4456 48988 4520 48992
rect 4456 48932 4460 48988
rect 4460 48932 4516 48988
rect 4516 48932 4520 48988
rect 4456 48928 4520 48932
rect 7480 48988 7544 48992
rect 7480 48932 7484 48988
rect 7484 48932 7540 48988
rect 7540 48932 7544 48988
rect 7480 48928 7544 48932
rect 7560 48988 7624 48992
rect 7560 48932 7564 48988
rect 7564 48932 7620 48988
rect 7620 48932 7624 48988
rect 7560 48928 7624 48932
rect 7640 48988 7704 48992
rect 7640 48932 7644 48988
rect 7644 48932 7700 48988
rect 7700 48932 7704 48988
rect 7640 48928 7704 48932
rect 7720 48988 7784 48992
rect 7720 48932 7724 48988
rect 7724 48932 7780 48988
rect 7780 48932 7784 48988
rect 7720 48928 7784 48932
rect 2584 48444 2648 48448
rect 2584 48388 2588 48444
rect 2588 48388 2644 48444
rect 2644 48388 2648 48444
rect 2584 48384 2648 48388
rect 2664 48444 2728 48448
rect 2664 48388 2668 48444
rect 2668 48388 2724 48444
rect 2724 48388 2728 48444
rect 2664 48384 2728 48388
rect 2744 48444 2808 48448
rect 2744 48388 2748 48444
rect 2748 48388 2804 48444
rect 2804 48388 2808 48444
rect 2744 48384 2808 48388
rect 2824 48444 2888 48448
rect 2824 48388 2828 48444
rect 2828 48388 2884 48444
rect 2884 48388 2888 48444
rect 2824 48384 2888 48388
rect 1164 48376 1228 48380
rect 1164 48320 1178 48376
rect 1178 48320 1228 48376
rect 1164 48316 1228 48320
rect 1900 48180 1964 48244
rect 1900 48044 1964 48108
rect 5580 48452 5644 48516
rect 5848 48444 5912 48448
rect 5848 48388 5852 48444
rect 5852 48388 5908 48444
rect 5908 48388 5912 48444
rect 5848 48384 5912 48388
rect 5928 48444 5992 48448
rect 5928 48388 5932 48444
rect 5932 48388 5988 48444
rect 5988 48388 5992 48444
rect 5928 48384 5992 48388
rect 6008 48444 6072 48448
rect 6008 48388 6012 48444
rect 6012 48388 6068 48444
rect 6068 48388 6072 48444
rect 6008 48384 6072 48388
rect 6088 48444 6152 48448
rect 6088 48388 6092 48444
rect 6092 48388 6148 48444
rect 6148 48388 6152 48444
rect 6088 48384 6152 48388
rect 9112 48444 9176 48448
rect 9112 48388 9116 48444
rect 9116 48388 9172 48444
rect 9172 48388 9176 48444
rect 9112 48384 9176 48388
rect 9192 48444 9256 48448
rect 9192 48388 9196 48444
rect 9196 48388 9252 48444
rect 9252 48388 9256 48444
rect 9192 48384 9256 48388
rect 9272 48444 9336 48448
rect 9272 48388 9276 48444
rect 9276 48388 9332 48444
rect 9332 48388 9336 48444
rect 9272 48384 9336 48388
rect 9352 48444 9416 48448
rect 9352 48388 9356 48444
rect 9356 48388 9412 48444
rect 9412 48388 9416 48444
rect 9352 48384 9416 48388
rect 3740 48240 3804 48244
rect 3740 48184 3790 48240
rect 3790 48184 3804 48240
rect 3740 48180 3804 48184
rect 2268 47908 2332 47972
rect 4216 47900 4280 47904
rect 4216 47844 4220 47900
rect 4220 47844 4276 47900
rect 4276 47844 4280 47900
rect 4216 47840 4280 47844
rect 4296 47900 4360 47904
rect 4296 47844 4300 47900
rect 4300 47844 4356 47900
rect 4356 47844 4360 47900
rect 4296 47840 4360 47844
rect 4376 47900 4440 47904
rect 4376 47844 4380 47900
rect 4380 47844 4436 47900
rect 4436 47844 4440 47900
rect 4376 47840 4440 47844
rect 4456 47900 4520 47904
rect 4456 47844 4460 47900
rect 4460 47844 4516 47900
rect 4516 47844 4520 47900
rect 4456 47840 4520 47844
rect 7480 47900 7544 47904
rect 7480 47844 7484 47900
rect 7484 47844 7540 47900
rect 7540 47844 7544 47900
rect 7480 47840 7544 47844
rect 7560 47900 7624 47904
rect 7560 47844 7564 47900
rect 7564 47844 7620 47900
rect 7620 47844 7624 47900
rect 7560 47840 7624 47844
rect 7640 47900 7704 47904
rect 7640 47844 7644 47900
rect 7644 47844 7700 47900
rect 7700 47844 7704 47900
rect 7640 47840 7704 47844
rect 7720 47900 7784 47904
rect 7720 47844 7724 47900
rect 7724 47844 7780 47900
rect 7780 47844 7784 47900
rect 7720 47840 7784 47844
rect 2406 47772 2470 47836
rect 3740 47772 3804 47836
rect 244 47364 308 47428
rect 2584 47356 2648 47360
rect 2584 47300 2588 47356
rect 2588 47300 2644 47356
rect 2644 47300 2648 47356
rect 2584 47296 2648 47300
rect 2664 47356 2728 47360
rect 2664 47300 2668 47356
rect 2668 47300 2724 47356
rect 2724 47300 2728 47356
rect 2664 47296 2728 47300
rect 2744 47356 2808 47360
rect 2744 47300 2748 47356
rect 2748 47300 2804 47356
rect 2804 47300 2808 47356
rect 2744 47296 2808 47300
rect 2824 47356 2888 47360
rect 2824 47300 2828 47356
rect 2828 47300 2884 47356
rect 2884 47300 2888 47356
rect 2824 47296 2888 47300
rect 6316 47500 6380 47564
rect 5848 47356 5912 47360
rect 5848 47300 5852 47356
rect 5852 47300 5908 47356
rect 5908 47300 5912 47356
rect 5848 47296 5912 47300
rect 5928 47356 5992 47360
rect 5928 47300 5932 47356
rect 5932 47300 5988 47356
rect 5988 47300 5992 47356
rect 5928 47296 5992 47300
rect 6008 47356 6072 47360
rect 6008 47300 6012 47356
rect 6012 47300 6068 47356
rect 6068 47300 6072 47356
rect 6008 47296 6072 47300
rect 6088 47356 6152 47360
rect 6088 47300 6092 47356
rect 6092 47300 6148 47356
rect 6148 47300 6152 47356
rect 6088 47296 6152 47300
rect 9112 47356 9176 47360
rect 9112 47300 9116 47356
rect 9116 47300 9172 47356
rect 9172 47300 9176 47356
rect 9112 47296 9176 47300
rect 9192 47356 9256 47360
rect 9192 47300 9196 47356
rect 9196 47300 9252 47356
rect 9252 47300 9256 47356
rect 9192 47296 9256 47300
rect 9272 47356 9336 47360
rect 9272 47300 9276 47356
rect 9276 47300 9332 47356
rect 9332 47300 9336 47356
rect 9272 47296 9336 47300
rect 9352 47356 9416 47360
rect 9352 47300 9356 47356
rect 9356 47300 9412 47356
rect 9412 47300 9416 47356
rect 9352 47296 9416 47300
rect 5580 47092 5644 47156
rect 4844 46956 4908 47020
rect 1532 46820 1596 46884
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 7480 46812 7544 46816
rect 7480 46756 7484 46812
rect 7484 46756 7540 46812
rect 7540 46756 7544 46812
rect 7480 46752 7544 46756
rect 7560 46812 7624 46816
rect 7560 46756 7564 46812
rect 7564 46756 7620 46812
rect 7620 46756 7624 46812
rect 7560 46752 7624 46756
rect 7640 46812 7704 46816
rect 7640 46756 7644 46812
rect 7644 46756 7700 46812
rect 7700 46756 7704 46812
rect 7640 46752 7704 46756
rect 7720 46812 7784 46816
rect 7720 46756 7724 46812
rect 7724 46756 7780 46812
rect 7780 46756 7784 46812
rect 7720 46752 7784 46756
rect 60 46574 124 46578
rect 60 46518 110 46574
rect 110 46518 124 46574
rect 1532 46548 1596 46612
rect 8340 46548 8404 46612
rect 60 46514 124 46518
rect 5028 46412 5092 46476
rect 6500 46412 6564 46476
rect 2584 46268 2648 46272
rect 2584 46212 2588 46268
rect 2588 46212 2644 46268
rect 2644 46212 2648 46268
rect 2584 46208 2648 46212
rect 2664 46268 2728 46272
rect 2664 46212 2668 46268
rect 2668 46212 2724 46268
rect 2724 46212 2728 46268
rect 2664 46208 2728 46212
rect 2744 46268 2808 46272
rect 2744 46212 2748 46268
rect 2748 46212 2804 46268
rect 2804 46212 2808 46268
rect 2744 46208 2808 46212
rect 2824 46268 2888 46272
rect 2824 46212 2828 46268
rect 2828 46212 2884 46268
rect 2884 46212 2888 46268
rect 2824 46208 2888 46212
rect 5848 46268 5912 46272
rect 5848 46212 5852 46268
rect 5852 46212 5908 46268
rect 5908 46212 5912 46268
rect 5848 46208 5912 46212
rect 5928 46268 5992 46272
rect 5928 46212 5932 46268
rect 5932 46212 5988 46268
rect 5988 46212 5992 46268
rect 5928 46208 5992 46212
rect 6008 46268 6072 46272
rect 6008 46212 6012 46268
rect 6012 46212 6068 46268
rect 6068 46212 6072 46268
rect 6008 46208 6072 46212
rect 6088 46268 6152 46272
rect 6088 46212 6092 46268
rect 6092 46212 6148 46268
rect 6148 46212 6152 46268
rect 6088 46208 6152 46212
rect 9112 46268 9176 46272
rect 9112 46212 9116 46268
rect 9116 46212 9172 46268
rect 9172 46212 9176 46268
rect 9112 46208 9176 46212
rect 9192 46268 9256 46272
rect 9192 46212 9196 46268
rect 9196 46212 9252 46268
rect 9252 46212 9256 46268
rect 9192 46208 9256 46212
rect 9272 46268 9336 46272
rect 9272 46212 9276 46268
rect 9276 46212 9332 46268
rect 9332 46212 9336 46268
rect 9272 46208 9336 46212
rect 9352 46268 9416 46272
rect 9352 46212 9356 46268
rect 9356 46212 9412 46268
rect 9412 46212 9416 46268
rect 9352 46208 9416 46212
rect 5028 46004 5092 46068
rect 3004 45732 3068 45796
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 7480 45724 7544 45728
rect 7480 45668 7484 45724
rect 7484 45668 7540 45724
rect 7540 45668 7544 45724
rect 7480 45664 7544 45668
rect 7560 45724 7624 45728
rect 7560 45668 7564 45724
rect 7564 45668 7620 45724
rect 7620 45668 7624 45724
rect 7560 45664 7624 45668
rect 7640 45724 7704 45728
rect 7640 45668 7644 45724
rect 7644 45668 7700 45724
rect 7700 45668 7704 45724
rect 7640 45664 7704 45668
rect 7720 45724 7784 45728
rect 7720 45668 7724 45724
rect 7724 45668 7780 45724
rect 7780 45668 7784 45724
rect 7720 45664 7784 45668
rect 2406 45596 2470 45660
rect 3004 45596 3068 45660
rect 4660 45596 4724 45660
rect 1348 45324 1412 45388
rect 2406 45324 2470 45388
rect 3188 45324 3252 45388
rect 2584 45180 2648 45184
rect 2584 45124 2588 45180
rect 2588 45124 2644 45180
rect 2644 45124 2648 45180
rect 2584 45120 2648 45124
rect 2664 45180 2728 45184
rect 2664 45124 2668 45180
rect 2668 45124 2724 45180
rect 2724 45124 2728 45180
rect 2664 45120 2728 45124
rect 2744 45180 2808 45184
rect 2744 45124 2748 45180
rect 2748 45124 2804 45180
rect 2804 45124 2808 45180
rect 2744 45120 2808 45124
rect 2824 45180 2888 45184
rect 2824 45124 2828 45180
rect 2828 45124 2884 45180
rect 2884 45124 2888 45180
rect 2824 45120 2888 45124
rect 5848 45180 5912 45184
rect 5848 45124 5852 45180
rect 5852 45124 5908 45180
rect 5908 45124 5912 45180
rect 5848 45120 5912 45124
rect 5928 45180 5992 45184
rect 5928 45124 5932 45180
rect 5932 45124 5988 45180
rect 5988 45124 5992 45180
rect 5928 45120 5992 45124
rect 6008 45180 6072 45184
rect 6008 45124 6012 45180
rect 6012 45124 6068 45180
rect 6068 45124 6072 45180
rect 6008 45120 6072 45124
rect 6088 45180 6152 45184
rect 6088 45124 6092 45180
rect 6092 45124 6148 45180
rect 6148 45124 6152 45180
rect 6088 45120 6152 45124
rect 9112 45180 9176 45184
rect 9112 45124 9116 45180
rect 9116 45124 9172 45180
rect 9172 45124 9176 45180
rect 9112 45120 9176 45124
rect 9192 45180 9256 45184
rect 9192 45124 9196 45180
rect 9196 45124 9252 45180
rect 9252 45124 9256 45180
rect 9192 45120 9256 45124
rect 9272 45180 9336 45184
rect 9272 45124 9276 45180
rect 9276 45124 9332 45180
rect 9332 45124 9336 45180
rect 9272 45120 9336 45124
rect 9352 45180 9416 45184
rect 9352 45124 9356 45180
rect 9356 45124 9412 45180
rect 9412 45124 9416 45180
rect 9352 45120 9416 45124
rect 3372 44644 3436 44708
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 7480 44636 7544 44640
rect 7480 44580 7484 44636
rect 7484 44580 7540 44636
rect 7540 44580 7544 44636
rect 7480 44576 7544 44580
rect 7560 44636 7624 44640
rect 7560 44580 7564 44636
rect 7564 44580 7620 44636
rect 7620 44580 7624 44636
rect 7560 44576 7624 44580
rect 7640 44636 7704 44640
rect 7640 44580 7644 44636
rect 7644 44580 7700 44636
rect 7700 44580 7704 44636
rect 7640 44576 7704 44580
rect 7720 44636 7784 44640
rect 7720 44580 7724 44636
rect 7724 44580 7780 44636
rect 7780 44580 7784 44636
rect 7720 44576 7784 44580
rect 428 44372 492 44436
rect 612 44372 676 44436
rect 980 44372 1044 44436
rect 3372 44372 3436 44436
rect 1164 44236 1228 44300
rect 2584 44092 2648 44096
rect 2584 44036 2588 44092
rect 2588 44036 2644 44092
rect 2644 44036 2648 44092
rect 2584 44032 2648 44036
rect 2664 44092 2728 44096
rect 2664 44036 2668 44092
rect 2668 44036 2724 44092
rect 2724 44036 2728 44092
rect 2664 44032 2728 44036
rect 2744 44092 2808 44096
rect 2744 44036 2748 44092
rect 2748 44036 2804 44092
rect 2804 44036 2808 44092
rect 2744 44032 2808 44036
rect 2824 44092 2888 44096
rect 2824 44036 2828 44092
rect 2828 44036 2884 44092
rect 2884 44036 2888 44092
rect 2824 44032 2888 44036
rect 5848 44092 5912 44096
rect 5848 44036 5852 44092
rect 5852 44036 5908 44092
rect 5908 44036 5912 44092
rect 5848 44032 5912 44036
rect 5928 44092 5992 44096
rect 5928 44036 5932 44092
rect 5932 44036 5988 44092
rect 5988 44036 5992 44092
rect 5928 44032 5992 44036
rect 6008 44092 6072 44096
rect 6008 44036 6012 44092
rect 6012 44036 6068 44092
rect 6068 44036 6072 44092
rect 6008 44032 6072 44036
rect 6088 44092 6152 44096
rect 6088 44036 6092 44092
rect 6092 44036 6148 44092
rect 6148 44036 6152 44092
rect 6088 44032 6152 44036
rect 9112 44092 9176 44096
rect 9112 44036 9116 44092
rect 9116 44036 9172 44092
rect 9172 44036 9176 44092
rect 9112 44032 9176 44036
rect 9192 44092 9256 44096
rect 9192 44036 9196 44092
rect 9196 44036 9252 44092
rect 9252 44036 9256 44092
rect 9192 44032 9256 44036
rect 9272 44092 9336 44096
rect 9272 44036 9276 44092
rect 9276 44036 9332 44092
rect 9332 44036 9336 44092
rect 9272 44032 9336 44036
rect 9352 44092 9416 44096
rect 9352 44036 9356 44092
rect 9356 44036 9412 44092
rect 9412 44036 9416 44092
rect 9352 44032 9416 44036
rect 2084 43828 2148 43892
rect 1532 43692 1596 43756
rect 2084 43692 2148 43756
rect 1532 43420 1596 43484
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 7480 43548 7544 43552
rect 7480 43492 7484 43548
rect 7484 43492 7540 43548
rect 7540 43492 7544 43548
rect 7480 43488 7544 43492
rect 7560 43548 7624 43552
rect 7560 43492 7564 43548
rect 7564 43492 7620 43548
rect 7620 43492 7624 43548
rect 7560 43488 7624 43492
rect 7640 43548 7704 43552
rect 7640 43492 7644 43548
rect 7644 43492 7700 43548
rect 7700 43492 7704 43548
rect 7640 43488 7704 43492
rect 7720 43548 7784 43552
rect 7720 43492 7724 43548
rect 7724 43492 7780 43548
rect 7780 43492 7784 43548
rect 7720 43488 7784 43492
rect 3556 43148 3620 43212
rect 1900 43012 1964 43076
rect 2584 43004 2648 43008
rect 2584 42948 2588 43004
rect 2588 42948 2644 43004
rect 2644 42948 2648 43004
rect 2584 42944 2648 42948
rect 2664 43004 2728 43008
rect 2664 42948 2668 43004
rect 2668 42948 2724 43004
rect 2724 42948 2728 43004
rect 2664 42944 2728 42948
rect 2744 43004 2808 43008
rect 2744 42948 2748 43004
rect 2748 42948 2804 43004
rect 2804 42948 2808 43004
rect 2744 42944 2808 42948
rect 2824 43004 2888 43008
rect 2824 42948 2828 43004
rect 2828 42948 2884 43004
rect 2884 42948 2888 43004
rect 2824 42944 2888 42948
rect 1900 42936 1964 42940
rect 1900 42880 1950 42936
rect 1950 42880 1964 42936
rect 1900 42876 1964 42880
rect 1348 42800 1412 42804
rect 1348 42744 1362 42800
rect 1362 42744 1412 42800
rect 1348 42740 1412 42744
rect 1716 42740 1780 42804
rect 3188 43012 3252 43076
rect 5848 43004 5912 43008
rect 5848 42948 5852 43004
rect 5852 42948 5908 43004
rect 5908 42948 5912 43004
rect 5848 42944 5912 42948
rect 5928 43004 5992 43008
rect 5928 42948 5932 43004
rect 5932 42948 5988 43004
rect 5988 42948 5992 43004
rect 5928 42944 5992 42948
rect 6008 43004 6072 43008
rect 6008 42948 6012 43004
rect 6012 42948 6068 43004
rect 6068 42948 6072 43004
rect 6008 42944 6072 42948
rect 6088 43004 6152 43008
rect 6088 42948 6092 43004
rect 6092 42948 6148 43004
rect 6148 42948 6152 43004
rect 6088 42944 6152 42948
rect 9112 43004 9176 43008
rect 9112 42948 9116 43004
rect 9116 42948 9172 43004
rect 9172 42948 9176 43004
rect 9112 42944 9176 42948
rect 9192 43004 9256 43008
rect 9192 42948 9196 43004
rect 9196 42948 9252 43004
rect 9252 42948 9256 43004
rect 9192 42944 9256 42948
rect 9272 43004 9336 43008
rect 9272 42948 9276 43004
rect 9276 42948 9332 43004
rect 9332 42948 9336 43004
rect 9272 42944 9336 42948
rect 9352 43004 9416 43008
rect 9352 42948 9356 43004
rect 9356 42948 9412 43004
rect 9412 42948 9416 43004
rect 9352 42944 9416 42948
rect 3188 42876 3252 42940
rect 3924 42740 3988 42804
rect 1348 42604 1412 42668
rect 2084 42604 2148 42668
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 7480 42460 7544 42464
rect 7480 42404 7484 42460
rect 7484 42404 7540 42460
rect 7540 42404 7544 42460
rect 7480 42400 7544 42404
rect 7560 42460 7624 42464
rect 7560 42404 7564 42460
rect 7564 42404 7620 42460
rect 7620 42404 7624 42460
rect 7560 42400 7624 42404
rect 7640 42460 7704 42464
rect 7640 42404 7644 42460
rect 7644 42404 7700 42460
rect 7700 42404 7704 42460
rect 7640 42400 7704 42404
rect 7720 42460 7784 42464
rect 7720 42404 7724 42460
rect 7724 42404 7780 42460
rect 7780 42404 7784 42460
rect 7720 42400 7784 42404
rect 1716 42392 1780 42396
rect 1716 42336 1766 42392
rect 1766 42336 1780 42392
rect 1716 42332 1780 42336
rect 5396 42060 5460 42124
rect 3372 41924 3436 41988
rect 4844 41924 4908 41988
rect 5396 41924 5460 41988
rect 2584 41916 2648 41920
rect 2584 41860 2588 41916
rect 2588 41860 2644 41916
rect 2644 41860 2648 41916
rect 2584 41856 2648 41860
rect 2664 41916 2728 41920
rect 2664 41860 2668 41916
rect 2668 41860 2724 41916
rect 2724 41860 2728 41916
rect 2664 41856 2728 41860
rect 2744 41916 2808 41920
rect 2744 41860 2748 41916
rect 2748 41860 2804 41916
rect 2804 41860 2808 41916
rect 2744 41856 2808 41860
rect 2824 41916 2888 41920
rect 2824 41860 2828 41916
rect 2828 41860 2884 41916
rect 2884 41860 2888 41916
rect 2824 41856 2888 41860
rect 5848 41916 5912 41920
rect 5848 41860 5852 41916
rect 5852 41860 5908 41916
rect 5908 41860 5912 41916
rect 5848 41856 5912 41860
rect 5928 41916 5992 41920
rect 5928 41860 5932 41916
rect 5932 41860 5988 41916
rect 5988 41860 5992 41916
rect 5928 41856 5992 41860
rect 6008 41916 6072 41920
rect 6008 41860 6012 41916
rect 6012 41860 6068 41916
rect 6068 41860 6072 41916
rect 6008 41856 6072 41860
rect 6088 41916 6152 41920
rect 6088 41860 6092 41916
rect 6092 41860 6148 41916
rect 6148 41860 6152 41916
rect 6088 41856 6152 41860
rect 9112 41916 9176 41920
rect 9112 41860 9116 41916
rect 9116 41860 9172 41916
rect 9172 41860 9176 41916
rect 9112 41856 9176 41860
rect 9192 41916 9256 41920
rect 9192 41860 9196 41916
rect 9196 41860 9252 41916
rect 9252 41860 9256 41916
rect 9192 41856 9256 41860
rect 9272 41916 9336 41920
rect 9272 41860 9276 41916
rect 9276 41860 9332 41916
rect 9332 41860 9336 41916
rect 9272 41856 9336 41860
rect 9352 41916 9416 41920
rect 9352 41860 9356 41916
rect 9356 41860 9412 41916
rect 9412 41860 9416 41916
rect 9352 41856 9416 41860
rect 2084 41788 2148 41852
rect 1348 41576 1412 41580
rect 1348 41520 1362 41576
rect 1362 41520 1412 41576
rect 1348 41516 1412 41520
rect 3740 41516 3804 41580
rect 5028 41516 5092 41580
rect 60 41380 124 41444
rect 3188 41380 3252 41444
rect 3924 41380 3988 41444
rect 4844 41380 4908 41444
rect 5212 41380 5276 41444
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 7480 41372 7544 41376
rect 7480 41316 7484 41372
rect 7484 41316 7540 41372
rect 7540 41316 7544 41372
rect 7480 41312 7544 41316
rect 7560 41372 7624 41376
rect 7560 41316 7564 41372
rect 7564 41316 7620 41372
rect 7620 41316 7624 41372
rect 7560 41312 7624 41316
rect 7640 41372 7704 41376
rect 7640 41316 7644 41372
rect 7644 41316 7700 41372
rect 7700 41316 7704 41372
rect 7640 41312 7704 41316
rect 7720 41372 7784 41376
rect 7720 41316 7724 41372
rect 7724 41316 7780 41372
rect 7780 41316 7784 41372
rect 7720 41312 7784 41316
rect 1348 41244 1412 41308
rect 1716 41244 1780 41308
rect 3556 41304 3620 41308
rect 3556 41248 3606 41304
rect 3606 41248 3620 41304
rect 3556 41244 3620 41248
rect 5212 41304 5276 41308
rect 5212 41248 5262 41304
rect 5262 41248 5276 41304
rect 3372 41108 3436 41172
rect 3372 41032 3436 41036
rect 3372 40976 3422 41032
rect 3422 40976 3436 41032
rect 3372 40972 3436 40976
rect 3556 40972 3620 41036
rect 5212 41244 5276 41248
rect 2584 40828 2648 40832
rect 2584 40772 2588 40828
rect 2588 40772 2644 40828
rect 2644 40772 2648 40828
rect 2584 40768 2648 40772
rect 2664 40828 2728 40832
rect 2664 40772 2668 40828
rect 2668 40772 2724 40828
rect 2724 40772 2728 40828
rect 2664 40768 2728 40772
rect 2744 40828 2808 40832
rect 2744 40772 2748 40828
rect 2748 40772 2804 40828
rect 2804 40772 2808 40828
rect 2744 40768 2808 40772
rect 2824 40828 2888 40832
rect 2824 40772 2828 40828
rect 2828 40772 2884 40828
rect 2884 40772 2888 40828
rect 2824 40768 2888 40772
rect 5848 40828 5912 40832
rect 5848 40772 5852 40828
rect 5852 40772 5908 40828
rect 5908 40772 5912 40828
rect 5848 40768 5912 40772
rect 5928 40828 5992 40832
rect 5928 40772 5932 40828
rect 5932 40772 5988 40828
rect 5988 40772 5992 40828
rect 5928 40768 5992 40772
rect 6008 40828 6072 40832
rect 6008 40772 6012 40828
rect 6012 40772 6068 40828
rect 6068 40772 6072 40828
rect 6008 40768 6072 40772
rect 6088 40828 6152 40832
rect 6088 40772 6092 40828
rect 6092 40772 6148 40828
rect 6148 40772 6152 40828
rect 6088 40768 6152 40772
rect 9112 40828 9176 40832
rect 9112 40772 9116 40828
rect 9116 40772 9172 40828
rect 9172 40772 9176 40828
rect 9112 40768 9176 40772
rect 9192 40828 9256 40832
rect 9192 40772 9196 40828
rect 9196 40772 9252 40828
rect 9252 40772 9256 40828
rect 9192 40768 9256 40772
rect 9272 40828 9336 40832
rect 9272 40772 9276 40828
rect 9276 40772 9332 40828
rect 9332 40772 9336 40828
rect 9272 40768 9336 40772
rect 9352 40828 9416 40832
rect 9352 40772 9356 40828
rect 9356 40772 9412 40828
rect 9412 40772 9416 40828
rect 9352 40768 9416 40772
rect 2406 40428 2470 40492
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 7480 40284 7544 40288
rect 7480 40228 7484 40284
rect 7484 40228 7540 40284
rect 7540 40228 7544 40284
rect 7480 40224 7544 40228
rect 7560 40284 7624 40288
rect 7560 40228 7564 40284
rect 7564 40228 7620 40284
rect 7620 40228 7624 40284
rect 7560 40224 7624 40228
rect 7640 40284 7704 40288
rect 7640 40228 7644 40284
rect 7644 40228 7700 40284
rect 7700 40228 7704 40284
rect 7640 40224 7704 40228
rect 7720 40284 7784 40288
rect 7720 40228 7724 40284
rect 7724 40228 7780 40284
rect 7780 40228 7784 40284
rect 7720 40224 7784 40228
rect 5396 39884 5460 39948
rect 2584 39740 2648 39744
rect 2584 39684 2588 39740
rect 2588 39684 2644 39740
rect 2644 39684 2648 39740
rect 2584 39680 2648 39684
rect 2664 39740 2728 39744
rect 2664 39684 2668 39740
rect 2668 39684 2724 39740
rect 2724 39684 2728 39740
rect 2664 39680 2728 39684
rect 2744 39740 2808 39744
rect 2744 39684 2748 39740
rect 2748 39684 2804 39740
rect 2804 39684 2808 39740
rect 2744 39680 2808 39684
rect 2824 39740 2888 39744
rect 2824 39684 2828 39740
rect 2828 39684 2884 39740
rect 2884 39684 2888 39740
rect 2824 39680 2888 39684
rect 5848 39740 5912 39744
rect 5848 39684 5852 39740
rect 5852 39684 5908 39740
rect 5908 39684 5912 39740
rect 5848 39680 5912 39684
rect 5928 39740 5992 39744
rect 5928 39684 5932 39740
rect 5932 39684 5988 39740
rect 5988 39684 5992 39740
rect 5928 39680 5992 39684
rect 6008 39740 6072 39744
rect 6008 39684 6012 39740
rect 6012 39684 6068 39740
rect 6068 39684 6072 39740
rect 6008 39680 6072 39684
rect 6088 39740 6152 39744
rect 6088 39684 6092 39740
rect 6092 39684 6148 39740
rect 6148 39684 6152 39740
rect 6088 39680 6152 39684
rect 9112 39740 9176 39744
rect 9112 39684 9116 39740
rect 9116 39684 9172 39740
rect 9172 39684 9176 39740
rect 9112 39680 9176 39684
rect 9192 39740 9256 39744
rect 9192 39684 9196 39740
rect 9196 39684 9252 39740
rect 9252 39684 9256 39740
rect 9192 39680 9256 39684
rect 9272 39740 9336 39744
rect 9272 39684 9276 39740
rect 9276 39684 9332 39740
rect 9332 39684 9336 39740
rect 9272 39680 9336 39684
rect 9352 39740 9416 39744
rect 9352 39684 9356 39740
rect 9356 39684 9412 39740
rect 9412 39684 9416 39740
rect 9352 39680 9416 39684
rect 3924 39476 3988 39540
rect 6500 39476 6564 39540
rect 1716 39340 1780 39404
rect 3188 39204 3252 39268
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 7480 39196 7544 39200
rect 7480 39140 7484 39196
rect 7484 39140 7540 39196
rect 7540 39140 7544 39196
rect 7480 39136 7544 39140
rect 7560 39196 7624 39200
rect 7560 39140 7564 39196
rect 7564 39140 7620 39196
rect 7620 39140 7624 39196
rect 7560 39136 7624 39140
rect 7640 39196 7704 39200
rect 7640 39140 7644 39196
rect 7644 39140 7700 39196
rect 7700 39140 7704 39196
rect 7640 39136 7704 39140
rect 7720 39196 7784 39200
rect 7720 39140 7724 39196
rect 7724 39140 7780 39196
rect 7780 39140 7784 39196
rect 7720 39136 7784 39140
rect 2084 38932 2148 38996
rect 6316 38932 6380 38996
rect 428 38796 492 38860
rect 2084 38796 2148 38860
rect 3556 38796 3620 38860
rect 2584 38652 2648 38656
rect 2584 38596 2588 38652
rect 2588 38596 2644 38652
rect 2644 38596 2648 38652
rect 2584 38592 2648 38596
rect 2664 38652 2728 38656
rect 2664 38596 2668 38652
rect 2668 38596 2724 38652
rect 2724 38596 2728 38652
rect 2664 38592 2728 38596
rect 2744 38652 2808 38656
rect 2744 38596 2748 38652
rect 2748 38596 2804 38652
rect 2804 38596 2808 38652
rect 2744 38592 2808 38596
rect 2824 38652 2888 38656
rect 2824 38596 2828 38652
rect 2828 38596 2884 38652
rect 2884 38596 2888 38652
rect 2824 38592 2888 38596
rect 5848 38652 5912 38656
rect 5848 38596 5852 38652
rect 5852 38596 5908 38652
rect 5908 38596 5912 38652
rect 5848 38592 5912 38596
rect 5928 38652 5992 38656
rect 5928 38596 5932 38652
rect 5932 38596 5988 38652
rect 5988 38596 5992 38652
rect 5928 38592 5992 38596
rect 6008 38652 6072 38656
rect 6008 38596 6012 38652
rect 6012 38596 6068 38652
rect 6068 38596 6072 38652
rect 6008 38592 6072 38596
rect 6088 38652 6152 38656
rect 6088 38596 6092 38652
rect 6092 38596 6148 38652
rect 6148 38596 6152 38652
rect 6088 38592 6152 38596
rect 9112 38652 9176 38656
rect 9112 38596 9116 38652
rect 9116 38596 9172 38652
rect 9172 38596 9176 38652
rect 9112 38592 9176 38596
rect 9192 38652 9256 38656
rect 9192 38596 9196 38652
rect 9196 38596 9252 38652
rect 9252 38596 9256 38652
rect 9192 38592 9256 38596
rect 9272 38652 9336 38656
rect 9272 38596 9276 38652
rect 9276 38596 9332 38652
rect 9332 38596 9336 38652
rect 9272 38592 9336 38596
rect 9352 38652 9416 38656
rect 9352 38596 9356 38652
rect 9356 38596 9412 38652
rect 9412 38596 9416 38652
rect 9352 38592 9416 38596
rect 3188 38252 3252 38316
rect 2084 38116 2148 38180
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 3372 37844 3436 37908
rect 7480 38108 7544 38112
rect 7480 38052 7484 38108
rect 7484 38052 7540 38108
rect 7540 38052 7544 38108
rect 7480 38048 7544 38052
rect 7560 38108 7624 38112
rect 7560 38052 7564 38108
rect 7564 38052 7620 38108
rect 7620 38052 7624 38108
rect 7560 38048 7624 38052
rect 7640 38108 7704 38112
rect 7640 38052 7644 38108
rect 7644 38052 7700 38108
rect 7700 38052 7704 38108
rect 7640 38048 7704 38052
rect 7720 38108 7784 38112
rect 7720 38052 7724 38108
rect 7724 38052 7780 38108
rect 7780 38052 7784 38108
rect 7720 38048 7784 38052
rect 2584 37564 2648 37568
rect 2584 37508 2588 37564
rect 2588 37508 2644 37564
rect 2644 37508 2648 37564
rect 2584 37504 2648 37508
rect 2664 37564 2728 37568
rect 2664 37508 2668 37564
rect 2668 37508 2724 37564
rect 2724 37508 2728 37564
rect 2664 37504 2728 37508
rect 2744 37564 2808 37568
rect 2744 37508 2748 37564
rect 2748 37508 2804 37564
rect 2804 37508 2808 37564
rect 2744 37504 2808 37508
rect 2824 37564 2888 37568
rect 2824 37508 2828 37564
rect 2828 37508 2884 37564
rect 2884 37508 2888 37564
rect 2824 37504 2888 37508
rect 5848 37564 5912 37568
rect 5848 37508 5852 37564
rect 5852 37508 5908 37564
rect 5908 37508 5912 37564
rect 5848 37504 5912 37508
rect 5928 37564 5992 37568
rect 5928 37508 5932 37564
rect 5932 37508 5988 37564
rect 5988 37508 5992 37564
rect 5928 37504 5992 37508
rect 6008 37564 6072 37568
rect 6008 37508 6012 37564
rect 6012 37508 6068 37564
rect 6068 37508 6072 37564
rect 6008 37504 6072 37508
rect 6088 37564 6152 37568
rect 6088 37508 6092 37564
rect 6092 37508 6148 37564
rect 6148 37508 6152 37564
rect 6088 37504 6152 37508
rect 9112 37564 9176 37568
rect 9112 37508 9116 37564
rect 9116 37508 9172 37564
rect 9172 37508 9176 37564
rect 9112 37504 9176 37508
rect 9192 37564 9256 37568
rect 9192 37508 9196 37564
rect 9196 37508 9252 37564
rect 9252 37508 9256 37564
rect 9192 37504 9256 37508
rect 9272 37564 9336 37568
rect 9272 37508 9276 37564
rect 9276 37508 9332 37564
rect 9332 37508 9336 37564
rect 9272 37504 9336 37508
rect 9352 37564 9416 37568
rect 9352 37508 9356 37564
rect 9356 37508 9412 37564
rect 9412 37508 9416 37564
rect 9352 37504 9416 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 7480 37020 7544 37024
rect 7480 36964 7484 37020
rect 7484 36964 7540 37020
rect 7540 36964 7544 37020
rect 7480 36960 7544 36964
rect 7560 37020 7624 37024
rect 7560 36964 7564 37020
rect 7564 36964 7620 37020
rect 7620 36964 7624 37020
rect 7560 36960 7624 36964
rect 7640 37020 7704 37024
rect 7640 36964 7644 37020
rect 7644 36964 7700 37020
rect 7700 36964 7704 37020
rect 7640 36960 7704 36964
rect 7720 37020 7784 37024
rect 7720 36964 7724 37020
rect 7724 36964 7780 37020
rect 7780 36964 7784 37020
rect 7720 36960 7784 36964
rect 2268 36756 2332 36820
rect 2268 36544 2332 36548
rect 5028 36756 5092 36820
rect 2268 36488 2318 36544
rect 2318 36488 2332 36544
rect 2268 36484 2332 36488
rect 2584 36476 2648 36480
rect 2584 36420 2588 36476
rect 2588 36420 2644 36476
rect 2644 36420 2648 36476
rect 2584 36416 2648 36420
rect 2664 36476 2728 36480
rect 2664 36420 2668 36476
rect 2668 36420 2724 36476
rect 2724 36420 2728 36476
rect 2664 36416 2728 36420
rect 2744 36476 2808 36480
rect 2744 36420 2748 36476
rect 2748 36420 2804 36476
rect 2804 36420 2808 36476
rect 2744 36416 2808 36420
rect 2824 36476 2888 36480
rect 2824 36420 2828 36476
rect 2828 36420 2884 36476
rect 2884 36420 2888 36476
rect 2824 36416 2888 36420
rect 5848 36476 5912 36480
rect 5848 36420 5852 36476
rect 5852 36420 5908 36476
rect 5908 36420 5912 36476
rect 5848 36416 5912 36420
rect 5928 36476 5992 36480
rect 5928 36420 5932 36476
rect 5932 36420 5988 36476
rect 5988 36420 5992 36476
rect 5928 36416 5992 36420
rect 6008 36476 6072 36480
rect 6008 36420 6012 36476
rect 6012 36420 6068 36476
rect 6068 36420 6072 36476
rect 6008 36416 6072 36420
rect 6088 36476 6152 36480
rect 6088 36420 6092 36476
rect 6092 36420 6148 36476
rect 6148 36420 6152 36476
rect 6088 36416 6152 36420
rect 9112 36476 9176 36480
rect 9112 36420 9116 36476
rect 9116 36420 9172 36476
rect 9172 36420 9176 36476
rect 9112 36416 9176 36420
rect 9192 36476 9256 36480
rect 9192 36420 9196 36476
rect 9196 36420 9252 36476
rect 9252 36420 9256 36476
rect 9192 36416 9256 36420
rect 9272 36476 9336 36480
rect 9272 36420 9276 36476
rect 9276 36420 9332 36476
rect 9332 36420 9336 36476
rect 9272 36416 9336 36420
rect 9352 36476 9416 36480
rect 9352 36420 9356 36476
rect 9356 36420 9412 36476
rect 9412 36420 9416 36476
rect 9352 36416 9416 36420
rect 1900 36076 1964 36140
rect 5028 35940 5092 36004
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 7480 35932 7544 35936
rect 7480 35876 7484 35932
rect 7484 35876 7540 35932
rect 7540 35876 7544 35932
rect 7480 35872 7544 35876
rect 7560 35932 7624 35936
rect 7560 35876 7564 35932
rect 7564 35876 7620 35932
rect 7620 35876 7624 35932
rect 7560 35872 7624 35876
rect 7640 35932 7704 35936
rect 7640 35876 7644 35932
rect 7644 35876 7700 35932
rect 7700 35876 7704 35932
rect 7640 35872 7704 35876
rect 7720 35932 7784 35936
rect 7720 35876 7724 35932
rect 7724 35876 7780 35932
rect 7780 35876 7784 35932
rect 7720 35872 7784 35876
rect 5396 35668 5460 35732
rect 2584 35388 2648 35392
rect 2584 35332 2588 35388
rect 2588 35332 2644 35388
rect 2644 35332 2648 35388
rect 2584 35328 2648 35332
rect 2664 35388 2728 35392
rect 2664 35332 2668 35388
rect 2668 35332 2724 35388
rect 2724 35332 2728 35388
rect 2664 35328 2728 35332
rect 2744 35388 2808 35392
rect 2744 35332 2748 35388
rect 2748 35332 2804 35388
rect 2804 35332 2808 35388
rect 2744 35328 2808 35332
rect 2824 35388 2888 35392
rect 2824 35332 2828 35388
rect 2828 35332 2884 35388
rect 2884 35332 2888 35388
rect 2824 35328 2888 35332
rect 5848 35388 5912 35392
rect 5848 35332 5852 35388
rect 5852 35332 5908 35388
rect 5908 35332 5912 35388
rect 5848 35328 5912 35332
rect 5928 35388 5992 35392
rect 5928 35332 5932 35388
rect 5932 35332 5988 35388
rect 5988 35332 5992 35388
rect 5928 35328 5992 35332
rect 6008 35388 6072 35392
rect 6008 35332 6012 35388
rect 6012 35332 6068 35388
rect 6068 35332 6072 35388
rect 6008 35328 6072 35332
rect 6088 35388 6152 35392
rect 6088 35332 6092 35388
rect 6092 35332 6148 35388
rect 6148 35332 6152 35388
rect 6088 35328 6152 35332
rect 9112 35388 9176 35392
rect 9112 35332 9116 35388
rect 9116 35332 9172 35388
rect 9172 35332 9176 35388
rect 9112 35328 9176 35332
rect 9192 35388 9256 35392
rect 9192 35332 9196 35388
rect 9196 35332 9252 35388
rect 9252 35332 9256 35388
rect 9192 35328 9256 35332
rect 9272 35388 9336 35392
rect 9272 35332 9276 35388
rect 9276 35332 9332 35388
rect 9332 35332 9336 35388
rect 9272 35328 9336 35332
rect 9352 35388 9416 35392
rect 9352 35332 9356 35388
rect 9356 35332 9412 35388
rect 9412 35332 9416 35388
rect 9352 35328 9416 35332
rect 3740 35320 3804 35324
rect 3740 35264 3790 35320
rect 3790 35264 3804 35320
rect 3740 35260 3804 35264
rect 3740 35184 3804 35188
rect 3740 35128 3754 35184
rect 3754 35128 3804 35184
rect 3740 35124 3804 35128
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 7480 34844 7544 34848
rect 7480 34788 7484 34844
rect 7484 34788 7540 34844
rect 7540 34788 7544 34844
rect 7480 34784 7544 34788
rect 7560 34844 7624 34848
rect 7560 34788 7564 34844
rect 7564 34788 7620 34844
rect 7620 34788 7624 34844
rect 7560 34784 7624 34788
rect 7640 34844 7704 34848
rect 7640 34788 7644 34844
rect 7644 34788 7700 34844
rect 7700 34788 7704 34844
rect 7640 34784 7704 34788
rect 7720 34844 7784 34848
rect 7720 34788 7724 34844
rect 7724 34788 7780 34844
rect 7780 34788 7784 34844
rect 7720 34784 7784 34788
rect 2584 34300 2648 34304
rect 2584 34244 2588 34300
rect 2588 34244 2644 34300
rect 2644 34244 2648 34300
rect 2584 34240 2648 34244
rect 2664 34300 2728 34304
rect 2664 34244 2668 34300
rect 2668 34244 2724 34300
rect 2724 34244 2728 34300
rect 2664 34240 2728 34244
rect 2744 34300 2808 34304
rect 2744 34244 2748 34300
rect 2748 34244 2804 34300
rect 2804 34244 2808 34300
rect 2744 34240 2808 34244
rect 2824 34300 2888 34304
rect 2824 34244 2828 34300
rect 2828 34244 2884 34300
rect 2884 34244 2888 34300
rect 2824 34240 2888 34244
rect 5848 34300 5912 34304
rect 5848 34244 5852 34300
rect 5852 34244 5908 34300
rect 5908 34244 5912 34300
rect 5848 34240 5912 34244
rect 5928 34300 5992 34304
rect 5928 34244 5932 34300
rect 5932 34244 5988 34300
rect 5988 34244 5992 34300
rect 5928 34240 5992 34244
rect 6008 34300 6072 34304
rect 6008 34244 6012 34300
rect 6012 34244 6068 34300
rect 6068 34244 6072 34300
rect 6008 34240 6072 34244
rect 6088 34300 6152 34304
rect 6088 34244 6092 34300
rect 6092 34244 6148 34300
rect 6148 34244 6152 34300
rect 6088 34240 6152 34244
rect 9112 34300 9176 34304
rect 9112 34244 9116 34300
rect 9116 34244 9172 34300
rect 9172 34244 9176 34300
rect 9112 34240 9176 34244
rect 9192 34300 9256 34304
rect 9192 34244 9196 34300
rect 9196 34244 9252 34300
rect 9252 34244 9256 34300
rect 9192 34240 9256 34244
rect 9272 34300 9336 34304
rect 9272 34244 9276 34300
rect 9276 34244 9332 34300
rect 9332 34244 9336 34300
rect 9272 34240 9336 34244
rect 9352 34300 9416 34304
rect 9352 34244 9356 34300
rect 9356 34244 9412 34300
rect 9412 34244 9416 34300
rect 9352 34240 9416 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 7480 33756 7544 33760
rect 7480 33700 7484 33756
rect 7484 33700 7540 33756
rect 7540 33700 7544 33756
rect 7480 33696 7544 33700
rect 7560 33756 7624 33760
rect 7560 33700 7564 33756
rect 7564 33700 7620 33756
rect 7620 33700 7624 33756
rect 7560 33696 7624 33700
rect 7640 33756 7704 33760
rect 7640 33700 7644 33756
rect 7644 33700 7700 33756
rect 7700 33700 7704 33756
rect 7640 33696 7704 33700
rect 7720 33756 7784 33760
rect 7720 33700 7724 33756
rect 7724 33700 7780 33756
rect 7780 33700 7784 33756
rect 7720 33696 7784 33700
rect 1348 33220 1412 33284
rect 2584 33212 2648 33216
rect 2584 33156 2588 33212
rect 2588 33156 2644 33212
rect 2644 33156 2648 33212
rect 2584 33152 2648 33156
rect 2664 33212 2728 33216
rect 2664 33156 2668 33212
rect 2668 33156 2724 33212
rect 2724 33156 2728 33212
rect 2664 33152 2728 33156
rect 2744 33212 2808 33216
rect 2744 33156 2748 33212
rect 2748 33156 2804 33212
rect 2804 33156 2808 33212
rect 2744 33152 2808 33156
rect 2824 33212 2888 33216
rect 2824 33156 2828 33212
rect 2828 33156 2884 33212
rect 2884 33156 2888 33212
rect 2824 33152 2888 33156
rect 5848 33212 5912 33216
rect 5848 33156 5852 33212
rect 5852 33156 5908 33212
rect 5908 33156 5912 33212
rect 5848 33152 5912 33156
rect 5928 33212 5992 33216
rect 5928 33156 5932 33212
rect 5932 33156 5988 33212
rect 5988 33156 5992 33212
rect 5928 33152 5992 33156
rect 6008 33212 6072 33216
rect 6008 33156 6012 33212
rect 6012 33156 6068 33212
rect 6068 33156 6072 33212
rect 6008 33152 6072 33156
rect 6088 33212 6152 33216
rect 6088 33156 6092 33212
rect 6092 33156 6148 33212
rect 6148 33156 6152 33212
rect 6088 33152 6152 33156
rect 9112 33212 9176 33216
rect 9112 33156 9116 33212
rect 9116 33156 9172 33212
rect 9172 33156 9176 33212
rect 9112 33152 9176 33156
rect 9192 33212 9256 33216
rect 9192 33156 9196 33212
rect 9196 33156 9252 33212
rect 9252 33156 9256 33212
rect 9192 33152 9256 33156
rect 9272 33212 9336 33216
rect 9272 33156 9276 33212
rect 9276 33156 9332 33212
rect 9332 33156 9336 33212
rect 9272 33152 9336 33156
rect 9352 33212 9416 33216
rect 9352 33156 9356 33212
rect 9356 33156 9412 33212
rect 9412 33156 9416 33212
rect 9352 33152 9416 33156
rect 796 32872 860 32876
rect 796 32816 810 32872
rect 810 32816 860 32872
rect 796 32812 860 32816
rect 1164 32812 1228 32876
rect 1532 32676 1596 32740
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 7480 32668 7544 32672
rect 7480 32612 7484 32668
rect 7484 32612 7540 32668
rect 7540 32612 7544 32668
rect 7480 32608 7544 32612
rect 7560 32668 7624 32672
rect 7560 32612 7564 32668
rect 7564 32612 7620 32668
rect 7620 32612 7624 32668
rect 7560 32608 7624 32612
rect 7640 32668 7704 32672
rect 7640 32612 7644 32668
rect 7644 32612 7700 32668
rect 7700 32612 7704 32668
rect 7640 32608 7704 32612
rect 7720 32668 7784 32672
rect 7720 32612 7724 32668
rect 7724 32612 7780 32668
rect 7780 32612 7784 32668
rect 7720 32608 7784 32612
rect 3924 32404 3988 32468
rect 1716 32192 1780 32196
rect 1716 32136 1730 32192
rect 1730 32136 1780 32192
rect 1716 32132 1780 32136
rect 2584 32124 2648 32128
rect 2584 32068 2588 32124
rect 2588 32068 2644 32124
rect 2644 32068 2648 32124
rect 2584 32064 2648 32068
rect 2664 32124 2728 32128
rect 2664 32068 2668 32124
rect 2668 32068 2724 32124
rect 2724 32068 2728 32124
rect 2664 32064 2728 32068
rect 2744 32124 2808 32128
rect 2744 32068 2748 32124
rect 2748 32068 2804 32124
rect 2804 32068 2808 32124
rect 2744 32064 2808 32068
rect 2824 32124 2888 32128
rect 2824 32068 2828 32124
rect 2828 32068 2884 32124
rect 2884 32068 2888 32124
rect 2824 32064 2888 32068
rect 5848 32124 5912 32128
rect 5848 32068 5852 32124
rect 5852 32068 5908 32124
rect 5908 32068 5912 32124
rect 5848 32064 5912 32068
rect 5928 32124 5992 32128
rect 5928 32068 5932 32124
rect 5932 32068 5988 32124
rect 5988 32068 5992 32124
rect 5928 32064 5992 32068
rect 6008 32124 6072 32128
rect 6008 32068 6012 32124
rect 6012 32068 6068 32124
rect 6068 32068 6072 32124
rect 6008 32064 6072 32068
rect 6088 32124 6152 32128
rect 6088 32068 6092 32124
rect 6092 32068 6148 32124
rect 6148 32068 6152 32124
rect 6088 32064 6152 32068
rect 9112 32124 9176 32128
rect 9112 32068 9116 32124
rect 9116 32068 9172 32124
rect 9172 32068 9176 32124
rect 9112 32064 9176 32068
rect 9192 32124 9256 32128
rect 9192 32068 9196 32124
rect 9196 32068 9252 32124
rect 9252 32068 9256 32124
rect 9192 32064 9256 32068
rect 9272 32124 9336 32128
rect 9272 32068 9276 32124
rect 9276 32068 9332 32124
rect 9332 32068 9336 32124
rect 9272 32064 9336 32068
rect 9352 32124 9416 32128
rect 9352 32068 9356 32124
rect 9356 32068 9412 32124
rect 9412 32068 9416 32124
rect 9352 32064 9416 32068
rect 3556 31996 3620 32060
rect 3924 32056 3988 32060
rect 3924 32000 3974 32056
rect 3974 32000 3988 32056
rect 3924 31996 3988 32000
rect 1532 31860 1596 31924
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 1532 31512 1596 31516
rect 1532 31456 1546 31512
rect 1546 31456 1596 31512
rect 1532 31452 1596 31456
rect 7480 31580 7544 31584
rect 7480 31524 7484 31580
rect 7484 31524 7540 31580
rect 7540 31524 7544 31580
rect 7480 31520 7544 31524
rect 7560 31580 7624 31584
rect 7560 31524 7564 31580
rect 7564 31524 7620 31580
rect 7620 31524 7624 31580
rect 7560 31520 7624 31524
rect 7640 31580 7704 31584
rect 7640 31524 7644 31580
rect 7644 31524 7700 31580
rect 7700 31524 7704 31580
rect 7640 31520 7704 31524
rect 7720 31580 7784 31584
rect 7720 31524 7724 31580
rect 7724 31524 7780 31580
rect 7780 31524 7784 31580
rect 7720 31520 7784 31524
rect 5396 31044 5460 31108
rect 2584 31036 2648 31040
rect 2584 30980 2588 31036
rect 2588 30980 2644 31036
rect 2644 30980 2648 31036
rect 2584 30976 2648 30980
rect 2664 31036 2728 31040
rect 2664 30980 2668 31036
rect 2668 30980 2724 31036
rect 2724 30980 2728 31036
rect 2664 30976 2728 30980
rect 2744 31036 2808 31040
rect 2744 30980 2748 31036
rect 2748 30980 2804 31036
rect 2804 30980 2808 31036
rect 2744 30976 2808 30980
rect 2824 31036 2888 31040
rect 2824 30980 2828 31036
rect 2828 30980 2884 31036
rect 2884 30980 2888 31036
rect 2824 30976 2888 30980
rect 5848 31036 5912 31040
rect 5848 30980 5852 31036
rect 5852 30980 5908 31036
rect 5908 30980 5912 31036
rect 5848 30976 5912 30980
rect 5928 31036 5992 31040
rect 5928 30980 5932 31036
rect 5932 30980 5988 31036
rect 5988 30980 5992 31036
rect 5928 30976 5992 30980
rect 6008 31036 6072 31040
rect 6008 30980 6012 31036
rect 6012 30980 6068 31036
rect 6068 30980 6072 31036
rect 6008 30976 6072 30980
rect 6088 31036 6152 31040
rect 6088 30980 6092 31036
rect 6092 30980 6148 31036
rect 6148 30980 6152 31036
rect 6088 30976 6152 30980
rect 9112 31036 9176 31040
rect 9112 30980 9116 31036
rect 9116 30980 9172 31036
rect 9172 30980 9176 31036
rect 9112 30976 9176 30980
rect 9192 31036 9256 31040
rect 9192 30980 9196 31036
rect 9196 30980 9252 31036
rect 9252 30980 9256 31036
rect 9192 30976 9256 30980
rect 9272 31036 9336 31040
rect 9272 30980 9276 31036
rect 9276 30980 9332 31036
rect 9332 30980 9336 31036
rect 9272 30976 9336 30980
rect 9352 31036 9416 31040
rect 9352 30980 9356 31036
rect 9356 30980 9412 31036
rect 9412 30980 9416 31036
rect 9352 30976 9416 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 7480 30492 7544 30496
rect 7480 30436 7484 30492
rect 7484 30436 7540 30492
rect 7540 30436 7544 30492
rect 7480 30432 7544 30436
rect 7560 30492 7624 30496
rect 7560 30436 7564 30492
rect 7564 30436 7620 30492
rect 7620 30436 7624 30492
rect 7560 30432 7624 30436
rect 7640 30492 7704 30496
rect 7640 30436 7644 30492
rect 7644 30436 7700 30492
rect 7700 30436 7704 30492
rect 7640 30432 7704 30436
rect 7720 30492 7784 30496
rect 7720 30436 7724 30492
rect 7724 30436 7780 30492
rect 7780 30436 7784 30492
rect 7720 30432 7784 30436
rect 980 30228 1044 30292
rect 2584 29948 2648 29952
rect 2584 29892 2588 29948
rect 2588 29892 2644 29948
rect 2644 29892 2648 29948
rect 2584 29888 2648 29892
rect 2664 29948 2728 29952
rect 2664 29892 2668 29948
rect 2668 29892 2724 29948
rect 2724 29892 2728 29948
rect 2664 29888 2728 29892
rect 2744 29948 2808 29952
rect 2744 29892 2748 29948
rect 2748 29892 2804 29948
rect 2804 29892 2808 29948
rect 2744 29888 2808 29892
rect 2824 29948 2888 29952
rect 2824 29892 2828 29948
rect 2828 29892 2884 29948
rect 2884 29892 2888 29948
rect 2824 29888 2888 29892
rect 5848 29948 5912 29952
rect 5848 29892 5852 29948
rect 5852 29892 5908 29948
rect 5908 29892 5912 29948
rect 5848 29888 5912 29892
rect 5928 29948 5992 29952
rect 5928 29892 5932 29948
rect 5932 29892 5988 29948
rect 5988 29892 5992 29948
rect 5928 29888 5992 29892
rect 6008 29948 6072 29952
rect 6008 29892 6012 29948
rect 6012 29892 6068 29948
rect 6068 29892 6072 29948
rect 6008 29888 6072 29892
rect 6088 29948 6152 29952
rect 6088 29892 6092 29948
rect 6092 29892 6148 29948
rect 6148 29892 6152 29948
rect 6088 29888 6152 29892
rect 9112 29948 9176 29952
rect 9112 29892 9116 29948
rect 9116 29892 9172 29948
rect 9172 29892 9176 29948
rect 9112 29888 9176 29892
rect 9192 29948 9256 29952
rect 9192 29892 9196 29948
rect 9196 29892 9252 29948
rect 9252 29892 9256 29948
rect 9192 29888 9256 29892
rect 9272 29948 9336 29952
rect 9272 29892 9276 29948
rect 9276 29892 9332 29948
rect 9332 29892 9336 29948
rect 9272 29888 9336 29892
rect 9352 29948 9416 29952
rect 9352 29892 9356 29948
rect 9356 29892 9412 29948
rect 9412 29892 9416 29948
rect 9352 29888 9416 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 7480 29404 7544 29408
rect 7480 29348 7484 29404
rect 7484 29348 7540 29404
rect 7540 29348 7544 29404
rect 7480 29344 7544 29348
rect 7560 29404 7624 29408
rect 7560 29348 7564 29404
rect 7564 29348 7620 29404
rect 7620 29348 7624 29404
rect 7560 29344 7624 29348
rect 7640 29404 7704 29408
rect 7640 29348 7644 29404
rect 7644 29348 7700 29404
rect 7700 29348 7704 29404
rect 7640 29344 7704 29348
rect 7720 29404 7784 29408
rect 7720 29348 7724 29404
rect 7724 29348 7780 29404
rect 7780 29348 7784 29404
rect 7720 29344 7784 29348
rect 3372 29276 3436 29340
rect 2584 28860 2648 28864
rect 2584 28804 2588 28860
rect 2588 28804 2644 28860
rect 2644 28804 2648 28860
rect 2584 28800 2648 28804
rect 2664 28860 2728 28864
rect 2664 28804 2668 28860
rect 2668 28804 2724 28860
rect 2724 28804 2728 28860
rect 2664 28800 2728 28804
rect 2744 28860 2808 28864
rect 2744 28804 2748 28860
rect 2748 28804 2804 28860
rect 2804 28804 2808 28860
rect 2744 28800 2808 28804
rect 2824 28860 2888 28864
rect 2824 28804 2828 28860
rect 2828 28804 2884 28860
rect 2884 28804 2888 28860
rect 2824 28800 2888 28804
rect 5848 28860 5912 28864
rect 5848 28804 5852 28860
rect 5852 28804 5908 28860
rect 5908 28804 5912 28860
rect 5848 28800 5912 28804
rect 5928 28860 5992 28864
rect 5928 28804 5932 28860
rect 5932 28804 5988 28860
rect 5988 28804 5992 28860
rect 5928 28800 5992 28804
rect 6008 28860 6072 28864
rect 6008 28804 6012 28860
rect 6012 28804 6068 28860
rect 6068 28804 6072 28860
rect 6008 28800 6072 28804
rect 6088 28860 6152 28864
rect 6088 28804 6092 28860
rect 6092 28804 6148 28860
rect 6148 28804 6152 28860
rect 6088 28800 6152 28804
rect 9112 28860 9176 28864
rect 9112 28804 9116 28860
rect 9116 28804 9172 28860
rect 9172 28804 9176 28860
rect 9112 28800 9176 28804
rect 9192 28860 9256 28864
rect 9192 28804 9196 28860
rect 9196 28804 9252 28860
rect 9252 28804 9256 28860
rect 9192 28800 9256 28804
rect 9272 28860 9336 28864
rect 9272 28804 9276 28860
rect 9276 28804 9332 28860
rect 9332 28804 9336 28860
rect 9272 28800 9336 28804
rect 9352 28860 9416 28864
rect 9352 28804 9356 28860
rect 9356 28804 9412 28860
rect 9412 28804 9416 28860
rect 9352 28800 9416 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 7480 28316 7544 28320
rect 7480 28260 7484 28316
rect 7484 28260 7540 28316
rect 7540 28260 7544 28316
rect 7480 28256 7544 28260
rect 7560 28316 7624 28320
rect 7560 28260 7564 28316
rect 7564 28260 7620 28316
rect 7620 28260 7624 28316
rect 7560 28256 7624 28260
rect 7640 28316 7704 28320
rect 7640 28260 7644 28316
rect 7644 28260 7700 28316
rect 7700 28260 7704 28316
rect 7640 28256 7704 28260
rect 7720 28316 7784 28320
rect 7720 28260 7724 28316
rect 7724 28260 7780 28316
rect 7780 28260 7784 28316
rect 7720 28256 7784 28260
rect 2084 28188 2148 28252
rect 5028 28052 5092 28116
rect 2584 27772 2648 27776
rect 2584 27716 2588 27772
rect 2588 27716 2644 27772
rect 2644 27716 2648 27772
rect 2584 27712 2648 27716
rect 2664 27772 2728 27776
rect 2664 27716 2668 27772
rect 2668 27716 2724 27772
rect 2724 27716 2728 27772
rect 2664 27712 2728 27716
rect 2744 27772 2808 27776
rect 2744 27716 2748 27772
rect 2748 27716 2804 27772
rect 2804 27716 2808 27772
rect 2744 27712 2808 27716
rect 2824 27772 2888 27776
rect 2824 27716 2828 27772
rect 2828 27716 2884 27772
rect 2884 27716 2888 27772
rect 2824 27712 2888 27716
rect 5848 27772 5912 27776
rect 5848 27716 5852 27772
rect 5852 27716 5908 27772
rect 5908 27716 5912 27772
rect 5848 27712 5912 27716
rect 5928 27772 5992 27776
rect 5928 27716 5932 27772
rect 5932 27716 5988 27772
rect 5988 27716 5992 27772
rect 5928 27712 5992 27716
rect 6008 27772 6072 27776
rect 6008 27716 6012 27772
rect 6012 27716 6068 27772
rect 6068 27716 6072 27772
rect 6008 27712 6072 27716
rect 6088 27772 6152 27776
rect 6088 27716 6092 27772
rect 6092 27716 6148 27772
rect 6148 27716 6152 27772
rect 6088 27712 6152 27716
rect 9112 27772 9176 27776
rect 9112 27716 9116 27772
rect 9116 27716 9172 27772
rect 9172 27716 9176 27772
rect 9112 27712 9176 27716
rect 9192 27772 9256 27776
rect 9192 27716 9196 27772
rect 9196 27716 9252 27772
rect 9252 27716 9256 27772
rect 9192 27712 9256 27716
rect 9272 27772 9336 27776
rect 9272 27716 9276 27772
rect 9276 27716 9332 27772
rect 9332 27716 9336 27772
rect 9272 27712 9336 27716
rect 9352 27772 9416 27776
rect 9352 27716 9356 27772
rect 9356 27716 9412 27772
rect 9412 27716 9416 27772
rect 9352 27712 9416 27716
rect 3372 27644 3436 27708
rect 3556 27508 3620 27572
rect 3372 27372 3436 27436
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 7480 27228 7544 27232
rect 7480 27172 7484 27228
rect 7484 27172 7540 27228
rect 7540 27172 7544 27228
rect 7480 27168 7544 27172
rect 7560 27228 7624 27232
rect 7560 27172 7564 27228
rect 7564 27172 7620 27228
rect 7620 27172 7624 27228
rect 7560 27168 7624 27172
rect 7640 27228 7704 27232
rect 7640 27172 7644 27228
rect 7644 27172 7700 27228
rect 7700 27172 7704 27228
rect 7640 27168 7704 27172
rect 7720 27228 7784 27232
rect 7720 27172 7724 27228
rect 7724 27172 7780 27228
rect 7780 27172 7784 27228
rect 7720 27168 7784 27172
rect 2584 26684 2648 26688
rect 2584 26628 2588 26684
rect 2588 26628 2644 26684
rect 2644 26628 2648 26684
rect 2584 26624 2648 26628
rect 2664 26684 2728 26688
rect 2664 26628 2668 26684
rect 2668 26628 2724 26684
rect 2724 26628 2728 26684
rect 2664 26624 2728 26628
rect 2744 26684 2808 26688
rect 2744 26628 2748 26684
rect 2748 26628 2804 26684
rect 2804 26628 2808 26684
rect 2744 26624 2808 26628
rect 2824 26684 2888 26688
rect 2824 26628 2828 26684
rect 2828 26628 2884 26684
rect 2884 26628 2888 26684
rect 2824 26624 2888 26628
rect 5848 26684 5912 26688
rect 5848 26628 5852 26684
rect 5852 26628 5908 26684
rect 5908 26628 5912 26684
rect 5848 26624 5912 26628
rect 5928 26684 5992 26688
rect 5928 26628 5932 26684
rect 5932 26628 5988 26684
rect 5988 26628 5992 26684
rect 5928 26624 5992 26628
rect 6008 26684 6072 26688
rect 6008 26628 6012 26684
rect 6012 26628 6068 26684
rect 6068 26628 6072 26684
rect 6008 26624 6072 26628
rect 6088 26684 6152 26688
rect 6088 26628 6092 26684
rect 6092 26628 6148 26684
rect 6148 26628 6152 26684
rect 6088 26624 6152 26628
rect 9112 26684 9176 26688
rect 9112 26628 9116 26684
rect 9116 26628 9172 26684
rect 9172 26628 9176 26684
rect 9112 26624 9176 26628
rect 9192 26684 9256 26688
rect 9192 26628 9196 26684
rect 9196 26628 9252 26684
rect 9252 26628 9256 26684
rect 9192 26624 9256 26628
rect 9272 26684 9336 26688
rect 9272 26628 9276 26684
rect 9276 26628 9332 26684
rect 9332 26628 9336 26684
rect 9272 26624 9336 26628
rect 9352 26684 9416 26688
rect 9352 26628 9356 26684
rect 9356 26628 9412 26684
rect 9412 26628 9416 26684
rect 9352 26624 9416 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 7480 26140 7544 26144
rect 7480 26084 7484 26140
rect 7484 26084 7540 26140
rect 7540 26084 7544 26140
rect 7480 26080 7544 26084
rect 7560 26140 7624 26144
rect 7560 26084 7564 26140
rect 7564 26084 7620 26140
rect 7620 26084 7624 26140
rect 7560 26080 7624 26084
rect 7640 26140 7704 26144
rect 7640 26084 7644 26140
rect 7644 26084 7700 26140
rect 7700 26084 7704 26140
rect 7640 26080 7704 26084
rect 7720 26140 7784 26144
rect 7720 26084 7724 26140
rect 7724 26084 7780 26140
rect 7780 26084 7784 26140
rect 7720 26080 7784 26084
rect 5212 25876 5276 25940
rect 2584 25596 2648 25600
rect 2584 25540 2588 25596
rect 2588 25540 2644 25596
rect 2644 25540 2648 25596
rect 2584 25536 2648 25540
rect 2664 25596 2728 25600
rect 2664 25540 2668 25596
rect 2668 25540 2724 25596
rect 2724 25540 2728 25596
rect 2664 25536 2728 25540
rect 2744 25596 2808 25600
rect 2744 25540 2748 25596
rect 2748 25540 2804 25596
rect 2804 25540 2808 25596
rect 2744 25536 2808 25540
rect 2824 25596 2888 25600
rect 2824 25540 2828 25596
rect 2828 25540 2884 25596
rect 2884 25540 2888 25596
rect 2824 25536 2888 25540
rect 5848 25596 5912 25600
rect 5848 25540 5852 25596
rect 5852 25540 5908 25596
rect 5908 25540 5912 25596
rect 5848 25536 5912 25540
rect 5928 25596 5992 25600
rect 5928 25540 5932 25596
rect 5932 25540 5988 25596
rect 5988 25540 5992 25596
rect 5928 25536 5992 25540
rect 6008 25596 6072 25600
rect 6008 25540 6012 25596
rect 6012 25540 6068 25596
rect 6068 25540 6072 25596
rect 6008 25536 6072 25540
rect 6088 25596 6152 25600
rect 6088 25540 6092 25596
rect 6092 25540 6148 25596
rect 6148 25540 6152 25596
rect 6088 25536 6152 25540
rect 9112 25596 9176 25600
rect 9112 25540 9116 25596
rect 9116 25540 9172 25596
rect 9172 25540 9176 25596
rect 9112 25536 9176 25540
rect 9192 25596 9256 25600
rect 9192 25540 9196 25596
rect 9196 25540 9252 25596
rect 9252 25540 9256 25596
rect 9192 25536 9256 25540
rect 9272 25596 9336 25600
rect 9272 25540 9276 25596
rect 9276 25540 9332 25596
rect 9332 25540 9336 25596
rect 9272 25536 9336 25540
rect 9352 25596 9416 25600
rect 9352 25540 9356 25596
rect 9356 25540 9412 25596
rect 9412 25540 9416 25596
rect 9352 25536 9416 25540
rect 3740 25196 3804 25260
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 7480 25052 7544 25056
rect 7480 24996 7484 25052
rect 7484 24996 7540 25052
rect 7540 24996 7544 25052
rect 7480 24992 7544 24996
rect 7560 25052 7624 25056
rect 7560 24996 7564 25052
rect 7564 24996 7620 25052
rect 7620 24996 7624 25052
rect 7560 24992 7624 24996
rect 7640 25052 7704 25056
rect 7640 24996 7644 25052
rect 7644 24996 7700 25052
rect 7700 24996 7704 25052
rect 7640 24992 7704 24996
rect 7720 25052 7784 25056
rect 7720 24996 7724 25052
rect 7724 24996 7780 25052
rect 7780 24996 7784 25052
rect 7720 24992 7784 24996
rect 3188 24788 3252 24852
rect 3924 24516 3988 24580
rect 2584 24508 2648 24512
rect 2584 24452 2588 24508
rect 2588 24452 2644 24508
rect 2644 24452 2648 24508
rect 2584 24448 2648 24452
rect 2664 24508 2728 24512
rect 2664 24452 2668 24508
rect 2668 24452 2724 24508
rect 2724 24452 2728 24508
rect 2664 24448 2728 24452
rect 2744 24508 2808 24512
rect 2744 24452 2748 24508
rect 2748 24452 2804 24508
rect 2804 24452 2808 24508
rect 2744 24448 2808 24452
rect 2824 24508 2888 24512
rect 2824 24452 2828 24508
rect 2828 24452 2884 24508
rect 2884 24452 2888 24508
rect 2824 24448 2888 24452
rect 5848 24508 5912 24512
rect 5848 24452 5852 24508
rect 5852 24452 5908 24508
rect 5908 24452 5912 24508
rect 5848 24448 5912 24452
rect 5928 24508 5992 24512
rect 5928 24452 5932 24508
rect 5932 24452 5988 24508
rect 5988 24452 5992 24508
rect 5928 24448 5992 24452
rect 6008 24508 6072 24512
rect 6008 24452 6012 24508
rect 6012 24452 6068 24508
rect 6068 24452 6072 24508
rect 6008 24448 6072 24452
rect 6088 24508 6152 24512
rect 6088 24452 6092 24508
rect 6092 24452 6148 24508
rect 6148 24452 6152 24508
rect 6088 24448 6152 24452
rect 9112 24508 9176 24512
rect 9112 24452 9116 24508
rect 9116 24452 9172 24508
rect 9172 24452 9176 24508
rect 9112 24448 9176 24452
rect 9192 24508 9256 24512
rect 9192 24452 9196 24508
rect 9196 24452 9252 24508
rect 9252 24452 9256 24508
rect 9192 24448 9256 24452
rect 9272 24508 9336 24512
rect 9272 24452 9276 24508
rect 9276 24452 9332 24508
rect 9332 24452 9336 24508
rect 9272 24448 9336 24452
rect 9352 24508 9416 24512
rect 9352 24452 9356 24508
rect 9356 24452 9412 24508
rect 9412 24452 9416 24508
rect 9352 24448 9416 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 7480 23964 7544 23968
rect 7480 23908 7484 23964
rect 7484 23908 7540 23964
rect 7540 23908 7544 23964
rect 7480 23904 7544 23908
rect 7560 23964 7624 23968
rect 7560 23908 7564 23964
rect 7564 23908 7620 23964
rect 7620 23908 7624 23964
rect 7560 23904 7624 23908
rect 7640 23964 7704 23968
rect 7640 23908 7644 23964
rect 7644 23908 7700 23964
rect 7700 23908 7704 23964
rect 7640 23904 7704 23908
rect 7720 23964 7784 23968
rect 7720 23908 7724 23964
rect 7724 23908 7780 23964
rect 7780 23908 7784 23964
rect 7720 23904 7784 23908
rect 2268 23836 2332 23900
rect 2584 23420 2648 23424
rect 2584 23364 2588 23420
rect 2588 23364 2644 23420
rect 2644 23364 2648 23420
rect 2584 23360 2648 23364
rect 2664 23420 2728 23424
rect 2664 23364 2668 23420
rect 2668 23364 2724 23420
rect 2724 23364 2728 23420
rect 2664 23360 2728 23364
rect 2744 23420 2808 23424
rect 2744 23364 2748 23420
rect 2748 23364 2804 23420
rect 2804 23364 2808 23420
rect 2744 23360 2808 23364
rect 2824 23420 2888 23424
rect 2824 23364 2828 23420
rect 2828 23364 2884 23420
rect 2884 23364 2888 23420
rect 2824 23360 2888 23364
rect 5848 23420 5912 23424
rect 5848 23364 5852 23420
rect 5852 23364 5908 23420
rect 5908 23364 5912 23420
rect 5848 23360 5912 23364
rect 5928 23420 5992 23424
rect 5928 23364 5932 23420
rect 5932 23364 5988 23420
rect 5988 23364 5992 23420
rect 5928 23360 5992 23364
rect 6008 23420 6072 23424
rect 6008 23364 6012 23420
rect 6012 23364 6068 23420
rect 6068 23364 6072 23420
rect 6008 23360 6072 23364
rect 6088 23420 6152 23424
rect 6088 23364 6092 23420
rect 6092 23364 6148 23420
rect 6148 23364 6152 23420
rect 6088 23360 6152 23364
rect 9112 23420 9176 23424
rect 9112 23364 9116 23420
rect 9116 23364 9172 23420
rect 9172 23364 9176 23420
rect 9112 23360 9176 23364
rect 9192 23420 9256 23424
rect 9192 23364 9196 23420
rect 9196 23364 9252 23420
rect 9252 23364 9256 23420
rect 9192 23360 9256 23364
rect 9272 23420 9336 23424
rect 9272 23364 9276 23420
rect 9276 23364 9332 23420
rect 9332 23364 9336 23420
rect 9272 23360 9336 23364
rect 9352 23420 9416 23424
rect 9352 23364 9356 23420
rect 9356 23364 9412 23420
rect 9412 23364 9416 23420
rect 9352 23360 9416 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 7480 22876 7544 22880
rect 7480 22820 7484 22876
rect 7484 22820 7540 22876
rect 7540 22820 7544 22876
rect 7480 22816 7544 22820
rect 7560 22876 7624 22880
rect 7560 22820 7564 22876
rect 7564 22820 7620 22876
rect 7620 22820 7624 22876
rect 7560 22816 7624 22820
rect 7640 22876 7704 22880
rect 7640 22820 7644 22876
rect 7644 22820 7700 22876
rect 7700 22820 7704 22876
rect 7640 22816 7704 22820
rect 7720 22876 7784 22880
rect 7720 22820 7724 22876
rect 7724 22820 7780 22876
rect 7780 22820 7784 22876
rect 7720 22816 7784 22820
rect 3372 22748 3436 22812
rect 2584 22332 2648 22336
rect 2584 22276 2588 22332
rect 2588 22276 2644 22332
rect 2644 22276 2648 22332
rect 2584 22272 2648 22276
rect 2664 22332 2728 22336
rect 2664 22276 2668 22332
rect 2668 22276 2724 22332
rect 2724 22276 2728 22332
rect 2664 22272 2728 22276
rect 2744 22332 2808 22336
rect 2744 22276 2748 22332
rect 2748 22276 2804 22332
rect 2804 22276 2808 22332
rect 2744 22272 2808 22276
rect 2824 22332 2888 22336
rect 2824 22276 2828 22332
rect 2828 22276 2884 22332
rect 2884 22276 2888 22332
rect 2824 22272 2888 22276
rect 5848 22332 5912 22336
rect 5848 22276 5852 22332
rect 5852 22276 5908 22332
rect 5908 22276 5912 22332
rect 5848 22272 5912 22276
rect 5928 22332 5992 22336
rect 5928 22276 5932 22332
rect 5932 22276 5988 22332
rect 5988 22276 5992 22332
rect 5928 22272 5992 22276
rect 6008 22332 6072 22336
rect 6008 22276 6012 22332
rect 6012 22276 6068 22332
rect 6068 22276 6072 22332
rect 6008 22272 6072 22276
rect 6088 22332 6152 22336
rect 6088 22276 6092 22332
rect 6092 22276 6148 22332
rect 6148 22276 6152 22332
rect 6088 22272 6152 22276
rect 9112 22332 9176 22336
rect 9112 22276 9116 22332
rect 9116 22276 9172 22332
rect 9172 22276 9176 22332
rect 9112 22272 9176 22276
rect 9192 22332 9256 22336
rect 9192 22276 9196 22332
rect 9196 22276 9252 22332
rect 9252 22276 9256 22332
rect 9192 22272 9256 22276
rect 9272 22332 9336 22336
rect 9272 22276 9276 22332
rect 9276 22276 9332 22332
rect 9332 22276 9336 22332
rect 9272 22272 9336 22276
rect 9352 22332 9416 22336
rect 9352 22276 9356 22332
rect 9356 22276 9412 22332
rect 9412 22276 9416 22332
rect 9352 22272 9416 22276
rect 2268 22264 2332 22268
rect 2268 22208 2318 22264
rect 2318 22208 2332 22264
rect 2268 22204 2332 22208
rect 3556 22204 3620 22268
rect 2268 21992 2332 21996
rect 2268 21936 2282 21992
rect 2282 21936 2332 21992
rect 2268 21932 2332 21936
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 7480 21788 7544 21792
rect 7480 21732 7484 21788
rect 7484 21732 7540 21788
rect 7540 21732 7544 21788
rect 7480 21728 7544 21732
rect 7560 21788 7624 21792
rect 7560 21732 7564 21788
rect 7564 21732 7620 21788
rect 7620 21732 7624 21788
rect 7560 21728 7624 21732
rect 7640 21788 7704 21792
rect 7640 21732 7644 21788
rect 7644 21732 7700 21788
rect 7700 21732 7704 21788
rect 7640 21728 7704 21732
rect 7720 21788 7784 21792
rect 7720 21732 7724 21788
rect 7724 21732 7780 21788
rect 7780 21732 7784 21788
rect 7720 21728 7784 21732
rect 2584 21244 2648 21248
rect 2584 21188 2588 21244
rect 2588 21188 2644 21244
rect 2644 21188 2648 21244
rect 2584 21184 2648 21188
rect 2664 21244 2728 21248
rect 2664 21188 2668 21244
rect 2668 21188 2724 21244
rect 2724 21188 2728 21244
rect 2664 21184 2728 21188
rect 2744 21244 2808 21248
rect 2744 21188 2748 21244
rect 2748 21188 2804 21244
rect 2804 21188 2808 21244
rect 2744 21184 2808 21188
rect 2824 21244 2888 21248
rect 2824 21188 2828 21244
rect 2828 21188 2884 21244
rect 2884 21188 2888 21244
rect 2824 21184 2888 21188
rect 5848 21244 5912 21248
rect 5848 21188 5852 21244
rect 5852 21188 5908 21244
rect 5908 21188 5912 21244
rect 5848 21184 5912 21188
rect 5928 21244 5992 21248
rect 5928 21188 5932 21244
rect 5932 21188 5988 21244
rect 5988 21188 5992 21244
rect 5928 21184 5992 21188
rect 6008 21244 6072 21248
rect 6008 21188 6012 21244
rect 6012 21188 6068 21244
rect 6068 21188 6072 21244
rect 6008 21184 6072 21188
rect 6088 21244 6152 21248
rect 6088 21188 6092 21244
rect 6092 21188 6148 21244
rect 6148 21188 6152 21244
rect 6088 21184 6152 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 9272 21244 9336 21248
rect 9272 21188 9276 21244
rect 9276 21188 9332 21244
rect 9332 21188 9336 21244
rect 9272 21184 9336 21188
rect 9352 21244 9416 21248
rect 9352 21188 9356 21244
rect 9356 21188 9412 21244
rect 9412 21188 9416 21244
rect 9352 21184 9416 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 7480 20700 7544 20704
rect 7480 20644 7484 20700
rect 7484 20644 7540 20700
rect 7540 20644 7544 20700
rect 7480 20640 7544 20644
rect 7560 20700 7624 20704
rect 7560 20644 7564 20700
rect 7564 20644 7620 20700
rect 7620 20644 7624 20700
rect 7560 20640 7624 20644
rect 7640 20700 7704 20704
rect 7640 20644 7644 20700
rect 7644 20644 7700 20700
rect 7700 20644 7704 20700
rect 7640 20640 7704 20644
rect 7720 20700 7784 20704
rect 7720 20644 7724 20700
rect 7724 20644 7780 20700
rect 7780 20644 7784 20700
rect 7720 20640 7784 20644
rect 2584 20156 2648 20160
rect 2584 20100 2588 20156
rect 2588 20100 2644 20156
rect 2644 20100 2648 20156
rect 2584 20096 2648 20100
rect 2664 20156 2728 20160
rect 2664 20100 2668 20156
rect 2668 20100 2724 20156
rect 2724 20100 2728 20156
rect 2664 20096 2728 20100
rect 2744 20156 2808 20160
rect 2744 20100 2748 20156
rect 2748 20100 2804 20156
rect 2804 20100 2808 20156
rect 2744 20096 2808 20100
rect 2824 20156 2888 20160
rect 2824 20100 2828 20156
rect 2828 20100 2884 20156
rect 2884 20100 2888 20156
rect 2824 20096 2888 20100
rect 5848 20156 5912 20160
rect 5848 20100 5852 20156
rect 5852 20100 5908 20156
rect 5908 20100 5912 20156
rect 5848 20096 5912 20100
rect 5928 20156 5992 20160
rect 5928 20100 5932 20156
rect 5932 20100 5988 20156
rect 5988 20100 5992 20156
rect 5928 20096 5992 20100
rect 6008 20156 6072 20160
rect 6008 20100 6012 20156
rect 6012 20100 6068 20156
rect 6068 20100 6072 20156
rect 6008 20096 6072 20100
rect 6088 20156 6152 20160
rect 6088 20100 6092 20156
rect 6092 20100 6148 20156
rect 6148 20100 6152 20156
rect 6088 20096 6152 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 9272 20156 9336 20160
rect 9272 20100 9276 20156
rect 9276 20100 9332 20156
rect 9332 20100 9336 20156
rect 9272 20096 9336 20100
rect 9352 20156 9416 20160
rect 9352 20100 9356 20156
rect 9356 20100 9412 20156
rect 9412 20100 9416 20156
rect 9352 20096 9416 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 7480 19612 7544 19616
rect 7480 19556 7484 19612
rect 7484 19556 7540 19612
rect 7540 19556 7544 19612
rect 7480 19552 7544 19556
rect 7560 19612 7624 19616
rect 7560 19556 7564 19612
rect 7564 19556 7620 19612
rect 7620 19556 7624 19612
rect 7560 19552 7624 19556
rect 7640 19612 7704 19616
rect 7640 19556 7644 19612
rect 7644 19556 7700 19612
rect 7700 19556 7704 19612
rect 7640 19552 7704 19556
rect 7720 19612 7784 19616
rect 7720 19556 7724 19612
rect 7724 19556 7780 19612
rect 7780 19556 7784 19612
rect 7720 19552 7784 19556
rect 2584 19068 2648 19072
rect 2584 19012 2588 19068
rect 2588 19012 2644 19068
rect 2644 19012 2648 19068
rect 2584 19008 2648 19012
rect 2664 19068 2728 19072
rect 2664 19012 2668 19068
rect 2668 19012 2724 19068
rect 2724 19012 2728 19068
rect 2664 19008 2728 19012
rect 2744 19068 2808 19072
rect 2744 19012 2748 19068
rect 2748 19012 2804 19068
rect 2804 19012 2808 19068
rect 2744 19008 2808 19012
rect 2824 19068 2888 19072
rect 2824 19012 2828 19068
rect 2828 19012 2884 19068
rect 2884 19012 2888 19068
rect 2824 19008 2888 19012
rect 5848 19068 5912 19072
rect 5848 19012 5852 19068
rect 5852 19012 5908 19068
rect 5908 19012 5912 19068
rect 5848 19008 5912 19012
rect 5928 19068 5992 19072
rect 5928 19012 5932 19068
rect 5932 19012 5988 19068
rect 5988 19012 5992 19068
rect 5928 19008 5992 19012
rect 6008 19068 6072 19072
rect 6008 19012 6012 19068
rect 6012 19012 6068 19068
rect 6068 19012 6072 19068
rect 6008 19008 6072 19012
rect 6088 19068 6152 19072
rect 6088 19012 6092 19068
rect 6092 19012 6148 19068
rect 6148 19012 6152 19068
rect 6088 19008 6152 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 9272 19068 9336 19072
rect 9272 19012 9276 19068
rect 9276 19012 9332 19068
rect 9332 19012 9336 19068
rect 9272 19008 9336 19012
rect 9352 19068 9416 19072
rect 9352 19012 9356 19068
rect 9356 19012 9412 19068
rect 9412 19012 9416 19068
rect 9352 19008 9416 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 7480 18524 7544 18528
rect 7480 18468 7484 18524
rect 7484 18468 7540 18524
rect 7540 18468 7544 18524
rect 7480 18464 7544 18468
rect 7560 18524 7624 18528
rect 7560 18468 7564 18524
rect 7564 18468 7620 18524
rect 7620 18468 7624 18524
rect 7560 18464 7624 18468
rect 7640 18524 7704 18528
rect 7640 18468 7644 18524
rect 7644 18468 7700 18524
rect 7700 18468 7704 18524
rect 7640 18464 7704 18468
rect 7720 18524 7784 18528
rect 7720 18468 7724 18524
rect 7724 18468 7780 18524
rect 7780 18468 7784 18524
rect 7720 18464 7784 18468
rect 2584 17980 2648 17984
rect 2584 17924 2588 17980
rect 2588 17924 2644 17980
rect 2644 17924 2648 17980
rect 2584 17920 2648 17924
rect 2664 17980 2728 17984
rect 2664 17924 2668 17980
rect 2668 17924 2724 17980
rect 2724 17924 2728 17980
rect 2664 17920 2728 17924
rect 2744 17980 2808 17984
rect 2744 17924 2748 17980
rect 2748 17924 2804 17980
rect 2804 17924 2808 17980
rect 2744 17920 2808 17924
rect 2824 17980 2888 17984
rect 2824 17924 2828 17980
rect 2828 17924 2884 17980
rect 2884 17924 2888 17980
rect 2824 17920 2888 17924
rect 5848 17980 5912 17984
rect 5848 17924 5852 17980
rect 5852 17924 5908 17980
rect 5908 17924 5912 17980
rect 5848 17920 5912 17924
rect 5928 17980 5992 17984
rect 5928 17924 5932 17980
rect 5932 17924 5988 17980
rect 5988 17924 5992 17980
rect 5928 17920 5992 17924
rect 6008 17980 6072 17984
rect 6008 17924 6012 17980
rect 6012 17924 6068 17980
rect 6068 17924 6072 17980
rect 6008 17920 6072 17924
rect 6088 17980 6152 17984
rect 6088 17924 6092 17980
rect 6092 17924 6148 17980
rect 6148 17924 6152 17980
rect 6088 17920 6152 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 9272 17980 9336 17984
rect 9272 17924 9276 17980
rect 9276 17924 9332 17980
rect 9332 17924 9336 17980
rect 9272 17920 9336 17924
rect 9352 17980 9416 17984
rect 9352 17924 9356 17980
rect 9356 17924 9412 17980
rect 9412 17924 9416 17980
rect 9352 17920 9416 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 7480 17436 7544 17440
rect 7480 17380 7484 17436
rect 7484 17380 7540 17436
rect 7540 17380 7544 17436
rect 7480 17376 7544 17380
rect 7560 17436 7624 17440
rect 7560 17380 7564 17436
rect 7564 17380 7620 17436
rect 7620 17380 7624 17436
rect 7560 17376 7624 17380
rect 7640 17436 7704 17440
rect 7640 17380 7644 17436
rect 7644 17380 7700 17436
rect 7700 17380 7704 17436
rect 7640 17376 7704 17380
rect 7720 17436 7784 17440
rect 7720 17380 7724 17436
rect 7724 17380 7780 17436
rect 7780 17380 7784 17436
rect 7720 17376 7784 17380
rect 2584 16892 2648 16896
rect 2584 16836 2588 16892
rect 2588 16836 2644 16892
rect 2644 16836 2648 16892
rect 2584 16832 2648 16836
rect 2664 16892 2728 16896
rect 2664 16836 2668 16892
rect 2668 16836 2724 16892
rect 2724 16836 2728 16892
rect 2664 16832 2728 16836
rect 2744 16892 2808 16896
rect 2744 16836 2748 16892
rect 2748 16836 2804 16892
rect 2804 16836 2808 16892
rect 2744 16832 2808 16836
rect 2824 16892 2888 16896
rect 2824 16836 2828 16892
rect 2828 16836 2884 16892
rect 2884 16836 2888 16892
rect 2824 16832 2888 16836
rect 5848 16892 5912 16896
rect 5848 16836 5852 16892
rect 5852 16836 5908 16892
rect 5908 16836 5912 16892
rect 5848 16832 5912 16836
rect 5928 16892 5992 16896
rect 5928 16836 5932 16892
rect 5932 16836 5988 16892
rect 5988 16836 5992 16892
rect 5928 16832 5992 16836
rect 6008 16892 6072 16896
rect 6008 16836 6012 16892
rect 6012 16836 6068 16892
rect 6068 16836 6072 16892
rect 6008 16832 6072 16836
rect 6088 16892 6152 16896
rect 6088 16836 6092 16892
rect 6092 16836 6148 16892
rect 6148 16836 6152 16892
rect 6088 16832 6152 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 9272 16892 9336 16896
rect 9272 16836 9276 16892
rect 9276 16836 9332 16892
rect 9332 16836 9336 16892
rect 9272 16832 9336 16836
rect 9352 16892 9416 16896
rect 9352 16836 9356 16892
rect 9356 16836 9412 16892
rect 9412 16836 9416 16892
rect 9352 16832 9416 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 7480 16348 7544 16352
rect 7480 16292 7484 16348
rect 7484 16292 7540 16348
rect 7540 16292 7544 16348
rect 7480 16288 7544 16292
rect 7560 16348 7624 16352
rect 7560 16292 7564 16348
rect 7564 16292 7620 16348
rect 7620 16292 7624 16348
rect 7560 16288 7624 16292
rect 7640 16348 7704 16352
rect 7640 16292 7644 16348
rect 7644 16292 7700 16348
rect 7700 16292 7704 16348
rect 7640 16288 7704 16292
rect 7720 16348 7784 16352
rect 7720 16292 7724 16348
rect 7724 16292 7780 16348
rect 7780 16292 7784 16348
rect 7720 16288 7784 16292
rect 2584 15804 2648 15808
rect 2584 15748 2588 15804
rect 2588 15748 2644 15804
rect 2644 15748 2648 15804
rect 2584 15744 2648 15748
rect 2664 15804 2728 15808
rect 2664 15748 2668 15804
rect 2668 15748 2724 15804
rect 2724 15748 2728 15804
rect 2664 15744 2728 15748
rect 2744 15804 2808 15808
rect 2744 15748 2748 15804
rect 2748 15748 2804 15804
rect 2804 15748 2808 15804
rect 2744 15744 2808 15748
rect 2824 15804 2888 15808
rect 2824 15748 2828 15804
rect 2828 15748 2884 15804
rect 2884 15748 2888 15804
rect 2824 15744 2888 15748
rect 5848 15804 5912 15808
rect 5848 15748 5852 15804
rect 5852 15748 5908 15804
rect 5908 15748 5912 15804
rect 5848 15744 5912 15748
rect 5928 15804 5992 15808
rect 5928 15748 5932 15804
rect 5932 15748 5988 15804
rect 5988 15748 5992 15804
rect 5928 15744 5992 15748
rect 6008 15804 6072 15808
rect 6008 15748 6012 15804
rect 6012 15748 6068 15804
rect 6068 15748 6072 15804
rect 6008 15744 6072 15748
rect 6088 15804 6152 15808
rect 6088 15748 6092 15804
rect 6092 15748 6148 15804
rect 6148 15748 6152 15804
rect 6088 15744 6152 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 9272 15804 9336 15808
rect 9272 15748 9276 15804
rect 9276 15748 9332 15804
rect 9332 15748 9336 15804
rect 9272 15744 9336 15748
rect 9352 15804 9416 15808
rect 9352 15748 9356 15804
rect 9356 15748 9412 15804
rect 9412 15748 9416 15804
rect 9352 15744 9416 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 7480 15260 7544 15264
rect 7480 15204 7484 15260
rect 7484 15204 7540 15260
rect 7540 15204 7544 15260
rect 7480 15200 7544 15204
rect 7560 15260 7624 15264
rect 7560 15204 7564 15260
rect 7564 15204 7620 15260
rect 7620 15204 7624 15260
rect 7560 15200 7624 15204
rect 7640 15260 7704 15264
rect 7640 15204 7644 15260
rect 7644 15204 7700 15260
rect 7700 15204 7704 15260
rect 7640 15200 7704 15204
rect 7720 15260 7784 15264
rect 7720 15204 7724 15260
rect 7724 15204 7780 15260
rect 7780 15204 7784 15260
rect 7720 15200 7784 15204
rect 5580 14996 5644 15060
rect 2584 14716 2648 14720
rect 2584 14660 2588 14716
rect 2588 14660 2644 14716
rect 2644 14660 2648 14716
rect 2584 14656 2648 14660
rect 2664 14716 2728 14720
rect 2664 14660 2668 14716
rect 2668 14660 2724 14716
rect 2724 14660 2728 14716
rect 2664 14656 2728 14660
rect 2744 14716 2808 14720
rect 2744 14660 2748 14716
rect 2748 14660 2804 14716
rect 2804 14660 2808 14716
rect 2744 14656 2808 14660
rect 2824 14716 2888 14720
rect 2824 14660 2828 14716
rect 2828 14660 2884 14716
rect 2884 14660 2888 14716
rect 2824 14656 2888 14660
rect 5848 14716 5912 14720
rect 5848 14660 5852 14716
rect 5852 14660 5908 14716
rect 5908 14660 5912 14716
rect 5848 14656 5912 14660
rect 5928 14716 5992 14720
rect 5928 14660 5932 14716
rect 5932 14660 5988 14716
rect 5988 14660 5992 14716
rect 5928 14656 5992 14660
rect 6008 14716 6072 14720
rect 6008 14660 6012 14716
rect 6012 14660 6068 14716
rect 6068 14660 6072 14716
rect 6008 14656 6072 14660
rect 6088 14716 6152 14720
rect 6088 14660 6092 14716
rect 6092 14660 6148 14716
rect 6148 14660 6152 14716
rect 6088 14656 6152 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 9272 14716 9336 14720
rect 9272 14660 9276 14716
rect 9276 14660 9332 14716
rect 9332 14660 9336 14716
rect 9272 14656 9336 14660
rect 9352 14716 9416 14720
rect 9352 14660 9356 14716
rect 9356 14660 9412 14716
rect 9412 14660 9416 14716
rect 9352 14656 9416 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 7480 14172 7544 14176
rect 7480 14116 7484 14172
rect 7484 14116 7540 14172
rect 7540 14116 7544 14172
rect 7480 14112 7544 14116
rect 7560 14172 7624 14176
rect 7560 14116 7564 14172
rect 7564 14116 7620 14172
rect 7620 14116 7624 14172
rect 7560 14112 7624 14116
rect 7640 14172 7704 14176
rect 7640 14116 7644 14172
rect 7644 14116 7700 14172
rect 7700 14116 7704 14172
rect 7640 14112 7704 14116
rect 7720 14172 7784 14176
rect 7720 14116 7724 14172
rect 7724 14116 7780 14172
rect 7780 14116 7784 14172
rect 7720 14112 7784 14116
rect 2584 13628 2648 13632
rect 2584 13572 2588 13628
rect 2588 13572 2644 13628
rect 2644 13572 2648 13628
rect 2584 13568 2648 13572
rect 2664 13628 2728 13632
rect 2664 13572 2668 13628
rect 2668 13572 2724 13628
rect 2724 13572 2728 13628
rect 2664 13568 2728 13572
rect 2744 13628 2808 13632
rect 2744 13572 2748 13628
rect 2748 13572 2804 13628
rect 2804 13572 2808 13628
rect 2744 13568 2808 13572
rect 2824 13628 2888 13632
rect 2824 13572 2828 13628
rect 2828 13572 2884 13628
rect 2884 13572 2888 13628
rect 2824 13568 2888 13572
rect 5848 13628 5912 13632
rect 5848 13572 5852 13628
rect 5852 13572 5908 13628
rect 5908 13572 5912 13628
rect 5848 13568 5912 13572
rect 5928 13628 5992 13632
rect 5928 13572 5932 13628
rect 5932 13572 5988 13628
rect 5988 13572 5992 13628
rect 5928 13568 5992 13572
rect 6008 13628 6072 13632
rect 6008 13572 6012 13628
rect 6012 13572 6068 13628
rect 6068 13572 6072 13628
rect 6008 13568 6072 13572
rect 6088 13628 6152 13632
rect 6088 13572 6092 13628
rect 6092 13572 6148 13628
rect 6148 13572 6152 13628
rect 6088 13568 6152 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 9272 13628 9336 13632
rect 9272 13572 9276 13628
rect 9276 13572 9332 13628
rect 9332 13572 9336 13628
rect 9272 13568 9336 13572
rect 9352 13628 9416 13632
rect 9352 13572 9356 13628
rect 9356 13572 9412 13628
rect 9412 13572 9416 13628
rect 9352 13568 9416 13572
rect 1900 13092 1964 13156
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 7480 13084 7544 13088
rect 7480 13028 7484 13084
rect 7484 13028 7540 13084
rect 7540 13028 7544 13084
rect 7480 13024 7544 13028
rect 7560 13084 7624 13088
rect 7560 13028 7564 13084
rect 7564 13028 7620 13084
rect 7620 13028 7624 13084
rect 7560 13024 7624 13028
rect 7640 13084 7704 13088
rect 7640 13028 7644 13084
rect 7644 13028 7700 13084
rect 7700 13028 7704 13084
rect 7640 13024 7704 13028
rect 7720 13084 7784 13088
rect 7720 13028 7724 13084
rect 7724 13028 7780 13084
rect 7780 13028 7784 13084
rect 7720 13024 7784 13028
rect 2584 12540 2648 12544
rect 2584 12484 2588 12540
rect 2588 12484 2644 12540
rect 2644 12484 2648 12540
rect 2584 12480 2648 12484
rect 2664 12540 2728 12544
rect 2664 12484 2668 12540
rect 2668 12484 2724 12540
rect 2724 12484 2728 12540
rect 2664 12480 2728 12484
rect 2744 12540 2808 12544
rect 2744 12484 2748 12540
rect 2748 12484 2804 12540
rect 2804 12484 2808 12540
rect 2744 12480 2808 12484
rect 2824 12540 2888 12544
rect 2824 12484 2828 12540
rect 2828 12484 2884 12540
rect 2884 12484 2888 12540
rect 2824 12480 2888 12484
rect 5848 12540 5912 12544
rect 5848 12484 5852 12540
rect 5852 12484 5908 12540
rect 5908 12484 5912 12540
rect 5848 12480 5912 12484
rect 5928 12540 5992 12544
rect 5928 12484 5932 12540
rect 5932 12484 5988 12540
rect 5988 12484 5992 12540
rect 5928 12480 5992 12484
rect 6008 12540 6072 12544
rect 6008 12484 6012 12540
rect 6012 12484 6068 12540
rect 6068 12484 6072 12540
rect 6008 12480 6072 12484
rect 6088 12540 6152 12544
rect 6088 12484 6092 12540
rect 6092 12484 6148 12540
rect 6148 12484 6152 12540
rect 6088 12480 6152 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 9272 12540 9336 12544
rect 9272 12484 9276 12540
rect 9276 12484 9332 12540
rect 9332 12484 9336 12540
rect 9272 12480 9336 12484
rect 9352 12540 9416 12544
rect 9352 12484 9356 12540
rect 9356 12484 9412 12540
rect 9412 12484 9416 12540
rect 9352 12480 9416 12484
rect 1900 12412 1964 12476
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 7480 11996 7544 12000
rect 7480 11940 7484 11996
rect 7484 11940 7540 11996
rect 7540 11940 7544 11996
rect 7480 11936 7544 11940
rect 7560 11996 7624 12000
rect 7560 11940 7564 11996
rect 7564 11940 7620 11996
rect 7620 11940 7624 11996
rect 7560 11936 7624 11940
rect 7640 11996 7704 12000
rect 7640 11940 7644 11996
rect 7644 11940 7700 11996
rect 7700 11940 7704 11996
rect 7640 11936 7704 11940
rect 7720 11996 7784 12000
rect 7720 11940 7724 11996
rect 7724 11940 7780 11996
rect 7780 11940 7784 11996
rect 7720 11936 7784 11940
rect 2584 11452 2648 11456
rect 2584 11396 2588 11452
rect 2588 11396 2644 11452
rect 2644 11396 2648 11452
rect 2584 11392 2648 11396
rect 2664 11452 2728 11456
rect 2664 11396 2668 11452
rect 2668 11396 2724 11452
rect 2724 11396 2728 11452
rect 2664 11392 2728 11396
rect 2744 11452 2808 11456
rect 2744 11396 2748 11452
rect 2748 11396 2804 11452
rect 2804 11396 2808 11452
rect 2744 11392 2808 11396
rect 2824 11452 2888 11456
rect 2824 11396 2828 11452
rect 2828 11396 2884 11452
rect 2884 11396 2888 11452
rect 2824 11392 2888 11396
rect 5848 11452 5912 11456
rect 5848 11396 5852 11452
rect 5852 11396 5908 11452
rect 5908 11396 5912 11452
rect 5848 11392 5912 11396
rect 5928 11452 5992 11456
rect 5928 11396 5932 11452
rect 5932 11396 5988 11452
rect 5988 11396 5992 11452
rect 5928 11392 5992 11396
rect 6008 11452 6072 11456
rect 6008 11396 6012 11452
rect 6012 11396 6068 11452
rect 6068 11396 6072 11452
rect 6008 11392 6072 11396
rect 6088 11452 6152 11456
rect 6088 11396 6092 11452
rect 6092 11396 6148 11452
rect 6148 11396 6152 11452
rect 6088 11392 6152 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 9272 11452 9336 11456
rect 9272 11396 9276 11452
rect 9276 11396 9332 11452
rect 9332 11396 9336 11452
rect 9272 11392 9336 11396
rect 9352 11452 9416 11456
rect 9352 11396 9356 11452
rect 9356 11396 9412 11452
rect 9412 11396 9416 11452
rect 9352 11392 9416 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 7480 10908 7544 10912
rect 7480 10852 7484 10908
rect 7484 10852 7540 10908
rect 7540 10852 7544 10908
rect 7480 10848 7544 10852
rect 7560 10908 7624 10912
rect 7560 10852 7564 10908
rect 7564 10852 7620 10908
rect 7620 10852 7624 10908
rect 7560 10848 7624 10852
rect 7640 10908 7704 10912
rect 7640 10852 7644 10908
rect 7644 10852 7700 10908
rect 7700 10852 7704 10908
rect 7640 10848 7704 10852
rect 7720 10908 7784 10912
rect 7720 10852 7724 10908
rect 7724 10852 7780 10908
rect 7780 10852 7784 10908
rect 7720 10848 7784 10852
rect 2584 10364 2648 10368
rect 2584 10308 2588 10364
rect 2588 10308 2644 10364
rect 2644 10308 2648 10364
rect 2584 10304 2648 10308
rect 2664 10364 2728 10368
rect 2664 10308 2668 10364
rect 2668 10308 2724 10364
rect 2724 10308 2728 10364
rect 2664 10304 2728 10308
rect 2744 10364 2808 10368
rect 2744 10308 2748 10364
rect 2748 10308 2804 10364
rect 2804 10308 2808 10364
rect 2744 10304 2808 10308
rect 2824 10364 2888 10368
rect 2824 10308 2828 10364
rect 2828 10308 2884 10364
rect 2884 10308 2888 10364
rect 2824 10304 2888 10308
rect 5848 10364 5912 10368
rect 5848 10308 5852 10364
rect 5852 10308 5908 10364
rect 5908 10308 5912 10364
rect 5848 10304 5912 10308
rect 5928 10364 5992 10368
rect 5928 10308 5932 10364
rect 5932 10308 5988 10364
rect 5988 10308 5992 10364
rect 5928 10304 5992 10308
rect 6008 10364 6072 10368
rect 6008 10308 6012 10364
rect 6012 10308 6068 10364
rect 6068 10308 6072 10364
rect 6008 10304 6072 10308
rect 6088 10364 6152 10368
rect 6088 10308 6092 10364
rect 6092 10308 6148 10364
rect 6148 10308 6152 10364
rect 6088 10304 6152 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 9272 10364 9336 10368
rect 9272 10308 9276 10364
rect 9276 10308 9332 10364
rect 9332 10308 9336 10364
rect 9272 10304 9336 10308
rect 9352 10364 9416 10368
rect 9352 10308 9356 10364
rect 9356 10308 9412 10364
rect 9412 10308 9416 10364
rect 9352 10304 9416 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 7480 9820 7544 9824
rect 7480 9764 7484 9820
rect 7484 9764 7540 9820
rect 7540 9764 7544 9820
rect 7480 9760 7544 9764
rect 7560 9820 7624 9824
rect 7560 9764 7564 9820
rect 7564 9764 7620 9820
rect 7620 9764 7624 9820
rect 7560 9760 7624 9764
rect 7640 9820 7704 9824
rect 7640 9764 7644 9820
rect 7644 9764 7700 9820
rect 7700 9764 7704 9820
rect 7640 9760 7704 9764
rect 7720 9820 7784 9824
rect 7720 9764 7724 9820
rect 7724 9764 7780 9820
rect 7780 9764 7784 9820
rect 7720 9760 7784 9764
rect 4844 9420 4908 9484
rect 2584 9276 2648 9280
rect 2584 9220 2588 9276
rect 2588 9220 2644 9276
rect 2644 9220 2648 9276
rect 2584 9216 2648 9220
rect 2664 9276 2728 9280
rect 2664 9220 2668 9276
rect 2668 9220 2724 9276
rect 2724 9220 2728 9276
rect 2664 9216 2728 9220
rect 2744 9276 2808 9280
rect 2744 9220 2748 9276
rect 2748 9220 2804 9276
rect 2804 9220 2808 9276
rect 2744 9216 2808 9220
rect 2824 9276 2888 9280
rect 2824 9220 2828 9276
rect 2828 9220 2884 9276
rect 2884 9220 2888 9276
rect 2824 9216 2888 9220
rect 5848 9276 5912 9280
rect 5848 9220 5852 9276
rect 5852 9220 5908 9276
rect 5908 9220 5912 9276
rect 5848 9216 5912 9220
rect 5928 9276 5992 9280
rect 5928 9220 5932 9276
rect 5932 9220 5988 9276
rect 5988 9220 5992 9276
rect 5928 9216 5992 9220
rect 6008 9276 6072 9280
rect 6008 9220 6012 9276
rect 6012 9220 6068 9276
rect 6068 9220 6072 9276
rect 6008 9216 6072 9220
rect 6088 9276 6152 9280
rect 6088 9220 6092 9276
rect 6092 9220 6148 9276
rect 6148 9220 6152 9276
rect 6088 9216 6152 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 9272 9276 9336 9280
rect 9272 9220 9276 9276
rect 9276 9220 9332 9276
rect 9332 9220 9336 9276
rect 9272 9216 9336 9220
rect 9352 9276 9416 9280
rect 9352 9220 9356 9276
rect 9356 9220 9412 9276
rect 9412 9220 9416 9276
rect 9352 9216 9416 9220
rect 3004 9208 3068 9212
rect 3004 9152 3018 9208
rect 3018 9152 3068 9208
rect 3004 9148 3068 9152
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 7480 8732 7544 8736
rect 7480 8676 7484 8732
rect 7484 8676 7540 8732
rect 7540 8676 7544 8732
rect 7480 8672 7544 8676
rect 7560 8732 7624 8736
rect 7560 8676 7564 8732
rect 7564 8676 7620 8732
rect 7620 8676 7624 8732
rect 7560 8672 7624 8676
rect 7640 8732 7704 8736
rect 7640 8676 7644 8732
rect 7644 8676 7700 8732
rect 7700 8676 7704 8732
rect 7640 8672 7704 8676
rect 7720 8732 7784 8736
rect 7720 8676 7724 8732
rect 7724 8676 7780 8732
rect 7780 8676 7784 8732
rect 7720 8672 7784 8676
rect 2584 8188 2648 8192
rect 2584 8132 2588 8188
rect 2588 8132 2644 8188
rect 2644 8132 2648 8188
rect 2584 8128 2648 8132
rect 2664 8188 2728 8192
rect 2664 8132 2668 8188
rect 2668 8132 2724 8188
rect 2724 8132 2728 8188
rect 2664 8128 2728 8132
rect 2744 8188 2808 8192
rect 2744 8132 2748 8188
rect 2748 8132 2804 8188
rect 2804 8132 2808 8188
rect 2744 8128 2808 8132
rect 2824 8188 2888 8192
rect 2824 8132 2828 8188
rect 2828 8132 2884 8188
rect 2884 8132 2888 8188
rect 2824 8128 2888 8132
rect 5848 8188 5912 8192
rect 5848 8132 5852 8188
rect 5852 8132 5908 8188
rect 5908 8132 5912 8188
rect 5848 8128 5912 8132
rect 5928 8188 5992 8192
rect 5928 8132 5932 8188
rect 5932 8132 5988 8188
rect 5988 8132 5992 8188
rect 5928 8128 5992 8132
rect 6008 8188 6072 8192
rect 6008 8132 6012 8188
rect 6012 8132 6068 8188
rect 6068 8132 6072 8188
rect 6008 8128 6072 8132
rect 6088 8188 6152 8192
rect 6088 8132 6092 8188
rect 6092 8132 6148 8188
rect 6148 8132 6152 8188
rect 6088 8128 6152 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 9272 8188 9336 8192
rect 9272 8132 9276 8188
rect 9276 8132 9332 8188
rect 9332 8132 9336 8188
rect 9272 8128 9336 8132
rect 9352 8188 9416 8192
rect 9352 8132 9356 8188
rect 9356 8132 9412 8188
rect 9412 8132 9416 8188
rect 9352 8128 9416 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 7480 7644 7544 7648
rect 7480 7588 7484 7644
rect 7484 7588 7540 7644
rect 7540 7588 7544 7644
rect 7480 7584 7544 7588
rect 7560 7644 7624 7648
rect 7560 7588 7564 7644
rect 7564 7588 7620 7644
rect 7620 7588 7624 7644
rect 7560 7584 7624 7588
rect 7640 7644 7704 7648
rect 7640 7588 7644 7644
rect 7644 7588 7700 7644
rect 7700 7588 7704 7644
rect 7640 7584 7704 7588
rect 7720 7644 7784 7648
rect 7720 7588 7724 7644
rect 7724 7588 7780 7644
rect 7780 7588 7784 7644
rect 7720 7584 7784 7588
rect 2584 7100 2648 7104
rect 2584 7044 2588 7100
rect 2588 7044 2644 7100
rect 2644 7044 2648 7100
rect 2584 7040 2648 7044
rect 2664 7100 2728 7104
rect 2664 7044 2668 7100
rect 2668 7044 2724 7100
rect 2724 7044 2728 7100
rect 2664 7040 2728 7044
rect 2744 7100 2808 7104
rect 2744 7044 2748 7100
rect 2748 7044 2804 7100
rect 2804 7044 2808 7100
rect 2744 7040 2808 7044
rect 2824 7100 2888 7104
rect 2824 7044 2828 7100
rect 2828 7044 2884 7100
rect 2884 7044 2888 7100
rect 2824 7040 2888 7044
rect 5848 7100 5912 7104
rect 5848 7044 5852 7100
rect 5852 7044 5908 7100
rect 5908 7044 5912 7100
rect 5848 7040 5912 7044
rect 5928 7100 5992 7104
rect 5928 7044 5932 7100
rect 5932 7044 5988 7100
rect 5988 7044 5992 7100
rect 5928 7040 5992 7044
rect 6008 7100 6072 7104
rect 6008 7044 6012 7100
rect 6012 7044 6068 7100
rect 6068 7044 6072 7100
rect 6008 7040 6072 7044
rect 6088 7100 6152 7104
rect 6088 7044 6092 7100
rect 6092 7044 6148 7100
rect 6148 7044 6152 7100
rect 6088 7040 6152 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 9272 7100 9336 7104
rect 9272 7044 9276 7100
rect 9276 7044 9332 7100
rect 9332 7044 9336 7100
rect 9272 7040 9336 7044
rect 9352 7100 9416 7104
rect 9352 7044 9356 7100
rect 9356 7044 9412 7100
rect 9412 7044 9416 7100
rect 9352 7040 9416 7044
rect 980 6700 1044 6764
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 7480 6556 7544 6560
rect 7480 6500 7484 6556
rect 7484 6500 7540 6556
rect 7540 6500 7544 6556
rect 7480 6496 7544 6500
rect 7560 6556 7624 6560
rect 7560 6500 7564 6556
rect 7564 6500 7620 6556
rect 7620 6500 7624 6556
rect 7560 6496 7624 6500
rect 7640 6556 7704 6560
rect 7640 6500 7644 6556
rect 7644 6500 7700 6556
rect 7700 6500 7704 6556
rect 7640 6496 7704 6500
rect 7720 6556 7784 6560
rect 7720 6500 7724 6556
rect 7724 6500 7780 6556
rect 7780 6500 7784 6556
rect 7720 6496 7784 6500
rect 2584 6012 2648 6016
rect 2584 5956 2588 6012
rect 2588 5956 2644 6012
rect 2644 5956 2648 6012
rect 2584 5952 2648 5956
rect 2664 6012 2728 6016
rect 2664 5956 2668 6012
rect 2668 5956 2724 6012
rect 2724 5956 2728 6012
rect 2664 5952 2728 5956
rect 2744 6012 2808 6016
rect 2744 5956 2748 6012
rect 2748 5956 2804 6012
rect 2804 5956 2808 6012
rect 2744 5952 2808 5956
rect 2824 6012 2888 6016
rect 2824 5956 2828 6012
rect 2828 5956 2884 6012
rect 2884 5956 2888 6012
rect 2824 5952 2888 5956
rect 5848 6012 5912 6016
rect 5848 5956 5852 6012
rect 5852 5956 5908 6012
rect 5908 5956 5912 6012
rect 5848 5952 5912 5956
rect 5928 6012 5992 6016
rect 5928 5956 5932 6012
rect 5932 5956 5988 6012
rect 5988 5956 5992 6012
rect 5928 5952 5992 5956
rect 6008 6012 6072 6016
rect 6008 5956 6012 6012
rect 6012 5956 6068 6012
rect 6068 5956 6072 6012
rect 6008 5952 6072 5956
rect 6088 6012 6152 6016
rect 6088 5956 6092 6012
rect 6092 5956 6148 6012
rect 6148 5956 6152 6012
rect 6088 5952 6152 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 9272 6012 9336 6016
rect 9272 5956 9276 6012
rect 9276 5956 9332 6012
rect 9332 5956 9336 6012
rect 9272 5952 9336 5956
rect 9352 6012 9416 6016
rect 9352 5956 9356 6012
rect 9356 5956 9412 6012
rect 9412 5956 9416 6012
rect 9352 5952 9416 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 7480 5468 7544 5472
rect 7480 5412 7484 5468
rect 7484 5412 7540 5468
rect 7540 5412 7544 5468
rect 7480 5408 7544 5412
rect 7560 5468 7624 5472
rect 7560 5412 7564 5468
rect 7564 5412 7620 5468
rect 7620 5412 7624 5468
rect 7560 5408 7624 5412
rect 7640 5468 7704 5472
rect 7640 5412 7644 5468
rect 7644 5412 7700 5468
rect 7700 5412 7704 5468
rect 7640 5408 7704 5412
rect 7720 5468 7784 5472
rect 7720 5412 7724 5468
rect 7724 5412 7780 5468
rect 7780 5412 7784 5468
rect 7720 5408 7784 5412
rect 8340 5204 8404 5268
rect 2584 4924 2648 4928
rect 2584 4868 2588 4924
rect 2588 4868 2644 4924
rect 2644 4868 2648 4924
rect 2584 4864 2648 4868
rect 2664 4924 2728 4928
rect 2664 4868 2668 4924
rect 2668 4868 2724 4924
rect 2724 4868 2728 4924
rect 2664 4864 2728 4868
rect 2744 4924 2808 4928
rect 2744 4868 2748 4924
rect 2748 4868 2804 4924
rect 2804 4868 2808 4924
rect 2744 4864 2808 4868
rect 2824 4924 2888 4928
rect 2824 4868 2828 4924
rect 2828 4868 2884 4924
rect 2884 4868 2888 4924
rect 2824 4864 2888 4868
rect 5848 4924 5912 4928
rect 5848 4868 5852 4924
rect 5852 4868 5908 4924
rect 5908 4868 5912 4924
rect 5848 4864 5912 4868
rect 5928 4924 5992 4928
rect 5928 4868 5932 4924
rect 5932 4868 5988 4924
rect 5988 4868 5992 4924
rect 5928 4864 5992 4868
rect 6008 4924 6072 4928
rect 6008 4868 6012 4924
rect 6012 4868 6068 4924
rect 6068 4868 6072 4924
rect 6008 4864 6072 4868
rect 6088 4924 6152 4928
rect 6088 4868 6092 4924
rect 6092 4868 6148 4924
rect 6148 4868 6152 4924
rect 6088 4864 6152 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 9272 4924 9336 4928
rect 9272 4868 9276 4924
rect 9276 4868 9332 4924
rect 9332 4868 9336 4924
rect 9272 4864 9336 4868
rect 9352 4924 9416 4928
rect 9352 4868 9356 4924
rect 9356 4868 9412 4924
rect 9412 4868 9416 4924
rect 9352 4864 9416 4868
rect 4660 4796 4724 4860
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 7480 4380 7544 4384
rect 7480 4324 7484 4380
rect 7484 4324 7540 4380
rect 7540 4324 7544 4380
rect 7480 4320 7544 4324
rect 7560 4380 7624 4384
rect 7560 4324 7564 4380
rect 7564 4324 7620 4380
rect 7620 4324 7624 4380
rect 7560 4320 7624 4324
rect 7640 4380 7704 4384
rect 7640 4324 7644 4380
rect 7644 4324 7700 4380
rect 7700 4324 7704 4380
rect 7640 4320 7704 4324
rect 7720 4380 7784 4384
rect 7720 4324 7724 4380
rect 7724 4324 7780 4380
rect 7780 4324 7784 4380
rect 7720 4320 7784 4324
rect 2584 3836 2648 3840
rect 2584 3780 2588 3836
rect 2588 3780 2644 3836
rect 2644 3780 2648 3836
rect 2584 3776 2648 3780
rect 2664 3836 2728 3840
rect 2664 3780 2668 3836
rect 2668 3780 2724 3836
rect 2724 3780 2728 3836
rect 2664 3776 2728 3780
rect 2744 3836 2808 3840
rect 2744 3780 2748 3836
rect 2748 3780 2804 3836
rect 2804 3780 2808 3836
rect 2744 3776 2808 3780
rect 2824 3836 2888 3840
rect 2824 3780 2828 3836
rect 2828 3780 2884 3836
rect 2884 3780 2888 3836
rect 2824 3776 2888 3780
rect 5848 3836 5912 3840
rect 5848 3780 5852 3836
rect 5852 3780 5908 3836
rect 5908 3780 5912 3836
rect 5848 3776 5912 3780
rect 5928 3836 5992 3840
rect 5928 3780 5932 3836
rect 5932 3780 5988 3836
rect 5988 3780 5992 3836
rect 5928 3776 5992 3780
rect 6008 3836 6072 3840
rect 6008 3780 6012 3836
rect 6012 3780 6068 3836
rect 6068 3780 6072 3836
rect 6008 3776 6072 3780
rect 6088 3836 6152 3840
rect 6088 3780 6092 3836
rect 6092 3780 6148 3836
rect 6148 3780 6152 3836
rect 6088 3776 6152 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 9272 3836 9336 3840
rect 9272 3780 9276 3836
rect 9276 3780 9332 3836
rect 9332 3780 9336 3836
rect 9272 3776 9336 3780
rect 9352 3836 9416 3840
rect 9352 3780 9356 3836
rect 9356 3780 9412 3836
rect 9412 3780 9416 3836
rect 9352 3776 9416 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 7480 3292 7544 3296
rect 7480 3236 7484 3292
rect 7484 3236 7540 3292
rect 7540 3236 7544 3292
rect 7480 3232 7544 3236
rect 7560 3292 7624 3296
rect 7560 3236 7564 3292
rect 7564 3236 7620 3292
rect 7620 3236 7624 3292
rect 7560 3232 7624 3236
rect 7640 3292 7704 3296
rect 7640 3236 7644 3292
rect 7644 3236 7700 3292
rect 7700 3236 7704 3292
rect 7640 3232 7704 3236
rect 7720 3292 7784 3296
rect 7720 3236 7724 3292
rect 7724 3236 7780 3292
rect 7780 3236 7784 3292
rect 7720 3232 7784 3236
rect 2584 2748 2648 2752
rect 2584 2692 2588 2748
rect 2588 2692 2644 2748
rect 2644 2692 2648 2748
rect 2584 2688 2648 2692
rect 2664 2748 2728 2752
rect 2664 2692 2668 2748
rect 2668 2692 2724 2748
rect 2724 2692 2728 2748
rect 2664 2688 2728 2692
rect 2744 2748 2808 2752
rect 2744 2692 2748 2748
rect 2748 2692 2804 2748
rect 2804 2692 2808 2748
rect 2744 2688 2808 2692
rect 2824 2748 2888 2752
rect 2824 2692 2828 2748
rect 2828 2692 2884 2748
rect 2884 2692 2888 2748
rect 2824 2688 2888 2692
rect 5848 2748 5912 2752
rect 5848 2692 5852 2748
rect 5852 2692 5908 2748
rect 5908 2692 5912 2748
rect 5848 2688 5912 2692
rect 5928 2748 5992 2752
rect 5928 2692 5932 2748
rect 5932 2692 5988 2748
rect 5988 2692 5992 2748
rect 5928 2688 5992 2692
rect 6008 2748 6072 2752
rect 6008 2692 6012 2748
rect 6012 2692 6068 2748
rect 6068 2692 6072 2748
rect 6008 2688 6072 2692
rect 6088 2748 6152 2752
rect 6088 2692 6092 2748
rect 6092 2692 6148 2748
rect 6148 2692 6152 2748
rect 6088 2688 6152 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 9272 2748 9336 2752
rect 9272 2692 9276 2748
rect 9276 2692 9332 2748
rect 9332 2692 9336 2748
rect 9272 2688 9336 2692
rect 9352 2748 9416 2752
rect 9352 2692 9356 2748
rect 9356 2692 9412 2748
rect 9412 2692 9416 2748
rect 9352 2688 9416 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 7480 2204 7544 2208
rect 7480 2148 7484 2204
rect 7484 2148 7540 2204
rect 7540 2148 7544 2204
rect 7480 2144 7544 2148
rect 7560 2204 7624 2208
rect 7560 2148 7564 2204
rect 7564 2148 7620 2204
rect 7620 2148 7624 2204
rect 7560 2144 7624 2148
rect 7640 2204 7704 2208
rect 7640 2148 7644 2204
rect 7644 2148 7700 2204
rect 7700 2148 7704 2204
rect 7640 2144 7704 2148
rect 7720 2204 7784 2208
rect 7720 2148 7724 2204
rect 7724 2148 7780 2204
rect 7780 2148 7784 2204
rect 7720 2144 7784 2148
<< metal4 >>
rect 2576 77824 2896 77840
rect 2576 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2576 76736 2896 77760
rect 2576 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2576 75648 2896 76672
rect 2576 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2576 74560 2896 75584
rect 4208 77280 4528 77840
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 76192 4528 77216
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 75104 4528 76128
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 3923 75036 3989 75037
rect 3923 74972 3924 75036
rect 3988 74972 3989 75036
rect 3923 74971 3989 74972
rect 2576 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2576 73472 2896 74496
rect 2576 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2576 72384 2896 73408
rect 2576 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2576 71296 2896 72320
rect 2576 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2576 70208 2896 71232
rect 2576 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2267 69324 2333 69325
rect 2267 69260 2268 69324
rect 2332 69260 2333 69324
rect 2267 69259 2333 69260
rect 1715 67692 1781 67693
rect 1715 67628 1716 67692
rect 1780 67628 1781 67692
rect 1715 67627 1781 67628
rect 1347 64972 1413 64973
rect 1347 64908 1348 64972
rect 1412 64908 1413 64972
rect 1347 64907 1413 64908
rect 59 56404 125 56405
rect 59 56340 60 56404
rect 124 56340 125 56404
rect 59 56339 125 56340
rect 62 50421 122 56339
rect 1163 55452 1229 55453
rect 1163 55388 1164 55452
rect 1228 55388 1229 55452
rect 1163 55387 1229 55388
rect 979 55180 1045 55181
rect 979 55178 980 55180
rect 798 55118 980 55178
rect 798 54770 858 55118
rect 979 55116 980 55118
rect 1044 55116 1045 55180
rect 979 55115 1045 55116
rect 1166 54909 1226 55387
rect 1163 54908 1229 54909
rect 1163 54844 1164 54908
rect 1228 54844 1229 54908
rect 1163 54843 1229 54844
rect 430 54710 858 54770
rect 979 54772 1045 54773
rect 59 50420 125 50421
rect 59 50356 60 50420
rect 124 50356 125 50420
rect 59 50355 125 50356
rect 243 47428 309 47429
rect 243 47364 244 47428
rect 308 47364 309 47428
rect 243 47363 309 47364
rect 59 46578 125 46579
rect 59 46514 60 46578
rect 124 46514 125 46578
rect 59 46513 125 46514
rect 62 41445 122 46513
rect 59 41444 125 41445
rect 59 41380 60 41444
rect 124 41380 125 41444
rect 59 41379 125 41380
rect 246 38670 306 47363
rect 430 44570 490 54710
rect 979 54708 980 54772
rect 1044 54708 1045 54772
rect 979 54707 1045 54708
rect 982 52730 1042 54707
rect 614 52670 1042 52730
rect 614 48330 674 52670
rect 979 51644 1045 51645
rect 979 51580 980 51644
rect 1044 51580 1045 51644
rect 979 51579 1045 51580
rect 982 50965 1042 51579
rect 1163 51372 1229 51373
rect 1163 51308 1164 51372
rect 1228 51308 1229 51372
rect 1163 51307 1229 51308
rect 979 50964 1045 50965
rect 979 50900 980 50964
rect 1044 50900 1045 50964
rect 979 50899 1045 50900
rect 979 50828 1045 50829
rect 979 50764 980 50828
rect 1044 50764 1045 50828
rect 979 50763 1045 50764
rect 614 48270 858 48330
rect 430 44510 674 44570
rect 614 44437 674 44510
rect 427 44436 493 44437
rect 427 44372 428 44436
rect 492 44372 493 44436
rect 427 44371 493 44372
rect 611 44436 677 44437
rect 611 44372 612 44436
rect 676 44372 677 44436
rect 611 44371 677 44372
rect 430 38861 490 44371
rect 427 38860 493 38861
rect 427 38796 428 38860
rect 492 38796 493 38860
rect 427 38795 493 38796
rect 246 38610 674 38670
rect 614 22110 674 38610
rect 798 32877 858 48270
rect 982 46882 1042 50763
rect 1166 48381 1226 51307
rect 1163 48380 1229 48381
rect 1163 48316 1164 48380
rect 1228 48316 1229 48380
rect 1163 48315 1229 48316
rect 982 46822 1226 46882
rect 1166 45250 1226 46822
rect 1350 45389 1410 64907
rect 1531 62252 1597 62253
rect 1531 62188 1532 62252
rect 1596 62188 1597 62252
rect 1531 62187 1597 62188
rect 1534 46885 1594 62187
rect 1718 50421 1778 67627
rect 2083 67420 2149 67421
rect 2083 67356 2084 67420
rect 2148 67356 2149 67420
rect 2083 67355 2149 67356
rect 1899 62932 1965 62933
rect 1899 62868 1900 62932
rect 1964 62868 1965 62932
rect 1899 62867 1965 62868
rect 1715 50420 1781 50421
rect 1715 50356 1716 50420
rect 1780 50356 1781 50420
rect 1715 50355 1781 50356
rect 1715 50284 1781 50285
rect 1715 50220 1716 50284
rect 1780 50220 1781 50284
rect 1715 50219 1781 50220
rect 1531 46884 1597 46885
rect 1531 46820 1532 46884
rect 1596 46820 1597 46884
rect 1531 46819 1597 46820
rect 1531 46612 1597 46613
rect 1531 46548 1532 46612
rect 1596 46548 1597 46612
rect 1531 46547 1597 46548
rect 1347 45388 1413 45389
rect 1347 45324 1348 45388
rect 1412 45324 1413 45388
rect 1347 45323 1413 45324
rect 1166 45190 1410 45250
rect 979 44436 1045 44437
rect 979 44372 980 44436
rect 1044 44372 1045 44436
rect 979 44371 1045 44372
rect 795 32876 861 32877
rect 795 32812 796 32876
rect 860 32812 861 32876
rect 795 32811 861 32812
rect 982 30293 1042 44371
rect 1163 44300 1229 44301
rect 1163 44236 1164 44300
rect 1228 44236 1229 44300
rect 1163 44235 1229 44236
rect 1166 32877 1226 44235
rect 1350 42805 1410 45190
rect 1534 43757 1594 46547
rect 1531 43756 1597 43757
rect 1531 43692 1532 43756
rect 1596 43692 1597 43756
rect 1531 43691 1597 43692
rect 1531 43484 1597 43485
rect 1531 43420 1532 43484
rect 1596 43420 1597 43484
rect 1531 43419 1597 43420
rect 1347 42804 1413 42805
rect 1347 42740 1348 42804
rect 1412 42740 1413 42804
rect 1347 42739 1413 42740
rect 1347 42668 1413 42669
rect 1347 42604 1348 42668
rect 1412 42604 1413 42668
rect 1347 42603 1413 42604
rect 1350 41581 1410 42603
rect 1347 41580 1413 41581
rect 1347 41516 1348 41580
rect 1412 41516 1413 41580
rect 1347 41515 1413 41516
rect 1347 41308 1413 41309
rect 1347 41244 1348 41308
rect 1412 41244 1413 41308
rect 1347 41243 1413 41244
rect 1350 33285 1410 41243
rect 1347 33284 1413 33285
rect 1347 33220 1348 33284
rect 1412 33220 1413 33284
rect 1347 33219 1413 33220
rect 1163 32876 1229 32877
rect 1163 32812 1164 32876
rect 1228 32812 1229 32876
rect 1163 32811 1229 32812
rect 1534 32741 1594 43419
rect 1718 42805 1778 50219
rect 1902 48245 1962 62867
rect 2086 61165 2146 67355
rect 2270 64157 2330 69259
rect 2576 69120 2896 70144
rect 2576 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2576 68032 2896 69056
rect 2576 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2576 66944 2896 67968
rect 2576 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2576 65856 2896 66880
rect 2576 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2576 64768 2896 65792
rect 2576 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2267 64156 2333 64157
rect 2267 64092 2268 64156
rect 2332 64092 2333 64156
rect 2267 64091 2333 64092
rect 2576 63680 2896 64704
rect 2576 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2576 62592 2896 63616
rect 3555 63476 3621 63477
rect 3555 63412 3556 63476
rect 3620 63412 3621 63476
rect 3555 63411 3621 63412
rect 2576 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2576 61504 2896 62528
rect 3371 61844 3437 61845
rect 3371 61780 3372 61844
rect 3436 61780 3437 61844
rect 3371 61779 3437 61780
rect 2576 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2267 61300 2333 61301
rect 2267 61236 2268 61300
rect 2332 61236 2333 61300
rect 2267 61235 2333 61236
rect 2083 61164 2149 61165
rect 2083 61100 2084 61164
rect 2148 61100 2149 61164
rect 2083 61099 2149 61100
rect 2083 61028 2149 61029
rect 2083 60964 2084 61028
rect 2148 60964 2149 61028
rect 2083 60963 2149 60964
rect 2086 55181 2146 60963
rect 2270 59533 2330 61235
rect 2576 60416 2896 61440
rect 3187 61028 3253 61029
rect 3187 60964 3188 61028
rect 3252 60964 3253 61028
rect 3187 60963 3253 60964
rect 3003 60892 3069 60893
rect 3003 60828 3004 60892
rect 3068 60828 3069 60892
rect 3003 60827 3069 60828
rect 3006 60485 3066 60827
rect 3003 60484 3069 60485
rect 3003 60420 3004 60484
rect 3068 60420 3069 60484
rect 3003 60419 3069 60420
rect 2576 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2267 59532 2333 59533
rect 2267 59468 2268 59532
rect 2332 59468 2333 59532
rect 2267 59467 2333 59468
rect 2576 59328 2896 60352
rect 2576 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2576 58240 2896 59264
rect 2576 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2267 57628 2333 57629
rect 2267 57564 2268 57628
rect 2332 57564 2333 57628
rect 2267 57563 2333 57564
rect 2270 57490 2330 57563
rect 2270 57430 2514 57490
rect 2267 57356 2333 57357
rect 2267 57292 2268 57356
rect 2332 57292 2333 57356
rect 2267 57291 2333 57292
rect 2083 55180 2149 55181
rect 2083 55116 2084 55180
rect 2148 55116 2149 55180
rect 2083 55115 2149 55116
rect 2083 54364 2149 54365
rect 2083 54300 2084 54364
rect 2148 54300 2149 54364
rect 2083 54299 2149 54300
rect 2086 51373 2146 54299
rect 2083 51372 2149 51373
rect 2083 51308 2084 51372
rect 2148 51308 2149 51372
rect 2083 51307 2149 51308
rect 2270 50690 2330 57291
rect 2086 50630 2330 50690
rect 1899 48244 1965 48245
rect 1899 48180 1900 48244
rect 1964 48180 1965 48244
rect 1899 48179 1965 48180
rect 1899 48108 1965 48109
rect 1899 48044 1900 48108
rect 1964 48044 1965 48108
rect 1899 48043 1965 48044
rect 1902 43077 1962 48043
rect 2086 43893 2146 50630
rect 2267 49196 2333 49197
rect 2267 49132 2268 49196
rect 2332 49194 2333 49196
rect 2454 49194 2514 57430
rect 2332 49134 2514 49194
rect 2576 57152 2896 58176
rect 2576 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2576 56064 2896 57088
rect 2576 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2576 54976 2896 56000
rect 3003 55180 3069 55181
rect 3003 55116 3004 55180
rect 3068 55116 3069 55180
rect 3003 55115 3069 55116
rect 2576 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2576 53888 2896 54912
rect 2576 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2576 52800 2896 53824
rect 2576 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2576 51712 2896 52736
rect 2576 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2576 50624 2896 51648
rect 2576 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2576 49536 2896 50560
rect 2576 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2332 49132 2333 49134
rect 2267 49131 2333 49132
rect 2576 48448 2896 49472
rect 2576 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2267 47972 2333 47973
rect 2267 47908 2268 47972
rect 2332 47908 2333 47972
rect 2267 47907 2333 47908
rect 2083 43892 2149 43893
rect 2083 43828 2084 43892
rect 2148 43828 2149 43892
rect 2083 43827 2149 43828
rect 2083 43756 2149 43757
rect 2083 43692 2084 43756
rect 2148 43692 2149 43756
rect 2083 43691 2149 43692
rect 1899 43076 1965 43077
rect 1899 43012 1900 43076
rect 1964 43012 1965 43076
rect 1899 43011 1965 43012
rect 1899 42940 1965 42941
rect 1899 42876 1900 42940
rect 1964 42876 1965 42940
rect 1899 42875 1965 42876
rect 1715 42804 1781 42805
rect 1715 42740 1716 42804
rect 1780 42740 1781 42804
rect 1715 42739 1781 42740
rect 1715 42396 1781 42397
rect 1715 42332 1716 42396
rect 1780 42332 1781 42396
rect 1715 42331 1781 42332
rect 1718 41309 1778 42331
rect 1715 41308 1781 41309
rect 1715 41244 1716 41308
rect 1780 41244 1781 41308
rect 1715 41243 1781 41244
rect 1715 39404 1781 39405
rect 1715 39340 1716 39404
rect 1780 39340 1781 39404
rect 1715 39339 1781 39340
rect 1531 32740 1597 32741
rect 1531 32676 1532 32740
rect 1596 32676 1597 32740
rect 1531 32675 1597 32676
rect 1718 32197 1778 39339
rect 1902 36141 1962 42875
rect 2086 42669 2146 43691
rect 2083 42668 2149 42669
rect 2083 42604 2084 42668
rect 2148 42604 2149 42668
rect 2083 42603 2149 42604
rect 2083 41852 2149 41853
rect 2083 41788 2084 41852
rect 2148 41788 2149 41852
rect 2083 41787 2149 41788
rect 2086 38997 2146 41787
rect 2083 38996 2149 38997
rect 2083 38932 2084 38996
rect 2148 38932 2149 38996
rect 2083 38931 2149 38932
rect 2083 38860 2149 38861
rect 2083 38796 2084 38860
rect 2148 38796 2149 38860
rect 2083 38795 2149 38796
rect 2086 38181 2146 38795
rect 2083 38180 2149 38181
rect 2083 38116 2084 38180
rect 2148 38116 2149 38180
rect 2083 38115 2149 38116
rect 1899 36140 1965 36141
rect 1899 36076 1900 36140
rect 1964 36076 1965 36140
rect 1899 36075 1965 36076
rect 1715 32196 1781 32197
rect 1715 32132 1716 32196
rect 1780 32132 1781 32196
rect 1715 32131 1781 32132
rect 1531 31924 1597 31925
rect 1531 31860 1532 31924
rect 1596 31860 1597 31924
rect 1531 31859 1597 31860
rect 1534 31517 1594 31859
rect 1531 31516 1597 31517
rect 1531 31452 1532 31516
rect 1596 31452 1597 31516
rect 1531 31451 1597 31452
rect 979 30292 1045 30293
rect 979 30228 980 30292
rect 1044 30228 1045 30292
rect 979 30227 1045 30228
rect 2086 28253 2146 38115
rect 2270 36821 2330 47907
rect 2405 47836 2471 47837
rect 2405 47772 2406 47836
rect 2470 47834 2471 47836
rect 2470 47772 2514 47834
rect 2405 47771 2514 47772
rect 2454 45661 2514 47771
rect 2405 45660 2514 45661
rect 2405 45596 2406 45660
rect 2470 45598 2514 45660
rect 2576 47360 2896 48384
rect 2576 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2576 46272 2896 47296
rect 2576 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2470 45596 2471 45598
rect 2405 45595 2471 45596
rect 2405 45388 2471 45389
rect 2405 45324 2406 45388
rect 2470 45386 2471 45388
rect 2470 45324 2514 45386
rect 2405 45323 2514 45324
rect 2454 40493 2514 45323
rect 2405 40492 2514 40493
rect 2405 40428 2406 40492
rect 2470 40430 2514 40492
rect 2576 45184 2896 46208
rect 3006 45797 3066 55115
rect 3190 53549 3250 60963
rect 3374 60349 3434 61779
rect 3371 60348 3437 60349
rect 3371 60284 3372 60348
rect 3436 60284 3437 60348
rect 3371 60283 3437 60284
rect 3558 58581 3618 63411
rect 3739 60620 3805 60621
rect 3739 60556 3740 60620
rect 3804 60556 3805 60620
rect 3739 60555 3805 60556
rect 3555 58580 3621 58581
rect 3555 58516 3556 58580
rect 3620 58516 3621 58580
rect 3555 58515 3621 58516
rect 3371 55724 3437 55725
rect 3371 55660 3372 55724
rect 3436 55660 3437 55724
rect 3371 55659 3437 55660
rect 3187 53548 3253 53549
rect 3187 53484 3188 53548
rect 3252 53484 3253 53548
rect 3187 53483 3253 53484
rect 3187 53412 3253 53413
rect 3187 53348 3188 53412
rect 3252 53348 3253 53412
rect 3187 53347 3253 53348
rect 3003 45796 3069 45797
rect 3003 45732 3004 45796
rect 3068 45732 3069 45796
rect 3003 45731 3069 45732
rect 3003 45660 3069 45661
rect 3003 45596 3004 45660
rect 3068 45596 3069 45660
rect 3003 45595 3069 45596
rect 2576 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2576 44096 2896 45120
rect 2576 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2576 43008 2896 44032
rect 2576 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2576 41920 2896 42944
rect 2576 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2576 40832 2896 41856
rect 2576 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2470 40428 2471 40430
rect 2405 40427 2471 40428
rect 2576 39744 2896 40768
rect 2576 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2576 38656 2896 39680
rect 2576 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2576 37568 2896 38592
rect 2576 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2267 36820 2333 36821
rect 2267 36756 2268 36820
rect 2332 36756 2333 36820
rect 2267 36755 2333 36756
rect 2267 36548 2333 36549
rect 2267 36484 2268 36548
rect 2332 36484 2333 36548
rect 2267 36483 2333 36484
rect 2083 28252 2149 28253
rect 2083 28188 2084 28252
rect 2148 28188 2149 28252
rect 2083 28187 2149 28188
rect 2270 23901 2330 36483
rect 2576 36480 2896 37504
rect 2576 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2576 35392 2896 36416
rect 2576 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2576 34304 2896 35328
rect 2576 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2576 33216 2896 34240
rect 2576 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2576 32128 2896 33152
rect 2576 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2576 31040 2896 32064
rect 2576 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2576 29952 2896 30976
rect 2576 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2576 28864 2896 29888
rect 2576 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2576 27776 2896 28800
rect 2576 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2576 26688 2896 27712
rect 2576 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2576 25600 2896 26624
rect 2576 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2576 24512 2896 25536
rect 2576 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2267 23900 2333 23901
rect 2267 23836 2268 23900
rect 2332 23836 2333 23900
rect 2267 23835 2333 23836
rect 2576 23424 2896 24448
rect 2576 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2576 22336 2896 23360
rect 2576 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2267 22268 2333 22269
rect 2267 22204 2268 22268
rect 2332 22204 2333 22268
rect 2267 22203 2333 22204
rect 614 22050 1042 22110
rect 982 6765 1042 22050
rect 2270 21997 2330 22203
rect 2267 21996 2333 21997
rect 2267 21932 2268 21996
rect 2332 21932 2333 21996
rect 2267 21931 2333 21932
rect 2576 21248 2896 22272
rect 2576 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2576 20160 2896 21184
rect 2576 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2576 19072 2896 20096
rect 2576 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2576 17984 2896 19008
rect 2576 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2576 16896 2896 17920
rect 2576 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2576 15808 2896 16832
rect 2576 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2576 14720 2896 15744
rect 2576 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2576 13632 2896 14656
rect 2576 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 1899 13156 1965 13157
rect 1899 13092 1900 13156
rect 1964 13092 1965 13156
rect 1899 13091 1965 13092
rect 1902 12477 1962 13091
rect 2576 12544 2896 13568
rect 2576 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 1899 12476 1965 12477
rect 1899 12412 1900 12476
rect 1964 12412 1965 12476
rect 1899 12411 1965 12412
rect 2576 11456 2896 12480
rect 2576 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2576 10368 2896 11392
rect 2576 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2576 9280 2896 10304
rect 2576 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2576 8192 2896 9216
rect 3006 9213 3066 45595
rect 3190 45389 3250 53347
rect 3374 51373 3434 55659
rect 3742 52733 3802 60555
rect 3739 52732 3805 52733
rect 3739 52668 3740 52732
rect 3804 52668 3805 52732
rect 3739 52667 3805 52668
rect 3371 51372 3437 51373
rect 3371 51308 3372 51372
rect 3436 51308 3437 51372
rect 3371 51307 3437 51308
rect 3371 51236 3437 51237
rect 3371 51172 3372 51236
rect 3436 51172 3437 51236
rect 3371 51171 3437 51172
rect 3374 50965 3434 51171
rect 3371 50964 3437 50965
rect 3371 50900 3372 50964
rect 3436 50900 3437 50964
rect 3371 50899 3437 50900
rect 3555 50964 3621 50965
rect 3555 50900 3556 50964
rect 3620 50900 3621 50964
rect 3555 50899 3621 50900
rect 3371 50148 3437 50149
rect 3371 50084 3372 50148
rect 3436 50084 3437 50148
rect 3371 50083 3437 50084
rect 3187 45388 3253 45389
rect 3187 45324 3188 45388
rect 3252 45324 3253 45388
rect 3187 45323 3253 45324
rect 3374 44709 3434 50083
rect 3371 44708 3437 44709
rect 3371 44644 3372 44708
rect 3436 44644 3437 44708
rect 3371 44643 3437 44644
rect 3558 44570 3618 50899
rect 3739 50012 3805 50013
rect 3739 49948 3740 50012
rect 3804 49948 3805 50012
rect 3739 49947 3805 49948
rect 3742 48245 3802 49947
rect 3739 48244 3805 48245
rect 3739 48180 3740 48244
rect 3804 48180 3805 48244
rect 3739 48179 3805 48180
rect 3739 47836 3805 47837
rect 3739 47772 3740 47836
rect 3804 47772 3805 47836
rect 3739 47771 3805 47772
rect 3190 44510 3618 44570
rect 3190 43077 3250 44510
rect 3371 44436 3437 44437
rect 3371 44372 3372 44436
rect 3436 44372 3437 44436
rect 3371 44371 3437 44372
rect 3187 43076 3253 43077
rect 3187 43012 3188 43076
rect 3252 43012 3253 43076
rect 3187 43011 3253 43012
rect 3187 42940 3253 42941
rect 3187 42876 3188 42940
rect 3252 42876 3253 42940
rect 3187 42875 3253 42876
rect 3190 41850 3250 42875
rect 3374 41989 3434 44371
rect 3555 43212 3621 43213
rect 3555 43148 3556 43212
rect 3620 43148 3621 43212
rect 3555 43147 3621 43148
rect 3371 41988 3437 41989
rect 3371 41924 3372 41988
rect 3436 41924 3437 41988
rect 3371 41923 3437 41924
rect 3190 41790 3434 41850
rect 3187 41444 3253 41445
rect 3187 41380 3188 41444
rect 3252 41380 3253 41444
rect 3187 41379 3253 41380
rect 3190 39269 3250 41379
rect 3374 41173 3434 41790
rect 3558 41309 3618 43147
rect 3742 41850 3802 47771
rect 3926 42805 3986 74971
rect 4208 74016 4528 75040
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 72928 4528 73952
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 71840 4528 72864
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 70752 4528 71776
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 69664 4528 70688
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 68576 4528 69600
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 67488 4528 68512
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 66400 4528 67424
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 65312 4528 66336
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 64224 4528 65248
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 63136 4528 64160
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 62048 4528 63072
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 60960 4528 61984
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 59872 4528 60896
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 58784 4528 59808
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 57696 4528 58720
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 56608 4528 57632
rect 5840 77824 6160 77840
rect 5840 77760 5848 77824
rect 5912 77760 5928 77824
rect 5992 77760 6008 77824
rect 6072 77760 6088 77824
rect 6152 77760 6160 77824
rect 5840 76736 6160 77760
rect 5840 76672 5848 76736
rect 5912 76672 5928 76736
rect 5992 76672 6008 76736
rect 6072 76672 6088 76736
rect 6152 76672 6160 76736
rect 5840 75648 6160 76672
rect 5840 75584 5848 75648
rect 5912 75584 5928 75648
rect 5992 75584 6008 75648
rect 6072 75584 6088 75648
rect 6152 75584 6160 75648
rect 5840 74560 6160 75584
rect 5840 74496 5848 74560
rect 5912 74496 5928 74560
rect 5992 74496 6008 74560
rect 6072 74496 6088 74560
rect 6152 74496 6160 74560
rect 5840 73472 6160 74496
rect 5840 73408 5848 73472
rect 5912 73408 5928 73472
rect 5992 73408 6008 73472
rect 6072 73408 6088 73472
rect 6152 73408 6160 73472
rect 5840 72384 6160 73408
rect 5840 72320 5848 72384
rect 5912 72320 5928 72384
rect 5992 72320 6008 72384
rect 6072 72320 6088 72384
rect 6152 72320 6160 72384
rect 5840 71296 6160 72320
rect 5840 71232 5848 71296
rect 5912 71232 5928 71296
rect 5992 71232 6008 71296
rect 6072 71232 6088 71296
rect 6152 71232 6160 71296
rect 5840 70208 6160 71232
rect 5840 70144 5848 70208
rect 5912 70144 5928 70208
rect 5992 70144 6008 70208
rect 6072 70144 6088 70208
rect 6152 70144 6160 70208
rect 5840 69120 6160 70144
rect 5840 69056 5848 69120
rect 5912 69056 5928 69120
rect 5992 69056 6008 69120
rect 6072 69056 6088 69120
rect 6152 69056 6160 69120
rect 5840 68032 6160 69056
rect 5840 67968 5848 68032
rect 5912 67968 5928 68032
rect 5992 67968 6008 68032
rect 6072 67968 6088 68032
rect 6152 67968 6160 68032
rect 5840 66944 6160 67968
rect 5840 66880 5848 66944
rect 5912 66880 5928 66944
rect 5992 66880 6008 66944
rect 6072 66880 6088 66944
rect 6152 66880 6160 66944
rect 5840 65856 6160 66880
rect 5840 65792 5848 65856
rect 5912 65792 5928 65856
rect 5992 65792 6008 65856
rect 6072 65792 6088 65856
rect 6152 65792 6160 65856
rect 5840 64768 6160 65792
rect 5840 64704 5848 64768
rect 5912 64704 5928 64768
rect 5992 64704 6008 64768
rect 6072 64704 6088 64768
rect 6152 64704 6160 64768
rect 5840 63680 6160 64704
rect 5840 63616 5848 63680
rect 5912 63616 5928 63680
rect 5992 63616 6008 63680
rect 6072 63616 6088 63680
rect 6152 63616 6160 63680
rect 5840 62592 6160 63616
rect 5840 62528 5848 62592
rect 5912 62528 5928 62592
rect 5992 62528 6008 62592
rect 6072 62528 6088 62592
rect 6152 62528 6160 62592
rect 5840 61504 6160 62528
rect 5840 61440 5848 61504
rect 5912 61440 5928 61504
rect 5992 61440 6008 61504
rect 6072 61440 6088 61504
rect 6152 61440 6160 61504
rect 5840 60416 6160 61440
rect 5840 60352 5848 60416
rect 5912 60352 5928 60416
rect 5992 60352 6008 60416
rect 6072 60352 6088 60416
rect 6152 60352 6160 60416
rect 5840 59328 6160 60352
rect 5840 59264 5848 59328
rect 5912 59264 5928 59328
rect 5992 59264 6008 59328
rect 6072 59264 6088 59328
rect 6152 59264 6160 59328
rect 5840 58240 6160 59264
rect 5840 58176 5848 58240
rect 5912 58176 5928 58240
rect 5992 58176 6008 58240
rect 6072 58176 6088 58240
rect 6152 58176 6160 58240
rect 5579 57492 5645 57493
rect 5579 57428 5580 57492
rect 5644 57428 5645 57492
rect 5579 57427 5645 57428
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 55520 4528 56544
rect 4659 55724 4725 55725
rect 4659 55660 4660 55724
rect 4724 55660 4725 55724
rect 4659 55659 4725 55660
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 54432 4528 55456
rect 4662 55181 4722 55659
rect 4659 55180 4725 55181
rect 4659 55116 4660 55180
rect 4724 55116 4725 55180
rect 4659 55115 4725 55116
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 53344 4528 54368
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 52256 4528 53280
rect 4662 52869 4722 55115
rect 4843 53548 4909 53549
rect 4843 53484 4844 53548
rect 4908 53484 4909 53548
rect 4843 53483 4909 53484
rect 4659 52868 4725 52869
rect 4659 52804 4660 52868
rect 4724 52804 4725 52868
rect 4659 52803 4725 52804
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 51168 4528 52192
rect 4659 51508 4725 51509
rect 4659 51444 4660 51508
rect 4724 51444 4725 51508
rect 4659 51443 4725 51444
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 50080 4528 51104
rect 4662 50693 4722 51443
rect 4659 50692 4725 50693
rect 4659 50628 4660 50692
rect 4724 50628 4725 50692
rect 4659 50627 4725 50628
rect 4659 50420 4725 50421
rect 4659 50356 4660 50420
rect 4724 50356 4725 50420
rect 4659 50355 4725 50356
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 48992 4528 50016
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 47904 4528 48928
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 46816 4528 47840
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4662 45661 4722 50355
rect 4846 50285 4906 53483
rect 5395 52732 5461 52733
rect 5395 52668 5396 52732
rect 5460 52668 5461 52732
rect 5395 52667 5461 52668
rect 5211 52188 5277 52189
rect 5211 52124 5212 52188
rect 5276 52124 5277 52188
rect 5211 52123 5277 52124
rect 5027 51092 5093 51093
rect 5027 51028 5028 51092
rect 5092 51028 5093 51092
rect 5027 51027 5093 51028
rect 4843 50284 4909 50285
rect 4843 50220 4844 50284
rect 4908 50220 4909 50284
rect 4843 50219 4909 50220
rect 4843 47020 4909 47021
rect 4843 46956 4844 47020
rect 4908 46956 4909 47020
rect 4843 46955 4909 46956
rect 4659 45660 4725 45661
rect 4659 45596 4660 45660
rect 4724 45596 4725 45660
rect 4659 45595 4725 45596
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 3923 42804 3989 42805
rect 3923 42740 3924 42804
rect 3988 42740 3989 42804
rect 3923 42739 3989 42740
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 3742 41790 3986 41850
rect 3739 41580 3805 41581
rect 3739 41516 3740 41580
rect 3804 41516 3805 41580
rect 3739 41515 3805 41516
rect 3555 41308 3621 41309
rect 3555 41244 3556 41308
rect 3620 41244 3621 41308
rect 3555 41243 3621 41244
rect 3371 41172 3437 41173
rect 3371 41108 3372 41172
rect 3436 41108 3437 41172
rect 3371 41107 3437 41108
rect 3371 41036 3437 41037
rect 3371 40972 3372 41036
rect 3436 40972 3437 41036
rect 3371 40971 3437 40972
rect 3555 41036 3621 41037
rect 3555 40972 3556 41036
rect 3620 40972 3621 41036
rect 3555 40971 3621 40972
rect 3187 39268 3253 39269
rect 3187 39204 3188 39268
rect 3252 39204 3253 39268
rect 3187 39203 3253 39204
rect 3187 38316 3253 38317
rect 3187 38252 3188 38316
rect 3252 38252 3253 38316
rect 3187 38251 3253 38252
rect 3190 24853 3250 38251
rect 3374 37909 3434 40971
rect 3558 38861 3618 40971
rect 3555 38860 3621 38861
rect 3555 38796 3556 38860
rect 3620 38796 3621 38860
rect 3555 38795 3621 38796
rect 3371 37908 3437 37909
rect 3371 37844 3372 37908
rect 3436 37844 3437 37908
rect 3371 37843 3437 37844
rect 3558 32061 3618 38795
rect 3742 35325 3802 41515
rect 3926 41445 3986 41790
rect 3923 41444 3989 41445
rect 3923 41380 3924 41444
rect 3988 41380 3989 41444
rect 3923 41379 3989 41380
rect 4208 41376 4528 42400
rect 4846 41989 4906 46955
rect 5030 46477 5090 51027
rect 5214 50829 5274 52123
rect 5211 50828 5277 50829
rect 5211 50764 5212 50828
rect 5276 50764 5277 50828
rect 5211 50763 5277 50764
rect 5398 50693 5458 52667
rect 5395 50692 5461 50693
rect 5395 50628 5396 50692
rect 5460 50628 5461 50692
rect 5395 50627 5461 50628
rect 5211 49332 5277 49333
rect 5211 49268 5212 49332
rect 5276 49268 5277 49332
rect 5211 49267 5277 49268
rect 5027 46476 5093 46477
rect 5027 46412 5028 46476
rect 5092 46412 5093 46476
rect 5027 46411 5093 46412
rect 5027 46068 5093 46069
rect 5027 46004 5028 46068
rect 5092 46004 5093 46068
rect 5027 46003 5093 46004
rect 4843 41988 4909 41989
rect 4843 41924 4844 41988
rect 4908 41924 4909 41988
rect 4843 41923 4909 41924
rect 5030 41850 5090 46003
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 3923 39540 3989 39541
rect 3923 39476 3924 39540
rect 3988 39476 3989 39540
rect 3923 39475 3989 39476
rect 3739 35324 3805 35325
rect 3739 35260 3740 35324
rect 3804 35260 3805 35324
rect 3739 35259 3805 35260
rect 3739 35188 3805 35189
rect 3739 35124 3740 35188
rect 3804 35124 3805 35188
rect 3739 35123 3805 35124
rect 3555 32060 3621 32061
rect 3555 31996 3556 32060
rect 3620 31996 3621 32060
rect 3555 31995 3621 31996
rect 3371 29340 3437 29341
rect 3371 29276 3372 29340
rect 3436 29276 3437 29340
rect 3371 29275 3437 29276
rect 3374 27709 3434 29275
rect 3371 27708 3437 27709
rect 3371 27644 3372 27708
rect 3436 27644 3437 27708
rect 3371 27643 3437 27644
rect 3555 27572 3621 27573
rect 3555 27508 3556 27572
rect 3620 27508 3621 27572
rect 3555 27507 3621 27508
rect 3371 27436 3437 27437
rect 3371 27372 3372 27436
rect 3436 27372 3437 27436
rect 3371 27371 3437 27372
rect 3187 24852 3253 24853
rect 3187 24788 3188 24852
rect 3252 24788 3253 24852
rect 3187 24787 3253 24788
rect 3374 22813 3434 27371
rect 3371 22812 3437 22813
rect 3371 22748 3372 22812
rect 3436 22748 3437 22812
rect 3371 22747 3437 22748
rect 3558 22269 3618 27507
rect 3742 25261 3802 35123
rect 3926 32469 3986 39475
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 3923 32468 3989 32469
rect 3923 32404 3924 32468
rect 3988 32404 3989 32468
rect 3923 32403 3989 32404
rect 3923 32060 3989 32061
rect 3923 31996 3924 32060
rect 3988 31996 3989 32060
rect 3923 31995 3989 31996
rect 3739 25260 3805 25261
rect 3739 25196 3740 25260
rect 3804 25196 3805 25260
rect 3739 25195 3805 25196
rect 3926 24581 3986 31995
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 3923 24580 3989 24581
rect 3923 24516 3924 24580
rect 3988 24516 3989 24580
rect 3923 24515 3989 24516
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 3555 22268 3621 22269
rect 3555 22204 3556 22268
rect 3620 22204 3621 22268
rect 3555 22203 3621 22204
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 3003 9212 3069 9213
rect 3003 9148 3004 9212
rect 3068 9148 3069 9212
rect 3003 9147 3069 9148
rect 2576 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2576 7104 2896 8128
rect 2576 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 979 6764 1045 6765
rect 979 6700 980 6764
rect 1044 6700 1045 6764
rect 979 6699 1045 6700
rect 2576 6016 2896 7040
rect 2576 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2576 4928 2896 5952
rect 2576 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2576 3840 2896 4864
rect 2576 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2576 2752 2896 3776
rect 2576 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2576 2128 2896 2688
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4662 41790 5090 41850
rect 4662 4861 4722 41790
rect 5027 41580 5093 41581
rect 5027 41516 5028 41580
rect 5092 41516 5093 41580
rect 5027 41515 5093 41516
rect 4843 41444 4909 41445
rect 4843 41380 4844 41444
rect 4908 41380 4909 41444
rect 4843 41379 4909 41380
rect 4846 9485 4906 41379
rect 5030 36821 5090 41515
rect 5214 41445 5274 49267
rect 5395 49196 5461 49197
rect 5395 49132 5396 49196
rect 5460 49132 5461 49196
rect 5395 49131 5461 49132
rect 5398 42125 5458 49131
rect 5582 48517 5642 57427
rect 5840 57152 6160 58176
rect 5840 57088 5848 57152
rect 5912 57088 5928 57152
rect 5992 57088 6008 57152
rect 6072 57088 6088 57152
rect 6152 57088 6160 57152
rect 5840 56064 6160 57088
rect 5840 56000 5848 56064
rect 5912 56000 5928 56064
rect 5992 56000 6008 56064
rect 6072 56000 6088 56064
rect 6152 56000 6160 56064
rect 5840 54976 6160 56000
rect 5840 54912 5848 54976
rect 5912 54912 5928 54976
rect 5992 54912 6008 54976
rect 6072 54912 6088 54976
rect 6152 54912 6160 54976
rect 5840 53888 6160 54912
rect 5840 53824 5848 53888
rect 5912 53824 5928 53888
rect 5992 53824 6008 53888
rect 6072 53824 6088 53888
rect 6152 53824 6160 53888
rect 5840 52800 6160 53824
rect 5840 52736 5848 52800
rect 5912 52736 5928 52800
rect 5992 52736 6008 52800
rect 6072 52736 6088 52800
rect 6152 52736 6160 52800
rect 5840 51712 6160 52736
rect 5840 51648 5848 51712
rect 5912 51648 5928 51712
rect 5992 51648 6008 51712
rect 6072 51648 6088 51712
rect 6152 51648 6160 51712
rect 5840 50624 6160 51648
rect 5840 50560 5848 50624
rect 5912 50560 5928 50624
rect 5992 50560 6008 50624
rect 6072 50560 6088 50624
rect 6152 50560 6160 50624
rect 5840 49536 6160 50560
rect 5840 49472 5848 49536
rect 5912 49472 5928 49536
rect 5992 49472 6008 49536
rect 6072 49472 6088 49536
rect 6152 49472 6160 49536
rect 5579 48516 5645 48517
rect 5579 48452 5580 48516
rect 5644 48452 5645 48516
rect 5579 48451 5645 48452
rect 5840 48448 6160 49472
rect 5840 48384 5848 48448
rect 5912 48384 5928 48448
rect 5992 48384 6008 48448
rect 6072 48384 6088 48448
rect 6152 48384 6160 48448
rect 5840 47360 6160 48384
rect 7472 77280 7792 77840
rect 7472 77216 7480 77280
rect 7544 77216 7560 77280
rect 7624 77216 7640 77280
rect 7704 77216 7720 77280
rect 7784 77216 7792 77280
rect 7472 76192 7792 77216
rect 7472 76128 7480 76192
rect 7544 76128 7560 76192
rect 7624 76128 7640 76192
rect 7704 76128 7720 76192
rect 7784 76128 7792 76192
rect 7472 75104 7792 76128
rect 7472 75040 7480 75104
rect 7544 75040 7560 75104
rect 7624 75040 7640 75104
rect 7704 75040 7720 75104
rect 7784 75040 7792 75104
rect 7472 74016 7792 75040
rect 7472 73952 7480 74016
rect 7544 73952 7560 74016
rect 7624 73952 7640 74016
rect 7704 73952 7720 74016
rect 7784 73952 7792 74016
rect 7472 72928 7792 73952
rect 7472 72864 7480 72928
rect 7544 72864 7560 72928
rect 7624 72864 7640 72928
rect 7704 72864 7720 72928
rect 7784 72864 7792 72928
rect 7472 71840 7792 72864
rect 7472 71776 7480 71840
rect 7544 71776 7560 71840
rect 7624 71776 7640 71840
rect 7704 71776 7720 71840
rect 7784 71776 7792 71840
rect 7472 70752 7792 71776
rect 7472 70688 7480 70752
rect 7544 70688 7560 70752
rect 7624 70688 7640 70752
rect 7704 70688 7720 70752
rect 7784 70688 7792 70752
rect 7472 69664 7792 70688
rect 7472 69600 7480 69664
rect 7544 69600 7560 69664
rect 7624 69600 7640 69664
rect 7704 69600 7720 69664
rect 7784 69600 7792 69664
rect 7472 68576 7792 69600
rect 7472 68512 7480 68576
rect 7544 68512 7560 68576
rect 7624 68512 7640 68576
rect 7704 68512 7720 68576
rect 7784 68512 7792 68576
rect 7472 67488 7792 68512
rect 7472 67424 7480 67488
rect 7544 67424 7560 67488
rect 7624 67424 7640 67488
rect 7704 67424 7720 67488
rect 7784 67424 7792 67488
rect 7472 66400 7792 67424
rect 7472 66336 7480 66400
rect 7544 66336 7560 66400
rect 7624 66336 7640 66400
rect 7704 66336 7720 66400
rect 7784 66336 7792 66400
rect 7472 65312 7792 66336
rect 7472 65248 7480 65312
rect 7544 65248 7560 65312
rect 7624 65248 7640 65312
rect 7704 65248 7720 65312
rect 7784 65248 7792 65312
rect 7472 64224 7792 65248
rect 7472 64160 7480 64224
rect 7544 64160 7560 64224
rect 7624 64160 7640 64224
rect 7704 64160 7720 64224
rect 7784 64160 7792 64224
rect 7472 63136 7792 64160
rect 7472 63072 7480 63136
rect 7544 63072 7560 63136
rect 7624 63072 7640 63136
rect 7704 63072 7720 63136
rect 7784 63072 7792 63136
rect 7472 62048 7792 63072
rect 7472 61984 7480 62048
rect 7544 61984 7560 62048
rect 7624 61984 7640 62048
rect 7704 61984 7720 62048
rect 7784 61984 7792 62048
rect 7472 60960 7792 61984
rect 7472 60896 7480 60960
rect 7544 60896 7560 60960
rect 7624 60896 7640 60960
rect 7704 60896 7720 60960
rect 7784 60896 7792 60960
rect 7472 59872 7792 60896
rect 7472 59808 7480 59872
rect 7544 59808 7560 59872
rect 7624 59808 7640 59872
rect 7704 59808 7720 59872
rect 7784 59808 7792 59872
rect 7472 58784 7792 59808
rect 7472 58720 7480 58784
rect 7544 58720 7560 58784
rect 7624 58720 7640 58784
rect 7704 58720 7720 58784
rect 7784 58720 7792 58784
rect 7472 57696 7792 58720
rect 7472 57632 7480 57696
rect 7544 57632 7560 57696
rect 7624 57632 7640 57696
rect 7704 57632 7720 57696
rect 7784 57632 7792 57696
rect 7472 56608 7792 57632
rect 7472 56544 7480 56608
rect 7544 56544 7560 56608
rect 7624 56544 7640 56608
rect 7704 56544 7720 56608
rect 7784 56544 7792 56608
rect 7472 55520 7792 56544
rect 7472 55456 7480 55520
rect 7544 55456 7560 55520
rect 7624 55456 7640 55520
rect 7704 55456 7720 55520
rect 7784 55456 7792 55520
rect 7472 54432 7792 55456
rect 7472 54368 7480 54432
rect 7544 54368 7560 54432
rect 7624 54368 7640 54432
rect 7704 54368 7720 54432
rect 7784 54368 7792 54432
rect 7472 53344 7792 54368
rect 7472 53280 7480 53344
rect 7544 53280 7560 53344
rect 7624 53280 7640 53344
rect 7704 53280 7720 53344
rect 7784 53280 7792 53344
rect 7472 52256 7792 53280
rect 7472 52192 7480 52256
rect 7544 52192 7560 52256
rect 7624 52192 7640 52256
rect 7704 52192 7720 52256
rect 7784 52192 7792 52256
rect 7472 51168 7792 52192
rect 7472 51104 7480 51168
rect 7544 51104 7560 51168
rect 7624 51104 7640 51168
rect 7704 51104 7720 51168
rect 7784 51104 7792 51168
rect 7472 50080 7792 51104
rect 7472 50016 7480 50080
rect 7544 50016 7560 50080
rect 7624 50016 7640 50080
rect 7704 50016 7720 50080
rect 7784 50016 7792 50080
rect 7472 48992 7792 50016
rect 7472 48928 7480 48992
rect 7544 48928 7560 48992
rect 7624 48928 7640 48992
rect 7704 48928 7720 48992
rect 7784 48928 7792 48992
rect 7472 47904 7792 48928
rect 7472 47840 7480 47904
rect 7544 47840 7560 47904
rect 7624 47840 7640 47904
rect 7704 47840 7720 47904
rect 7784 47840 7792 47904
rect 6315 47564 6381 47565
rect 6315 47500 6316 47564
rect 6380 47500 6381 47564
rect 6315 47499 6381 47500
rect 5840 47296 5848 47360
rect 5912 47296 5928 47360
rect 5992 47296 6008 47360
rect 6072 47296 6088 47360
rect 6152 47296 6160 47360
rect 5579 47156 5645 47157
rect 5579 47092 5580 47156
rect 5644 47092 5645 47156
rect 5579 47091 5645 47092
rect 5395 42124 5461 42125
rect 5395 42060 5396 42124
rect 5460 42060 5461 42124
rect 5395 42059 5461 42060
rect 5395 41988 5461 41989
rect 5395 41924 5396 41988
rect 5460 41924 5461 41988
rect 5395 41923 5461 41924
rect 5211 41444 5277 41445
rect 5211 41380 5212 41444
rect 5276 41380 5277 41444
rect 5211 41379 5277 41380
rect 5211 41308 5277 41309
rect 5211 41244 5212 41308
rect 5276 41244 5277 41308
rect 5211 41243 5277 41244
rect 5027 36820 5093 36821
rect 5027 36756 5028 36820
rect 5092 36756 5093 36820
rect 5027 36755 5093 36756
rect 5027 36004 5093 36005
rect 5027 35940 5028 36004
rect 5092 35940 5093 36004
rect 5027 35939 5093 35940
rect 5030 28117 5090 35939
rect 5027 28116 5093 28117
rect 5027 28052 5028 28116
rect 5092 28052 5093 28116
rect 5027 28051 5093 28052
rect 5214 25941 5274 41243
rect 5398 39949 5458 41923
rect 5395 39948 5461 39949
rect 5395 39884 5396 39948
rect 5460 39884 5461 39948
rect 5395 39883 5461 39884
rect 5395 35732 5461 35733
rect 5395 35668 5396 35732
rect 5460 35668 5461 35732
rect 5395 35667 5461 35668
rect 5398 31109 5458 35667
rect 5395 31108 5461 31109
rect 5395 31044 5396 31108
rect 5460 31044 5461 31108
rect 5395 31043 5461 31044
rect 5211 25940 5277 25941
rect 5211 25876 5212 25940
rect 5276 25876 5277 25940
rect 5211 25875 5277 25876
rect 5582 15061 5642 47091
rect 5840 46272 6160 47296
rect 5840 46208 5848 46272
rect 5912 46208 5928 46272
rect 5992 46208 6008 46272
rect 6072 46208 6088 46272
rect 6152 46208 6160 46272
rect 5840 45184 6160 46208
rect 5840 45120 5848 45184
rect 5912 45120 5928 45184
rect 5992 45120 6008 45184
rect 6072 45120 6088 45184
rect 6152 45120 6160 45184
rect 5840 44096 6160 45120
rect 5840 44032 5848 44096
rect 5912 44032 5928 44096
rect 5992 44032 6008 44096
rect 6072 44032 6088 44096
rect 6152 44032 6160 44096
rect 5840 43008 6160 44032
rect 5840 42944 5848 43008
rect 5912 42944 5928 43008
rect 5992 42944 6008 43008
rect 6072 42944 6088 43008
rect 6152 42944 6160 43008
rect 5840 41920 6160 42944
rect 5840 41856 5848 41920
rect 5912 41856 5928 41920
rect 5992 41856 6008 41920
rect 6072 41856 6088 41920
rect 6152 41856 6160 41920
rect 5840 40832 6160 41856
rect 5840 40768 5848 40832
rect 5912 40768 5928 40832
rect 5992 40768 6008 40832
rect 6072 40768 6088 40832
rect 6152 40768 6160 40832
rect 5840 39744 6160 40768
rect 5840 39680 5848 39744
rect 5912 39680 5928 39744
rect 5992 39680 6008 39744
rect 6072 39680 6088 39744
rect 6152 39680 6160 39744
rect 5840 38656 6160 39680
rect 6318 38997 6378 47499
rect 7472 46816 7792 47840
rect 7472 46752 7480 46816
rect 7544 46752 7560 46816
rect 7624 46752 7640 46816
rect 7704 46752 7720 46816
rect 7784 46752 7792 46816
rect 6499 46476 6565 46477
rect 6499 46412 6500 46476
rect 6564 46412 6565 46476
rect 6499 46411 6565 46412
rect 6502 39541 6562 46411
rect 7472 45728 7792 46752
rect 9104 77824 9424 77840
rect 9104 77760 9112 77824
rect 9176 77760 9192 77824
rect 9256 77760 9272 77824
rect 9336 77760 9352 77824
rect 9416 77760 9424 77824
rect 9104 76736 9424 77760
rect 9104 76672 9112 76736
rect 9176 76672 9192 76736
rect 9256 76672 9272 76736
rect 9336 76672 9352 76736
rect 9416 76672 9424 76736
rect 9104 75648 9424 76672
rect 9104 75584 9112 75648
rect 9176 75584 9192 75648
rect 9256 75584 9272 75648
rect 9336 75584 9352 75648
rect 9416 75584 9424 75648
rect 9104 74560 9424 75584
rect 9104 74496 9112 74560
rect 9176 74496 9192 74560
rect 9256 74496 9272 74560
rect 9336 74496 9352 74560
rect 9416 74496 9424 74560
rect 9104 73472 9424 74496
rect 9104 73408 9112 73472
rect 9176 73408 9192 73472
rect 9256 73408 9272 73472
rect 9336 73408 9352 73472
rect 9416 73408 9424 73472
rect 9104 72384 9424 73408
rect 9104 72320 9112 72384
rect 9176 72320 9192 72384
rect 9256 72320 9272 72384
rect 9336 72320 9352 72384
rect 9416 72320 9424 72384
rect 9104 71296 9424 72320
rect 9104 71232 9112 71296
rect 9176 71232 9192 71296
rect 9256 71232 9272 71296
rect 9336 71232 9352 71296
rect 9416 71232 9424 71296
rect 9104 70208 9424 71232
rect 9104 70144 9112 70208
rect 9176 70144 9192 70208
rect 9256 70144 9272 70208
rect 9336 70144 9352 70208
rect 9416 70144 9424 70208
rect 9104 69120 9424 70144
rect 9104 69056 9112 69120
rect 9176 69056 9192 69120
rect 9256 69056 9272 69120
rect 9336 69056 9352 69120
rect 9416 69056 9424 69120
rect 9104 68032 9424 69056
rect 9104 67968 9112 68032
rect 9176 67968 9192 68032
rect 9256 67968 9272 68032
rect 9336 67968 9352 68032
rect 9416 67968 9424 68032
rect 9104 66944 9424 67968
rect 9104 66880 9112 66944
rect 9176 66880 9192 66944
rect 9256 66880 9272 66944
rect 9336 66880 9352 66944
rect 9416 66880 9424 66944
rect 9104 65856 9424 66880
rect 9104 65792 9112 65856
rect 9176 65792 9192 65856
rect 9256 65792 9272 65856
rect 9336 65792 9352 65856
rect 9416 65792 9424 65856
rect 9104 64768 9424 65792
rect 9104 64704 9112 64768
rect 9176 64704 9192 64768
rect 9256 64704 9272 64768
rect 9336 64704 9352 64768
rect 9416 64704 9424 64768
rect 9104 63680 9424 64704
rect 9104 63616 9112 63680
rect 9176 63616 9192 63680
rect 9256 63616 9272 63680
rect 9336 63616 9352 63680
rect 9416 63616 9424 63680
rect 9104 62592 9424 63616
rect 9104 62528 9112 62592
rect 9176 62528 9192 62592
rect 9256 62528 9272 62592
rect 9336 62528 9352 62592
rect 9416 62528 9424 62592
rect 9104 61504 9424 62528
rect 9104 61440 9112 61504
rect 9176 61440 9192 61504
rect 9256 61440 9272 61504
rect 9336 61440 9352 61504
rect 9416 61440 9424 61504
rect 9104 60416 9424 61440
rect 9104 60352 9112 60416
rect 9176 60352 9192 60416
rect 9256 60352 9272 60416
rect 9336 60352 9352 60416
rect 9416 60352 9424 60416
rect 9104 59328 9424 60352
rect 9104 59264 9112 59328
rect 9176 59264 9192 59328
rect 9256 59264 9272 59328
rect 9336 59264 9352 59328
rect 9416 59264 9424 59328
rect 9104 58240 9424 59264
rect 9104 58176 9112 58240
rect 9176 58176 9192 58240
rect 9256 58176 9272 58240
rect 9336 58176 9352 58240
rect 9416 58176 9424 58240
rect 9104 57152 9424 58176
rect 9104 57088 9112 57152
rect 9176 57088 9192 57152
rect 9256 57088 9272 57152
rect 9336 57088 9352 57152
rect 9416 57088 9424 57152
rect 9104 56064 9424 57088
rect 9104 56000 9112 56064
rect 9176 56000 9192 56064
rect 9256 56000 9272 56064
rect 9336 56000 9352 56064
rect 9416 56000 9424 56064
rect 9104 54976 9424 56000
rect 9104 54912 9112 54976
rect 9176 54912 9192 54976
rect 9256 54912 9272 54976
rect 9336 54912 9352 54976
rect 9416 54912 9424 54976
rect 9104 53888 9424 54912
rect 9104 53824 9112 53888
rect 9176 53824 9192 53888
rect 9256 53824 9272 53888
rect 9336 53824 9352 53888
rect 9416 53824 9424 53888
rect 9104 52800 9424 53824
rect 9104 52736 9112 52800
rect 9176 52736 9192 52800
rect 9256 52736 9272 52800
rect 9336 52736 9352 52800
rect 9416 52736 9424 52800
rect 9104 51712 9424 52736
rect 9104 51648 9112 51712
rect 9176 51648 9192 51712
rect 9256 51648 9272 51712
rect 9336 51648 9352 51712
rect 9416 51648 9424 51712
rect 9104 50624 9424 51648
rect 9104 50560 9112 50624
rect 9176 50560 9192 50624
rect 9256 50560 9272 50624
rect 9336 50560 9352 50624
rect 9416 50560 9424 50624
rect 9104 49536 9424 50560
rect 9104 49472 9112 49536
rect 9176 49472 9192 49536
rect 9256 49472 9272 49536
rect 9336 49472 9352 49536
rect 9416 49472 9424 49536
rect 9104 48448 9424 49472
rect 9104 48384 9112 48448
rect 9176 48384 9192 48448
rect 9256 48384 9272 48448
rect 9336 48384 9352 48448
rect 9416 48384 9424 48448
rect 9104 47360 9424 48384
rect 9104 47296 9112 47360
rect 9176 47296 9192 47360
rect 9256 47296 9272 47360
rect 9336 47296 9352 47360
rect 9416 47296 9424 47360
rect 8339 46612 8405 46613
rect 8339 46548 8340 46612
rect 8404 46548 8405 46612
rect 8339 46547 8405 46548
rect 7472 45664 7480 45728
rect 7544 45664 7560 45728
rect 7624 45664 7640 45728
rect 7704 45664 7720 45728
rect 7784 45664 7792 45728
rect 7472 44640 7792 45664
rect 7472 44576 7480 44640
rect 7544 44576 7560 44640
rect 7624 44576 7640 44640
rect 7704 44576 7720 44640
rect 7784 44576 7792 44640
rect 7472 43552 7792 44576
rect 7472 43488 7480 43552
rect 7544 43488 7560 43552
rect 7624 43488 7640 43552
rect 7704 43488 7720 43552
rect 7784 43488 7792 43552
rect 7472 42464 7792 43488
rect 7472 42400 7480 42464
rect 7544 42400 7560 42464
rect 7624 42400 7640 42464
rect 7704 42400 7720 42464
rect 7784 42400 7792 42464
rect 7472 41376 7792 42400
rect 7472 41312 7480 41376
rect 7544 41312 7560 41376
rect 7624 41312 7640 41376
rect 7704 41312 7720 41376
rect 7784 41312 7792 41376
rect 7472 40288 7792 41312
rect 7472 40224 7480 40288
rect 7544 40224 7560 40288
rect 7624 40224 7640 40288
rect 7704 40224 7720 40288
rect 7784 40224 7792 40288
rect 6499 39540 6565 39541
rect 6499 39476 6500 39540
rect 6564 39476 6565 39540
rect 6499 39475 6565 39476
rect 7472 39200 7792 40224
rect 7472 39136 7480 39200
rect 7544 39136 7560 39200
rect 7624 39136 7640 39200
rect 7704 39136 7720 39200
rect 7784 39136 7792 39200
rect 6315 38996 6381 38997
rect 6315 38932 6316 38996
rect 6380 38932 6381 38996
rect 6315 38931 6381 38932
rect 5840 38592 5848 38656
rect 5912 38592 5928 38656
rect 5992 38592 6008 38656
rect 6072 38592 6088 38656
rect 6152 38592 6160 38656
rect 5840 37568 6160 38592
rect 5840 37504 5848 37568
rect 5912 37504 5928 37568
rect 5992 37504 6008 37568
rect 6072 37504 6088 37568
rect 6152 37504 6160 37568
rect 5840 36480 6160 37504
rect 5840 36416 5848 36480
rect 5912 36416 5928 36480
rect 5992 36416 6008 36480
rect 6072 36416 6088 36480
rect 6152 36416 6160 36480
rect 5840 35392 6160 36416
rect 5840 35328 5848 35392
rect 5912 35328 5928 35392
rect 5992 35328 6008 35392
rect 6072 35328 6088 35392
rect 6152 35328 6160 35392
rect 5840 34304 6160 35328
rect 5840 34240 5848 34304
rect 5912 34240 5928 34304
rect 5992 34240 6008 34304
rect 6072 34240 6088 34304
rect 6152 34240 6160 34304
rect 5840 33216 6160 34240
rect 5840 33152 5848 33216
rect 5912 33152 5928 33216
rect 5992 33152 6008 33216
rect 6072 33152 6088 33216
rect 6152 33152 6160 33216
rect 5840 32128 6160 33152
rect 5840 32064 5848 32128
rect 5912 32064 5928 32128
rect 5992 32064 6008 32128
rect 6072 32064 6088 32128
rect 6152 32064 6160 32128
rect 5840 31040 6160 32064
rect 5840 30976 5848 31040
rect 5912 30976 5928 31040
rect 5992 30976 6008 31040
rect 6072 30976 6088 31040
rect 6152 30976 6160 31040
rect 5840 29952 6160 30976
rect 5840 29888 5848 29952
rect 5912 29888 5928 29952
rect 5992 29888 6008 29952
rect 6072 29888 6088 29952
rect 6152 29888 6160 29952
rect 5840 28864 6160 29888
rect 5840 28800 5848 28864
rect 5912 28800 5928 28864
rect 5992 28800 6008 28864
rect 6072 28800 6088 28864
rect 6152 28800 6160 28864
rect 5840 27776 6160 28800
rect 5840 27712 5848 27776
rect 5912 27712 5928 27776
rect 5992 27712 6008 27776
rect 6072 27712 6088 27776
rect 6152 27712 6160 27776
rect 5840 26688 6160 27712
rect 5840 26624 5848 26688
rect 5912 26624 5928 26688
rect 5992 26624 6008 26688
rect 6072 26624 6088 26688
rect 6152 26624 6160 26688
rect 5840 25600 6160 26624
rect 5840 25536 5848 25600
rect 5912 25536 5928 25600
rect 5992 25536 6008 25600
rect 6072 25536 6088 25600
rect 6152 25536 6160 25600
rect 5840 24512 6160 25536
rect 5840 24448 5848 24512
rect 5912 24448 5928 24512
rect 5992 24448 6008 24512
rect 6072 24448 6088 24512
rect 6152 24448 6160 24512
rect 5840 23424 6160 24448
rect 5840 23360 5848 23424
rect 5912 23360 5928 23424
rect 5992 23360 6008 23424
rect 6072 23360 6088 23424
rect 6152 23360 6160 23424
rect 5840 22336 6160 23360
rect 5840 22272 5848 22336
rect 5912 22272 5928 22336
rect 5992 22272 6008 22336
rect 6072 22272 6088 22336
rect 6152 22272 6160 22336
rect 5840 21248 6160 22272
rect 5840 21184 5848 21248
rect 5912 21184 5928 21248
rect 5992 21184 6008 21248
rect 6072 21184 6088 21248
rect 6152 21184 6160 21248
rect 5840 20160 6160 21184
rect 5840 20096 5848 20160
rect 5912 20096 5928 20160
rect 5992 20096 6008 20160
rect 6072 20096 6088 20160
rect 6152 20096 6160 20160
rect 5840 19072 6160 20096
rect 5840 19008 5848 19072
rect 5912 19008 5928 19072
rect 5992 19008 6008 19072
rect 6072 19008 6088 19072
rect 6152 19008 6160 19072
rect 5840 17984 6160 19008
rect 5840 17920 5848 17984
rect 5912 17920 5928 17984
rect 5992 17920 6008 17984
rect 6072 17920 6088 17984
rect 6152 17920 6160 17984
rect 5840 16896 6160 17920
rect 5840 16832 5848 16896
rect 5912 16832 5928 16896
rect 5992 16832 6008 16896
rect 6072 16832 6088 16896
rect 6152 16832 6160 16896
rect 5840 15808 6160 16832
rect 5840 15744 5848 15808
rect 5912 15744 5928 15808
rect 5992 15744 6008 15808
rect 6072 15744 6088 15808
rect 6152 15744 6160 15808
rect 5579 15060 5645 15061
rect 5579 14996 5580 15060
rect 5644 14996 5645 15060
rect 5579 14995 5645 14996
rect 5840 14720 6160 15744
rect 5840 14656 5848 14720
rect 5912 14656 5928 14720
rect 5992 14656 6008 14720
rect 6072 14656 6088 14720
rect 6152 14656 6160 14720
rect 5840 13632 6160 14656
rect 5840 13568 5848 13632
rect 5912 13568 5928 13632
rect 5992 13568 6008 13632
rect 6072 13568 6088 13632
rect 6152 13568 6160 13632
rect 5840 12544 6160 13568
rect 5840 12480 5848 12544
rect 5912 12480 5928 12544
rect 5992 12480 6008 12544
rect 6072 12480 6088 12544
rect 6152 12480 6160 12544
rect 5840 11456 6160 12480
rect 5840 11392 5848 11456
rect 5912 11392 5928 11456
rect 5992 11392 6008 11456
rect 6072 11392 6088 11456
rect 6152 11392 6160 11456
rect 5840 10368 6160 11392
rect 5840 10304 5848 10368
rect 5912 10304 5928 10368
rect 5992 10304 6008 10368
rect 6072 10304 6088 10368
rect 6152 10304 6160 10368
rect 4843 9484 4909 9485
rect 4843 9420 4844 9484
rect 4908 9420 4909 9484
rect 4843 9419 4909 9420
rect 5840 9280 6160 10304
rect 5840 9216 5848 9280
rect 5912 9216 5928 9280
rect 5992 9216 6008 9280
rect 6072 9216 6088 9280
rect 6152 9216 6160 9280
rect 5840 8192 6160 9216
rect 5840 8128 5848 8192
rect 5912 8128 5928 8192
rect 5992 8128 6008 8192
rect 6072 8128 6088 8192
rect 6152 8128 6160 8192
rect 5840 7104 6160 8128
rect 5840 7040 5848 7104
rect 5912 7040 5928 7104
rect 5992 7040 6008 7104
rect 6072 7040 6088 7104
rect 6152 7040 6160 7104
rect 5840 6016 6160 7040
rect 5840 5952 5848 6016
rect 5912 5952 5928 6016
rect 5992 5952 6008 6016
rect 6072 5952 6088 6016
rect 6152 5952 6160 6016
rect 5840 4928 6160 5952
rect 5840 4864 5848 4928
rect 5912 4864 5928 4928
rect 5992 4864 6008 4928
rect 6072 4864 6088 4928
rect 6152 4864 6160 4928
rect 4659 4860 4725 4861
rect 4659 4796 4660 4860
rect 4724 4796 4725 4860
rect 4659 4795 4725 4796
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 5840 3840 6160 4864
rect 5840 3776 5848 3840
rect 5912 3776 5928 3840
rect 5992 3776 6008 3840
rect 6072 3776 6088 3840
rect 6152 3776 6160 3840
rect 5840 2752 6160 3776
rect 5840 2688 5848 2752
rect 5912 2688 5928 2752
rect 5992 2688 6008 2752
rect 6072 2688 6088 2752
rect 6152 2688 6160 2752
rect 5840 2128 6160 2688
rect 7472 38112 7792 39136
rect 7472 38048 7480 38112
rect 7544 38048 7560 38112
rect 7624 38048 7640 38112
rect 7704 38048 7720 38112
rect 7784 38048 7792 38112
rect 7472 37024 7792 38048
rect 7472 36960 7480 37024
rect 7544 36960 7560 37024
rect 7624 36960 7640 37024
rect 7704 36960 7720 37024
rect 7784 36960 7792 37024
rect 7472 35936 7792 36960
rect 7472 35872 7480 35936
rect 7544 35872 7560 35936
rect 7624 35872 7640 35936
rect 7704 35872 7720 35936
rect 7784 35872 7792 35936
rect 7472 34848 7792 35872
rect 7472 34784 7480 34848
rect 7544 34784 7560 34848
rect 7624 34784 7640 34848
rect 7704 34784 7720 34848
rect 7784 34784 7792 34848
rect 7472 33760 7792 34784
rect 7472 33696 7480 33760
rect 7544 33696 7560 33760
rect 7624 33696 7640 33760
rect 7704 33696 7720 33760
rect 7784 33696 7792 33760
rect 7472 32672 7792 33696
rect 7472 32608 7480 32672
rect 7544 32608 7560 32672
rect 7624 32608 7640 32672
rect 7704 32608 7720 32672
rect 7784 32608 7792 32672
rect 7472 31584 7792 32608
rect 7472 31520 7480 31584
rect 7544 31520 7560 31584
rect 7624 31520 7640 31584
rect 7704 31520 7720 31584
rect 7784 31520 7792 31584
rect 7472 30496 7792 31520
rect 7472 30432 7480 30496
rect 7544 30432 7560 30496
rect 7624 30432 7640 30496
rect 7704 30432 7720 30496
rect 7784 30432 7792 30496
rect 7472 29408 7792 30432
rect 7472 29344 7480 29408
rect 7544 29344 7560 29408
rect 7624 29344 7640 29408
rect 7704 29344 7720 29408
rect 7784 29344 7792 29408
rect 7472 28320 7792 29344
rect 7472 28256 7480 28320
rect 7544 28256 7560 28320
rect 7624 28256 7640 28320
rect 7704 28256 7720 28320
rect 7784 28256 7792 28320
rect 7472 27232 7792 28256
rect 7472 27168 7480 27232
rect 7544 27168 7560 27232
rect 7624 27168 7640 27232
rect 7704 27168 7720 27232
rect 7784 27168 7792 27232
rect 7472 26144 7792 27168
rect 7472 26080 7480 26144
rect 7544 26080 7560 26144
rect 7624 26080 7640 26144
rect 7704 26080 7720 26144
rect 7784 26080 7792 26144
rect 7472 25056 7792 26080
rect 7472 24992 7480 25056
rect 7544 24992 7560 25056
rect 7624 24992 7640 25056
rect 7704 24992 7720 25056
rect 7784 24992 7792 25056
rect 7472 23968 7792 24992
rect 7472 23904 7480 23968
rect 7544 23904 7560 23968
rect 7624 23904 7640 23968
rect 7704 23904 7720 23968
rect 7784 23904 7792 23968
rect 7472 22880 7792 23904
rect 7472 22816 7480 22880
rect 7544 22816 7560 22880
rect 7624 22816 7640 22880
rect 7704 22816 7720 22880
rect 7784 22816 7792 22880
rect 7472 21792 7792 22816
rect 7472 21728 7480 21792
rect 7544 21728 7560 21792
rect 7624 21728 7640 21792
rect 7704 21728 7720 21792
rect 7784 21728 7792 21792
rect 7472 20704 7792 21728
rect 7472 20640 7480 20704
rect 7544 20640 7560 20704
rect 7624 20640 7640 20704
rect 7704 20640 7720 20704
rect 7784 20640 7792 20704
rect 7472 19616 7792 20640
rect 7472 19552 7480 19616
rect 7544 19552 7560 19616
rect 7624 19552 7640 19616
rect 7704 19552 7720 19616
rect 7784 19552 7792 19616
rect 7472 18528 7792 19552
rect 7472 18464 7480 18528
rect 7544 18464 7560 18528
rect 7624 18464 7640 18528
rect 7704 18464 7720 18528
rect 7784 18464 7792 18528
rect 7472 17440 7792 18464
rect 7472 17376 7480 17440
rect 7544 17376 7560 17440
rect 7624 17376 7640 17440
rect 7704 17376 7720 17440
rect 7784 17376 7792 17440
rect 7472 16352 7792 17376
rect 7472 16288 7480 16352
rect 7544 16288 7560 16352
rect 7624 16288 7640 16352
rect 7704 16288 7720 16352
rect 7784 16288 7792 16352
rect 7472 15264 7792 16288
rect 7472 15200 7480 15264
rect 7544 15200 7560 15264
rect 7624 15200 7640 15264
rect 7704 15200 7720 15264
rect 7784 15200 7792 15264
rect 7472 14176 7792 15200
rect 7472 14112 7480 14176
rect 7544 14112 7560 14176
rect 7624 14112 7640 14176
rect 7704 14112 7720 14176
rect 7784 14112 7792 14176
rect 7472 13088 7792 14112
rect 7472 13024 7480 13088
rect 7544 13024 7560 13088
rect 7624 13024 7640 13088
rect 7704 13024 7720 13088
rect 7784 13024 7792 13088
rect 7472 12000 7792 13024
rect 7472 11936 7480 12000
rect 7544 11936 7560 12000
rect 7624 11936 7640 12000
rect 7704 11936 7720 12000
rect 7784 11936 7792 12000
rect 7472 10912 7792 11936
rect 7472 10848 7480 10912
rect 7544 10848 7560 10912
rect 7624 10848 7640 10912
rect 7704 10848 7720 10912
rect 7784 10848 7792 10912
rect 7472 9824 7792 10848
rect 7472 9760 7480 9824
rect 7544 9760 7560 9824
rect 7624 9760 7640 9824
rect 7704 9760 7720 9824
rect 7784 9760 7792 9824
rect 7472 8736 7792 9760
rect 7472 8672 7480 8736
rect 7544 8672 7560 8736
rect 7624 8672 7640 8736
rect 7704 8672 7720 8736
rect 7784 8672 7792 8736
rect 7472 7648 7792 8672
rect 7472 7584 7480 7648
rect 7544 7584 7560 7648
rect 7624 7584 7640 7648
rect 7704 7584 7720 7648
rect 7784 7584 7792 7648
rect 7472 6560 7792 7584
rect 7472 6496 7480 6560
rect 7544 6496 7560 6560
rect 7624 6496 7640 6560
rect 7704 6496 7720 6560
rect 7784 6496 7792 6560
rect 7472 5472 7792 6496
rect 7472 5408 7480 5472
rect 7544 5408 7560 5472
rect 7624 5408 7640 5472
rect 7704 5408 7720 5472
rect 7784 5408 7792 5472
rect 7472 4384 7792 5408
rect 8342 5269 8402 46547
rect 9104 46272 9424 47296
rect 9104 46208 9112 46272
rect 9176 46208 9192 46272
rect 9256 46208 9272 46272
rect 9336 46208 9352 46272
rect 9416 46208 9424 46272
rect 9104 45184 9424 46208
rect 9104 45120 9112 45184
rect 9176 45120 9192 45184
rect 9256 45120 9272 45184
rect 9336 45120 9352 45184
rect 9416 45120 9424 45184
rect 9104 44096 9424 45120
rect 9104 44032 9112 44096
rect 9176 44032 9192 44096
rect 9256 44032 9272 44096
rect 9336 44032 9352 44096
rect 9416 44032 9424 44096
rect 9104 43008 9424 44032
rect 9104 42944 9112 43008
rect 9176 42944 9192 43008
rect 9256 42944 9272 43008
rect 9336 42944 9352 43008
rect 9416 42944 9424 43008
rect 9104 41920 9424 42944
rect 9104 41856 9112 41920
rect 9176 41856 9192 41920
rect 9256 41856 9272 41920
rect 9336 41856 9352 41920
rect 9416 41856 9424 41920
rect 9104 40832 9424 41856
rect 9104 40768 9112 40832
rect 9176 40768 9192 40832
rect 9256 40768 9272 40832
rect 9336 40768 9352 40832
rect 9416 40768 9424 40832
rect 9104 39744 9424 40768
rect 9104 39680 9112 39744
rect 9176 39680 9192 39744
rect 9256 39680 9272 39744
rect 9336 39680 9352 39744
rect 9416 39680 9424 39744
rect 9104 38656 9424 39680
rect 9104 38592 9112 38656
rect 9176 38592 9192 38656
rect 9256 38592 9272 38656
rect 9336 38592 9352 38656
rect 9416 38592 9424 38656
rect 9104 37568 9424 38592
rect 9104 37504 9112 37568
rect 9176 37504 9192 37568
rect 9256 37504 9272 37568
rect 9336 37504 9352 37568
rect 9416 37504 9424 37568
rect 9104 36480 9424 37504
rect 9104 36416 9112 36480
rect 9176 36416 9192 36480
rect 9256 36416 9272 36480
rect 9336 36416 9352 36480
rect 9416 36416 9424 36480
rect 9104 35392 9424 36416
rect 9104 35328 9112 35392
rect 9176 35328 9192 35392
rect 9256 35328 9272 35392
rect 9336 35328 9352 35392
rect 9416 35328 9424 35392
rect 9104 34304 9424 35328
rect 9104 34240 9112 34304
rect 9176 34240 9192 34304
rect 9256 34240 9272 34304
rect 9336 34240 9352 34304
rect 9416 34240 9424 34304
rect 9104 33216 9424 34240
rect 9104 33152 9112 33216
rect 9176 33152 9192 33216
rect 9256 33152 9272 33216
rect 9336 33152 9352 33216
rect 9416 33152 9424 33216
rect 9104 32128 9424 33152
rect 9104 32064 9112 32128
rect 9176 32064 9192 32128
rect 9256 32064 9272 32128
rect 9336 32064 9352 32128
rect 9416 32064 9424 32128
rect 9104 31040 9424 32064
rect 9104 30976 9112 31040
rect 9176 30976 9192 31040
rect 9256 30976 9272 31040
rect 9336 30976 9352 31040
rect 9416 30976 9424 31040
rect 9104 29952 9424 30976
rect 9104 29888 9112 29952
rect 9176 29888 9192 29952
rect 9256 29888 9272 29952
rect 9336 29888 9352 29952
rect 9416 29888 9424 29952
rect 9104 28864 9424 29888
rect 9104 28800 9112 28864
rect 9176 28800 9192 28864
rect 9256 28800 9272 28864
rect 9336 28800 9352 28864
rect 9416 28800 9424 28864
rect 9104 27776 9424 28800
rect 9104 27712 9112 27776
rect 9176 27712 9192 27776
rect 9256 27712 9272 27776
rect 9336 27712 9352 27776
rect 9416 27712 9424 27776
rect 9104 26688 9424 27712
rect 9104 26624 9112 26688
rect 9176 26624 9192 26688
rect 9256 26624 9272 26688
rect 9336 26624 9352 26688
rect 9416 26624 9424 26688
rect 9104 25600 9424 26624
rect 9104 25536 9112 25600
rect 9176 25536 9192 25600
rect 9256 25536 9272 25600
rect 9336 25536 9352 25600
rect 9416 25536 9424 25600
rect 9104 24512 9424 25536
rect 9104 24448 9112 24512
rect 9176 24448 9192 24512
rect 9256 24448 9272 24512
rect 9336 24448 9352 24512
rect 9416 24448 9424 24512
rect 9104 23424 9424 24448
rect 9104 23360 9112 23424
rect 9176 23360 9192 23424
rect 9256 23360 9272 23424
rect 9336 23360 9352 23424
rect 9416 23360 9424 23424
rect 9104 22336 9424 23360
rect 9104 22272 9112 22336
rect 9176 22272 9192 22336
rect 9256 22272 9272 22336
rect 9336 22272 9352 22336
rect 9416 22272 9424 22336
rect 9104 21248 9424 22272
rect 9104 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9272 21248
rect 9336 21184 9352 21248
rect 9416 21184 9424 21248
rect 9104 20160 9424 21184
rect 9104 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9272 20160
rect 9336 20096 9352 20160
rect 9416 20096 9424 20160
rect 9104 19072 9424 20096
rect 9104 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9272 19072
rect 9336 19008 9352 19072
rect 9416 19008 9424 19072
rect 9104 17984 9424 19008
rect 9104 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9272 17984
rect 9336 17920 9352 17984
rect 9416 17920 9424 17984
rect 9104 16896 9424 17920
rect 9104 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9272 16896
rect 9336 16832 9352 16896
rect 9416 16832 9424 16896
rect 9104 15808 9424 16832
rect 9104 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9272 15808
rect 9336 15744 9352 15808
rect 9416 15744 9424 15808
rect 9104 14720 9424 15744
rect 9104 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9272 14720
rect 9336 14656 9352 14720
rect 9416 14656 9424 14720
rect 9104 13632 9424 14656
rect 9104 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9272 13632
rect 9336 13568 9352 13632
rect 9416 13568 9424 13632
rect 9104 12544 9424 13568
rect 9104 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9272 12544
rect 9336 12480 9352 12544
rect 9416 12480 9424 12544
rect 9104 11456 9424 12480
rect 9104 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9272 11456
rect 9336 11392 9352 11456
rect 9416 11392 9424 11456
rect 9104 10368 9424 11392
rect 9104 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9272 10368
rect 9336 10304 9352 10368
rect 9416 10304 9424 10368
rect 9104 9280 9424 10304
rect 9104 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9272 9280
rect 9336 9216 9352 9280
rect 9416 9216 9424 9280
rect 9104 8192 9424 9216
rect 9104 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9272 8192
rect 9336 8128 9352 8192
rect 9416 8128 9424 8192
rect 9104 7104 9424 8128
rect 9104 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9272 7104
rect 9336 7040 9352 7104
rect 9416 7040 9424 7104
rect 9104 6016 9424 7040
rect 9104 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9272 6016
rect 9336 5952 9352 6016
rect 9416 5952 9424 6016
rect 8339 5268 8405 5269
rect 8339 5204 8340 5268
rect 8404 5204 8405 5268
rect 8339 5203 8405 5204
rect 7472 4320 7480 4384
rect 7544 4320 7560 4384
rect 7624 4320 7640 4384
rect 7704 4320 7720 4384
rect 7784 4320 7792 4384
rect 7472 3296 7792 4320
rect 7472 3232 7480 3296
rect 7544 3232 7560 3296
rect 7624 3232 7640 3296
rect 7704 3232 7720 3296
rect 7784 3232 7792 3296
rect 7472 2208 7792 3232
rect 7472 2144 7480 2208
rect 7544 2144 7560 2208
rect 7624 2144 7640 2208
rect 7704 2144 7720 2208
rect 7784 2144 7792 2208
rect 7472 2128 7792 2144
rect 9104 4928 9424 5952
rect 9104 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9272 4928
rect 9336 4864 9352 4928
rect 9416 4864 9424 4928
rect 9104 3840 9424 4864
rect 9104 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9272 3840
rect 9336 3776 9352 3840
rect 9416 3776 9424 3840
rect 9104 2752 9424 3776
rect 9104 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9272 2752
rect 9336 2688 9352 2752
rect 9416 2688 9424 2752
rect 9104 2128 9424 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 2300 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39
timestamp 1644511149
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46
timestamp 1644511149
transform 1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91
timestamp 1644511149
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_14
timestamp 1644511149
transform 1 0 2392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1644511149
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1644511149
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1644511149
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_91
timestamp 1644511149
transform 1 0 9476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_99
timestamp 1644511149
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_34
timestamp 1644511149
transform 1 0 4232 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_46
timestamp 1644511149
transform 1 0 5336 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_58
timestamp 1644511149
transform 1 0 6440 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_70
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1644511149
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1644511149
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1644511149
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_22
timestamp 1644511149
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_31
timestamp 1644511149
transform 1 0 3956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_38
timestamp 1644511149
transform 1 0 4600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_45
timestamp 1644511149
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1644511149
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1644511149
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_11
timestamp 1644511149
transform 1 0 2116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_17
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1644511149
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_33
timestamp 1644511149
transform 1 0 4140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_40
timestamp 1644511149
transform 1 0 4784 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_52
timestamp 1644511149
transform 1 0 5888 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_64
timestamp 1644511149
transform 1 0 6992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1644511149
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1644511149
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_99
timestamp 1644511149
transform 1 0 10212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1644511149
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_22
timestamp 1644511149
transform 1 0 3128 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_30
timestamp 1644511149
transform 1 0 3864 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_42
timestamp 1644511149
transform 1 0 4968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1644511149
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 1644511149
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_91
timestamp 1644511149
transform 1 0 9476 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1644511149
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1644511149
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 1644511149
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_34
timestamp 1644511149
transform 1 0 4232 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_46
timestamp 1644511149
transform 1 0 5336 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_58
timestamp 1644511149
transform 1 0 6440 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_70
timestamp 1644511149
transform 1 0 7544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1644511149
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1644511149
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1644511149
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_11
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_18
timestamp 1644511149
transform 1 0 2760 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_25
timestamp 1644511149
transform 1 0 3404 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_37
timestamp 1644511149
transform 1 0 4508 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp 1644511149
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1644511149
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1644511149
transform 1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1644511149
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1644511149
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_99
timestamp 1644511149
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_33
timestamp 1644511149
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1644511149
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1644511149
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1644511149
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1644511149
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1644511149
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_13
timestamp 1644511149
transform 1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_22
timestamp 1644511149
transform 1 0 3128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_29
timestamp 1644511149
transform 1 0 3772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_41
timestamp 1644511149
transform 1 0 4876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1644511149
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1644511149
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1644511149
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1644511149
transform 1 0 4048 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1644511149
transform 1 0 5152 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1644511149
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1644511149
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1644511149
transform 1 0 9660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_99
timestamp 1644511149
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1644511149
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1644511149
transform 1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_28
timestamp 1644511149
transform 1 0 3680 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_40
timestamp 1644511149
transform 1 0 4784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1644511149
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_99
timestamp 1644511149
transform 1 0 10212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1644511149
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1644511149
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1644511149
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1644511149
transform 1 0 3036 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_28
timestamp 1644511149
transform 1 0 3680 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_40
timestamp 1644511149
transform 1 0 4784 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1644511149
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1644511149
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp 1644511149
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1644511149
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1644511149
transform 1 0 4048 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1644511149
transform 1 0 5152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1644511149
transform 1 0 6256 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1644511149
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1644511149
transform 1 0 9660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_99
timestamp 1644511149
transform 1 0 10212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1644511149
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1644511149
transform 1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_28
timestamp 1644511149
transform 1 0 3680 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_40
timestamp 1644511149
transform 1 0 4784 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1644511149
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1644511149
transform 1 0 10396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_9
timestamp 1644511149
transform 1 0 1932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_17
timestamp 1644511149
transform 1 0 2668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1644511149
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_91
timestamp 1644511149
transform 1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_99
timestamp 1644511149
transform 1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_6
timestamp 1644511149
transform 1 0 1656 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_21
timestamp 1644511149
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_33
timestamp 1644511149
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1644511149
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1644511149
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_87
timestamp 1644511149
transform 1 0 9108 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_91
timestamp 1644511149
transform 1 0 9476 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1644511149
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_6
timestamp 1644511149
transform 1 0 1656 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_17
timestamp 1644511149
transform 1 0 2668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1644511149
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1644511149
transform 1 0 4048 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1644511149
transform 1 0 5152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1644511149
transform 1 0 6256 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1644511149
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_92
timestamp 1644511149
transform 1 0 9568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99
timestamp 1644511149
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_6
timestamp 1644511149
transform 1 0 1656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_24
timestamp 1644511149
transform 1 0 3312 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1644511149
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_43
timestamp 1644511149
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1644511149
transform 1 0 10212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_9
timestamp 1644511149
transform 1 0 1932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1644511149
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1644511149
transform 1 0 4048 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1644511149
transform 1 0 5152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1644511149
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1644511149
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1644511149
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1644511149
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1644511149
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_13
timestamp 1644511149
transform 1 0 2300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_21
timestamp 1644511149
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_33
timestamp 1644511149
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1644511149
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1644511149
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_99
timestamp 1644511149
transform 1 0 10212 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_13
timestamp 1644511149
transform 1 0 2300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1644511149
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1644511149
transform 1 0 4048 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1644511149
transform 1 0 5152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1644511149
transform 1 0 6256 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1644511149
transform 1 0 7360 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1644511149
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1644511149
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_99
timestamp 1644511149
transform 1 0 10212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_12
timestamp 1644511149
transform 1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_20
timestamp 1644511149
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_32
timestamp 1644511149
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_44
timestamp 1644511149
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 1644511149
transform 1 0 9108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_91
timestamp 1644511149
transform 1 0 9476 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1644511149
transform 1 0 10212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 1644511149
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1644511149
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1644511149
transform 1 0 4048 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1644511149
transform 1 0 5152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1644511149
transform 1 0 6256 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1644511149
transform 1 0 7360 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1644511149
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1644511149
transform 1 0 10212 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_6
timestamp 1644511149
transform 1 0 1656 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_14
timestamp 1644511149
transform 1 0 2392 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_22
timestamp 1644511149
transform 1 0 3128 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_34
timestamp 1644511149
transform 1 0 4232 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_46
timestamp 1644511149
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1644511149
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_99
timestamp 1644511149
transform 1 0 10212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_6
timestamp 1644511149
transform 1 0 1656 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_10
timestamp 1644511149
transform 1 0 2024 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1644511149
transform 1 0 5152 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1644511149
transform 1 0 6256 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1644511149
transform 1 0 7360 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1644511149
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1644511149
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_99
timestamp 1644511149
transform 1 0 10212 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_6
timestamp 1644511149
transform 1 0 1656 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_12
timestamp 1644511149
transform 1 0 2208 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_18
timestamp 1644511149
transform 1 0 2760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_30
timestamp 1644511149
transform 1 0 3864 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_42
timestamp 1644511149
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1644511149
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_87
timestamp 1644511149
transform 1 0 9108 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_91
timestamp 1644511149
transform 1 0 9476 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_99
timestamp 1644511149
transform 1 0 10212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_6
timestamp 1644511149
transform 1 0 1656 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_13
timestamp 1644511149
transform 1 0 2300 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 1644511149
transform 1 0 2944 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1644511149
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_99
timestamp 1644511149
transform 1 0 10212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_11
timestamp 1644511149
transform 1 0 2116 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_18
timestamp 1644511149
transform 1 0 2760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_30
timestamp 1644511149
transform 1 0 3864 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_42
timestamp 1644511149
transform 1 0 4968 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1644511149
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_98
timestamp 1644511149
transform 1 0 10120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_102
timestamp 1644511149
transform 1 0 10488 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_12
timestamp 1644511149
transform 1 0 2208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1644511149
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1644511149
transform 1 0 4048 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1644511149
transform 1 0 5152 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1644511149
transform 1 0 6256 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1644511149
transform 1 0 7360 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1644511149
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1644511149
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1644511149
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_13
timestamp 1644511149
transform 1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_22
timestamp 1644511149
transform 1 0 3128 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_34
timestamp 1644511149
transform 1 0 4232 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 1644511149
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1644511149
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_99
timestamp 1644511149
transform 1 0 10212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_13
timestamp 1644511149
transform 1 0 2300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1644511149
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_13
timestamp 1644511149
transform 1 0 2300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_23
timestamp 1644511149
transform 1 0 3220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1644511149
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1644511149
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_99
timestamp 1644511149
transform 1 0 10212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1644511149
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_22
timestamp 1644511149
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_34
timestamp 1644511149
transform 1 0 4232 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_46
timestamp 1644511149
transform 1 0 5336 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_58
timestamp 1644511149
transform 1 0 6440 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_70
timestamp 1644511149
transform 1 0 7544 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1644511149
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_93
timestamp 1644511149
transform 1 0 9660 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1644511149
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_13
timestamp 1644511149
transform 1 0 2300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_22
timestamp 1644511149
transform 1 0 3128 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_30
timestamp 1644511149
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_38
timestamp 1644511149
transform 1 0 4600 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_50
timestamp 1644511149
transform 1 0 5704 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_99
timestamp 1644511149
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_13
timestamp 1644511149
transform 1 0 2300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1644511149
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_13
timestamp 1644511149
transform 1 0 2300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_99
timestamp 1644511149
transform 1 0 10212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_13
timestamp 1644511149
transform 1 0 2300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1644511149
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_93
timestamp 1644511149
transform 1 0 9660 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1644511149
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_11
timestamp 1644511149
transform 1 0 2116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_19
timestamp 1644511149
transform 1 0 2852 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_101
timestamp 1644511149
transform 1 0 10396 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_13
timestamp 1644511149
transform 1 0 2300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_17
timestamp 1644511149
transform 1 0 2668 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_23
timestamp 1644511149
transform 1 0 3220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_93
timestamp 1644511149
transform 1 0 9660 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1644511149
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_13
timestamp 1644511149
transform 1 0 2300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_22
timestamp 1644511149
transform 1 0 3128 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_34
timestamp 1644511149
transform 1 0 4232 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_46
timestamp 1644511149
transform 1 0 5336 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1644511149
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_99
timestamp 1644511149
transform 1 0 10212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_11
timestamp 1644511149
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1644511149
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_37
timestamp 1644511149
transform 1 0 4508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_49
timestamp 1644511149
transform 1 0 5612 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_61
timestamp 1644511149
transform 1 0 6716 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_73
timestamp 1644511149
transform 1 0 7820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1644511149
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_7
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_13
timestamp 1644511149
transform 1 0 2300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_22
timestamp 1644511149
transform 1 0 3128 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_30
timestamp 1644511149
transform 1 0 3864 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_42
timestamp 1644511149
transform 1 0 4968 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1644511149
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_99
timestamp 1644511149
transform 1 0 10212 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_13
timestamp 1644511149
transform 1 0 2300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_22
timestamp 1644511149
transform 1 0 3128 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_37
timestamp 1644511149
transform 1 0 4508 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_49
timestamp 1644511149
transform 1 0 5612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_61
timestamp 1644511149
transform 1 0 6716 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_73
timestamp 1644511149
transform 1 0 7820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1644511149
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_93
timestamp 1644511149
transform 1 0 9660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_99
timestamp 1644511149
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_13
timestamp 1644511149
transform 1 0 2300 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_22
timestamp 1644511149
transform 1 0 3128 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_30
timestamp 1644511149
transform 1 0 3864 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_37
timestamp 1644511149
transform 1 0 4508 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_49
timestamp 1644511149
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_99
timestamp 1644511149
transform 1 0 10212 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_11
timestamp 1644511149
transform 1 0 2116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1644511149
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_33
timestamp 1644511149
transform 1 0 4140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_45
timestamp 1644511149
transform 1 0 5244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_57
timestamp 1644511149
transform 1 0 6348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_69
timestamp 1644511149
transform 1 0 7452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_81
timestamp 1644511149
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_13
timestamp 1644511149
transform 1 0 2300 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_21
timestamp 1644511149
transform 1 0 3036 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_33
timestamp 1644511149
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1644511149
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1644511149
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_99
timestamp 1644511149
transform 1 0 10212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_11
timestamp 1644511149
transform 1 0 2116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1644511149
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_74
timestamp 1644511149
transform 1 0 7912 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1644511149
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_93
timestamp 1644511149
transform 1 0 9660 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_99
timestamp 1644511149
transform 1 0 10212 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_9
timestamp 1644511149
transform 1 0 1932 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_18
timestamp 1644511149
transform 1 0 2760 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_26
timestamp 1644511149
transform 1 0 3496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_33
timestamp 1644511149
transform 1 0 4140 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_40
timestamp 1644511149
transform 1 0 4784 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1644511149
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_101
timestamp 1644511149
transform 1 0 10396 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_11
timestamp 1644511149
transform 1 0 2116 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_19
timestamp 1644511149
transform 1 0 2852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_93
timestamp 1644511149
transform 1 0 9660 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_99
timestamp 1644511149
transform 1 0 10212 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_10
timestamp 1644511149
transform 1 0 2024 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_16
timestamp 1644511149
transform 1 0 2576 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_22
timestamp 1644511149
transform 1 0 3128 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_31
timestamp 1644511149
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_43
timestamp 1644511149
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_99
timestamp 1644511149
transform 1 0 10212 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_11
timestamp 1644511149
transform 1 0 2116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 1644511149
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_33
timestamp 1644511149
transform 1 0 4140 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_40
timestamp 1644511149
transform 1 0 4784 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_52
timestamp 1644511149
transform 1 0 5888 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_64
timestamp 1644511149
transform 1 0 6992 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_76
timestamp 1644511149
transform 1 0 8096 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_93
timestamp 1644511149
transform 1 0 9660 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_99
timestamp 1644511149
transform 1 0 10212 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_9
timestamp 1644511149
transform 1 0 1932 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_23
timestamp 1644511149
transform 1 0 3220 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_30
timestamp 1644511149
transform 1 0 3864 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_37
timestamp 1644511149
transform 1 0 4508 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_49
timestamp 1644511149
transform 1 0 5612 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_101
timestamp 1644511149
transform 1 0 10396 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_23
timestamp 1644511149
transform 1 0 3220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1644511149
transform 1 0 4048 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1644511149
transform 1 0 5152 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1644511149
transform 1 0 6256 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_68
timestamp 1644511149
transform 1 0 7360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1644511149
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_93
timestamp 1644511149
transform 1 0 9660 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_99
timestamp 1644511149
transform 1 0 10212 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_7
timestamp 1644511149
transform 1 0 1748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_21
timestamp 1644511149
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_38
timestamp 1644511149
transform 1 0 4600 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_50
timestamp 1644511149
transform 1 0 5704 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_99
timestamp 1644511149
transform 1 0 10212 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_11
timestamp 1644511149
transform 1 0 2116 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_22
timestamp 1644511149
transform 1 0 3128 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_32
timestamp 1644511149
transform 1 0 4048 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_44
timestamp 1644511149
transform 1 0 5152 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_56
timestamp 1644511149
transform 1 0 6256 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_68
timestamp 1644511149
transform 1 0 7360 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_80
timestamp 1644511149
transform 1 0 8464 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_93
timestamp 1644511149
transform 1 0 9660 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_99
timestamp 1644511149
transform 1 0 10212 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_7
timestamp 1644511149
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_23
timestamp 1644511149
transform 1 0 3220 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_36
timestamp 1644511149
transform 1 0 4416 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_48
timestamp 1644511149
transform 1 0 5520 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_99
timestamp 1644511149
transform 1 0 10212 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_10
timestamp 1644511149
transform 1 0 2024 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_18
timestamp 1644511149
transform 1 0 2760 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1644511149
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_42
timestamp 1644511149
transform 1 0 4968 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_54
timestamp 1644511149
transform 1 0 6072 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_66
timestamp 1644511149
transform 1 0 7176 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_78
timestamp 1644511149
transform 1 0 8280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_93
timestamp 1644511149
transform 1 0 9660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_99
timestamp 1644511149
transform 1 0 10212 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_7
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_33
timestamp 1644511149
transform 1 0 4140 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_37
timestamp 1644511149
transform 1 0 4508 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_43
timestamp 1644511149
transform 1 0 5060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_99
timestamp 1644511149
transform 1 0 10212 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_14
timestamp 1644511149
transform 1 0 2392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_22
timestamp 1644511149
transform 1 0 3128 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_91
timestamp 1644511149
transform 1 0 9476 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_99
timestamp 1644511149
transform 1 0 10212 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_10
timestamp 1644511149
transform 1 0 2024 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_17
timestamp 1644511149
transform 1 0 2668 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_21
timestamp 1644511149
transform 1 0 3036 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_33
timestamp 1644511149
transform 1 0 4140 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_99
timestamp 1644511149
transform 1 0 10212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_22
timestamp 1644511149
transform 1 0 3128 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_33
timestamp 1644511149
transform 1 0 4140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_45
timestamp 1644511149
transform 1 0 5244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_69
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1644511149
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_93
timestamp 1644511149
transform 1 0 9660 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_99
timestamp 1644511149
transform 1 0 10212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_10
timestamp 1644511149
transform 1 0 2024 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_19
timestamp 1644511149
transform 1 0 2852 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_35
timestamp 1644511149
transform 1 0 4324 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_47
timestamp 1644511149
transform 1 0 5428 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_99
timestamp 1644511149
transform 1 0 10212 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_7
timestamp 1644511149
transform 1 0 1748 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_20
timestamp 1644511149
transform 1 0 2944 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_33
timestamp 1644511149
transform 1 0 4140 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_39
timestamp 1644511149
transform 1 0 4692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_51
timestamp 1644511149
transform 1 0 5796 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_63
timestamp 1644511149
transform 1 0 6900 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_75
timestamp 1644511149
transform 1 0 8004 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_93
timestamp 1644511149
transform 1 0 9660 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_99
timestamp 1644511149
transform 1 0 10212 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_14
timestamp 1644511149
transform 1 0 2392 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_28
timestamp 1644511149
transform 1 0 3680 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_36
timestamp 1644511149
transform 1 0 4416 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_44
timestamp 1644511149
transform 1 0 5152 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_99
timestamp 1644511149
transform 1 0 10212 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_14
timestamp 1644511149
transform 1 0 2392 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_23
timestamp 1644511149
transform 1 0 3220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_34
timestamp 1644511149
transform 1 0 4232 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_42
timestamp 1644511149
transform 1 0 4968 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_49
timestamp 1644511149
transform 1 0 5612 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_61
timestamp 1644511149
transform 1 0 6716 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_73
timestamp 1644511149
transform 1 0 7820 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_81
timestamp 1644511149
transform 1 0 8556 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_93
timestamp 1644511149
transform 1 0 9660 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_99
timestamp 1644511149
transform 1 0 10212 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_10
timestamp 1644511149
transform 1 0 2024 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_24
timestamp 1644511149
transform 1 0 3312 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_32
timestamp 1644511149
transform 1 0 4048 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_40
timestamp 1644511149
transform 1 0 4784 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_52
timestamp 1644511149
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_60
timestamp 1644511149
transform 1 0 6624 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_72
timestamp 1644511149
transform 1 0 7728 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_84
timestamp 1644511149
transform 1 0 8832 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_92
timestamp 1644511149
transform 1 0 9568 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_99
timestamp 1644511149
transform 1 0 10212 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_9
timestamp 1644511149
transform 1 0 1932 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_20
timestamp 1644511149
transform 1 0 2944 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_33
timestamp 1644511149
transform 1 0 4140 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_45
timestamp 1644511149
transform 1 0 5244 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_57
timestamp 1644511149
transform 1 0 6348 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_69
timestamp 1644511149
transform 1 0 7452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_81
timestamp 1644511149
transform 1 0 8556 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_91
timestamp 1644511149
transform 1 0 9476 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_99
timestamp 1644511149
transform 1 0 10212 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_10
timestamp 1644511149
transform 1 0 2024 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_19
timestamp 1644511149
transform 1 0 2852 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_40
timestamp 1644511149
transform 1 0 4784 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_99
timestamp 1644511149
transform 1 0 10212 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_17
timestamp 1644511149
transform 1 0 2668 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_25
timestamp 1644511149
transform 1 0 3404 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_33
timestamp 1644511149
transform 1 0 4140 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_39
timestamp 1644511149
transform 1 0 4692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_51
timestamp 1644511149
transform 1 0 5796 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_63
timestamp 1644511149
transform 1 0 6900 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_75
timestamp 1644511149
transform 1 0 8004 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_13
timestamp 1644511149
transform 1 0 2300 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_22
timestamp 1644511149
transform 1 0 3128 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_43
timestamp 1644511149
transform 1 0 5060 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_50
timestamp 1644511149
transform 1 0 5704 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_99
timestamp 1644511149
transform 1 0 10212 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_14
timestamp 1644511149
transform 1 0 2392 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_22
timestamp 1644511149
transform 1 0 3128 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_33
timestamp 1644511149
transform 1 0 4140 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_45
timestamp 1644511149
transform 1 0 5244 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_57
timestamp 1644511149
transform 1 0 6348 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_69
timestamp 1644511149
transform 1 0 7452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_81
timestamp 1644511149
transform 1 0 8556 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_93
timestamp 1644511149
transform 1 0 9660 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_99
timestamp 1644511149
transform 1 0 10212 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_7
timestamp 1644511149
transform 1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_25
timestamp 1644511149
transform 1 0 3404 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1644511149
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1644511149
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_99
timestamp 1644511149
transform 1 0 10212 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_16
timestamp 1644511149
transform 1 0 2576 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_24
timestamp 1644511149
transform 1 0 3312 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_34
timestamp 1644511149
transform 1 0 4232 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_42
timestamp 1644511149
transform 1 0 4968 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_54
timestamp 1644511149
transform 1 0 6072 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_66
timestamp 1644511149
transform 1 0 7176 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_78
timestamp 1644511149
transform 1 0 8280 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_91
timestamp 1644511149
transform 1 0 9476 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_99
timestamp 1644511149
transform 1 0 10212 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_7
timestamp 1644511149
transform 1 0 1748 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_23
timestamp 1644511149
transform 1 0 3220 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_31
timestamp 1644511149
transform 1 0 3956 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_42
timestamp 1644511149
transform 1 0 4968 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_54
timestamp 1644511149
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_99
timestamp 1644511149
transform 1 0 10212 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_7
timestamp 1644511149
transform 1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_16
timestamp 1644511149
transform 1 0 2576 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_52
timestamp 1644511149
transform 1 0 5888 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_64
timestamp 1644511149
transform 1 0 6992 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_76
timestamp 1644511149
transform 1 0 8096 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_93
timestamp 1644511149
transform 1 0 9660 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_99
timestamp 1644511149
transform 1 0 10212 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_7
timestamp 1644511149
transform 1 0 1748 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_18
timestamp 1644511149
transform 1 0 2760 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_30
timestamp 1644511149
transform 1 0 3864 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_42
timestamp 1644511149
transform 1 0 4968 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_54
timestamp 1644511149
transform 1 0 6072 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_101
timestamp 1644511149
transform 1 0 10396 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_13
timestamp 1644511149
transform 1 0 2300 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1644511149
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_33
timestamp 1644511149
transform 1 0 4140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_45
timestamp 1644511149
transform 1 0 5244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_57
timestamp 1644511149
transform 1 0 6348 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_69
timestamp 1644511149
transform 1 0 7452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_81
timestamp 1644511149
transform 1 0 8556 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_93
timestamp 1644511149
transform 1 0 9660 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_99
timestamp 1644511149
transform 1 0 10212 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_10
timestamp 1644511149
transform 1 0 2024 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_18
timestamp 1644511149
transform 1 0 2760 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_24
timestamp 1644511149
transform 1 0 3312 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_32
timestamp 1644511149
transform 1 0 4048 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_44
timestamp 1644511149
transform 1 0 5152 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_99
timestamp 1644511149
transform 1 0 10212 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_14
timestamp 1644511149
transform 1 0 2392 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_23
timestamp 1644511149
transform 1 0 3220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_33
timestamp 1644511149
transform 1 0 4140 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_41
timestamp 1644511149
transform 1 0 4876 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_47
timestamp 1644511149
transform 1 0 5428 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_59
timestamp 1644511149
transform 1 0 6532 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_67
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_72
timestamp 1644511149
transform 1 0 7728 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_99
timestamp 1644511149
transform 1 0 10212 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_8
timestamp 1644511149
transform 1 0 1840 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_22
timestamp 1644511149
transform 1 0 3128 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_30
timestamp 1644511149
transform 1 0 3864 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_42
timestamp 1644511149
transform 1 0 4968 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_54
timestamp 1644511149
transform 1 0 6072 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1644511149
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1644511149
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_93
timestamp 1644511149
transform 1 0 9660 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_99
timestamp 1644511149
transform 1 0 10212 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_7
timestamp 1644511149
transform 1 0 1748 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_13
timestamp 1644511149
transform 1 0 2300 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_19
timestamp 1644511149
transform 1 0 2852 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1644511149
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_29
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_33
timestamp 1644511149
transform 1 0 4140 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_39
timestamp 1644511149
transform 1 0 4692 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_48
timestamp 1644511149
transform 1 0 5520 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_60
timestamp 1644511149
transform 1 0 6624 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1644511149
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1644511149
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1644511149
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_91
timestamp 1644511149
transform 1 0 9476 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_99
timestamp 1644511149
transform 1 0 10212 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_7
timestamp 1644511149
transform 1 0 1748 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_23
timestamp 1644511149
transform 1 0 3220 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_32
timestamp 1644511149
transform 1 0 4048 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_44
timestamp 1644511149
transform 1 0 5152 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1644511149
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_81
timestamp 1644511149
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_93
timestamp 1644511149
transform 1 0 9660 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_99
timestamp 1644511149
transform 1 0 10212 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_7
timestamp 1644511149
transform 1 0 1748 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1644511149
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1644511149
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_29
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_41
timestamp 1644511149
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_53
timestamp 1644511149
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_65
timestamp 1644511149
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1644511149
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1644511149
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_86_85
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_91
timestamp 1644511149
transform 1 0 9476 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_99
timestamp 1644511149
transform 1 0 10212 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_10
timestamp 1644511149
transform 1 0 2024 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_18
timestamp 1644511149
transform 1 0 2760 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_30
timestamp 1644511149
transform 1 0 3864 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_42
timestamp 1644511149
transform 1 0 4968 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_54
timestamp 1644511149
transform 1 0 6072 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1644511149
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1644511149
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1644511149
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_93
timestamp 1644511149
transform 1 0 9660 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_99
timestamp 1644511149
transform 1 0 10212 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_10
timestamp 1644511149
transform 1 0 2024 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_18
timestamp 1644511149
transform 1 0 2760 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1644511149
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_88_29
timestamp 1644511149
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_41
timestamp 1644511149
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_53
timestamp 1644511149
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_65
timestamp 1644511149
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1644511149
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1644511149
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_85
timestamp 1644511149
transform 1 0 8924 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_93
timestamp 1644511149
transform 1 0 9660 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_99
timestamp 1644511149
transform 1 0 10212 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_10
timestamp 1644511149
transform 1 0 2024 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_14
timestamp 1644511149
transform 1 0 2392 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_20
timestamp 1644511149
transform 1 0 2944 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_29
timestamp 1644511149
transform 1 0 3772 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_41
timestamp 1644511149
transform 1 0 4876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_53
timestamp 1644511149
transform 1 0 5980 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1644511149
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1644511149
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1644511149
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_93
timestamp 1644511149
transform 1 0 9660 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_99
timestamp 1644511149
transform 1 0 10212 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_7
timestamp 1644511149
transform 1 0 1748 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_16
timestamp 1644511149
transform 1 0 2576 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_23
timestamp 1644511149
transform 1 0 3220 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1644511149
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1644511149
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_41
timestamp 1644511149
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_53
timestamp 1644511149
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_65
timestamp 1644511149
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1644511149
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1644511149
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_85
timestamp 1644511149
transform 1 0 8924 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_93
timestamp 1644511149
transform 1 0 9660 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_99
timestamp 1644511149
transform 1 0 10212 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_7
timestamp 1644511149
transform 1 0 1748 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_15
timestamp 1644511149
transform 1 0 2484 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_23
timestamp 1644511149
transform 1 0 3220 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_35
timestamp 1644511149
transform 1 0 4324 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_47
timestamp 1644511149
transform 1 0 5428 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1644511149
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1644511149
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1644511149
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1644511149
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_93
timestamp 1644511149
transform 1 0 9660 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_99
timestamp 1644511149
transform 1 0 10212 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_7
timestamp 1644511149
transform 1 0 1748 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_14
timestamp 1644511149
transform 1 0 2392 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_26
timestamp 1644511149
transform 1 0 3496 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1644511149
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_41
timestamp 1644511149
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_53
timestamp 1644511149
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_65
timestamp 1644511149
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1644511149
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1644511149
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_85
timestamp 1644511149
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_97
timestamp 1644511149
transform 1 0 10028 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_7
timestamp 1644511149
transform 1 0 1748 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_19
timestamp 1644511149
transform 1 0 2852 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_31
timestamp 1644511149
transform 1 0 3956 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_43
timestamp 1644511149
transform 1 0 5060 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1644511149
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1644511149
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1644511149
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_81
timestamp 1644511149
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_93
timestamp 1644511149
transform 1 0 9660 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_99
timestamp 1644511149
transform 1 0 10212 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_7
timestamp 1644511149
transform 1 0 1748 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1644511149
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1644511149
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1644511149
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1644511149
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_53
timestamp 1644511149
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1644511149
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1644511149
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1644511149
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_85
timestamp 1644511149
transform 1 0 8924 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_93
timestamp 1644511149
transform 1 0 9660 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_99
timestamp 1644511149
transform 1 0 10212 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_11
timestamp 1644511149
transform 1 0 2116 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_19
timestamp 1644511149
transform 1 0 2852 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_31
timestamp 1644511149
transform 1 0 3956 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_43
timestamp 1644511149
transform 1 0 5060 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1644511149
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1644511149
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1644511149
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_81
timestamp 1644511149
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_93
timestamp 1644511149
transform 1 0 9660 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_99
timestamp 1644511149
transform 1 0 10212 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_11
timestamp 1644511149
transform 1 0 2116 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_19
timestamp 1644511149
transform 1 0 2852 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1644511149
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1644511149
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1644511149
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1644511149
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1644511149
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1644511149
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1644511149
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_85
timestamp 1644511149
transform 1 0 8924 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_92
timestamp 1644511149
transform 1 0 9568 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_99
timestamp 1644511149
transform 1 0 10212 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_97_7
timestamp 1644511149
transform 1 0 1748 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_13
timestamp 1644511149
transform 1 0 2300 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_19
timestamp 1644511149
transform 1 0 2852 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_28
timestamp 1644511149
transform 1 0 3680 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_37
timestamp 1644511149
transform 1 0 4508 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_49
timestamp 1644511149
transform 1 0 5612 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1644511149
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1644511149
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1644511149
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_81
timestamp 1644511149
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_93
timestamp 1644511149
transform 1 0 9660 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_99
timestamp 1644511149
transform 1 0 10212 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_7
timestamp 1644511149
transform 1 0 1748 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_15
timestamp 1644511149
transform 1 0 2484 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_24
timestamp 1644511149
transform 1 0 3312 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_34
timestamp 1644511149
transform 1 0 4232 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_46
timestamp 1644511149
transform 1 0 5336 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_58
timestamp 1644511149
transform 1 0 6440 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_70
timestamp 1644511149
transform 1 0 7544 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_98_82
timestamp 1644511149
transform 1 0 8648 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_98_85
timestamp 1644511149
transform 1 0 8924 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_93
timestamp 1644511149
transform 1 0 9660 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_99
timestamp 1644511149
transform 1 0 10212 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_7
timestamp 1644511149
transform 1 0 1748 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_15
timestamp 1644511149
transform 1 0 2484 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_23
timestamp 1644511149
transform 1 0 3220 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_30
timestamp 1644511149
transform 1 0 3864 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_42
timestamp 1644511149
transform 1 0 4968 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_54
timestamp 1644511149
transform 1 0 6072 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_57
timestamp 1644511149
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_69
timestamp 1644511149
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_81
timestamp 1644511149
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_93
timestamp 1644511149
transform 1 0 9660 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_99
timestamp 1644511149
transform 1 0 10212 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_11
timestamp 1644511149
transform 1 0 2116 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_18
timestamp 1644511149
transform 1 0 2760 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_26
timestamp 1644511149
transform 1 0 3496 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_29
timestamp 1644511149
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_41
timestamp 1644511149
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_53
timestamp 1644511149
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_65
timestamp 1644511149
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1644511149
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1644511149
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_85
timestamp 1644511149
transform 1 0 8924 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_99
timestamp 1644511149
transform 1 0 10212 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_11
timestamp 1644511149
transform 1 0 2116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_23
timestamp 1644511149
transform 1 0 3220 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_35
timestamp 1644511149
transform 1 0 4324 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_47
timestamp 1644511149
transform 1 0 5428 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1644511149
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1644511149
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1644511149
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_81
timestamp 1644511149
transform 1 0 8556 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_99
timestamp 1644511149
transform 1 0 10212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_7
timestamp 1644511149
transform 1 0 1748 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_15
timestamp 1644511149
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1644511149
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_29
timestamp 1644511149
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_41
timestamp 1644511149
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_53
timestamp 1644511149
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_65
timestamp 1644511149
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1644511149
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1644511149
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_85
timestamp 1644511149
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_97
timestamp 1644511149
transform 1 0 10028 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_103_7
timestamp 1644511149
transform 1 0 1748 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_103_20
timestamp 1644511149
transform 1 0 2944 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_28
timestamp 1644511149
transform 1 0 3680 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_40
timestamp 1644511149
transform 1 0 4784 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_52
timestamp 1644511149
transform 1 0 5888 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_57
timestamp 1644511149
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_69
timestamp 1644511149
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_81
timestamp 1644511149
transform 1 0 8556 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_103_99
timestamp 1644511149
transform 1 0 10212 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_6
timestamp 1644511149
transform 1 0 1656 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_104_18
timestamp 1644511149
transform 1 0 2760 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_104_26
timestamp 1644511149
transform 1 0 3496 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_104_33
timestamp 1644511149
transform 1 0 4140 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_45
timestamp 1644511149
transform 1 0 5244 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_57
timestamp 1644511149
transform 1 0 6348 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_69
timestamp 1644511149
transform 1 0 7452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_104_81
timestamp 1644511149
transform 1 0 8556 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_104_85
timestamp 1644511149
transform 1 0 8924 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_104_93
timestamp 1644511149
transform 1 0 9660 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_104_99
timestamp 1644511149
transform 1 0 10212 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_19
timestamp 1644511149
transform 1 0 2852 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_31
timestamp 1644511149
transform 1 0 3956 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_43
timestamp 1644511149
transform 1 0 5060 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1644511149
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_57
timestamp 1644511149
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_69
timestamp 1644511149
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_81
timestamp 1644511149
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_105_93
timestamp 1644511149
transform 1 0 9660 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_99
timestamp 1644511149
transform 1 0 10212 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_106_3
timestamp 1644511149
transform 1 0 1380 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_13
timestamp 1644511149
transform 1 0 2300 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_106_19
timestamp 1644511149
transform 1 0 2852 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1644511149
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1644511149
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1644511149
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_53
timestamp 1644511149
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_65
timestamp 1644511149
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1644511149
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1644511149
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_85
timestamp 1644511149
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_97
timestamp 1644511149
transform 1 0 10028 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_107_7
timestamp 1644511149
transform 1 0 1748 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_15
timestamp 1644511149
transform 1 0 2484 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_23
timestamp 1644511149
transform 1 0 3220 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_35
timestamp 1644511149
transform 1 0 4324 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_47
timestamp 1644511149
transform 1 0 5428 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1644511149
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_57
timestamp 1644511149
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_69
timestamp 1644511149
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_81
timestamp 1644511149
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_107_93
timestamp 1644511149
transform 1 0 9660 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_99
timestamp 1644511149
transform 1 0 10212 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_11
timestamp 1644511149
transform 1 0 2116 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_19
timestamp 1644511149
transform 1 0 2852 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1644511149
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_29
timestamp 1644511149
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_41
timestamp 1644511149
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_53
timestamp 1644511149
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_65
timestamp 1644511149
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1644511149
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1644511149
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_85
timestamp 1644511149
transform 1 0 8924 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_108_93
timestamp 1644511149
transform 1 0 9660 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_99
timestamp 1644511149
transform 1 0 10212 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_11
timestamp 1644511149
transform 1 0 2116 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_15
timestamp 1644511149
transform 1 0 2484 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_109_22
timestamp 1644511149
transform 1 0 3128 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_109_30
timestamp 1644511149
transform 1 0 3864 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_42
timestamp 1644511149
transform 1 0 4968 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_54
timestamp 1644511149
transform 1 0 6072 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_57
timestamp 1644511149
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_69
timestamp 1644511149
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_81
timestamp 1644511149
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_93
timestamp 1644511149
transform 1 0 9660 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_101
timestamp 1644511149
transform 1 0 10396 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_110_3
timestamp 1644511149
transform 1 0 1380 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_110_17
timestamp 1644511149
transform 1 0 2668 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_110_25
timestamp 1644511149
transform 1 0 3404 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_29
timestamp 1644511149
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_41
timestamp 1644511149
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_53
timestamp 1644511149
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_65
timestamp 1644511149
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1644511149
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1644511149
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_85
timestamp 1644511149
transform 1 0 8924 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_110_93
timestamp 1644511149
transform 1 0 9660 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_110_99
timestamp 1644511149
transform 1 0 10212 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_111_7
timestamp 1644511149
transform 1 0 1748 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_15
timestamp 1644511149
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_27
timestamp 1644511149
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_39
timestamp 1644511149
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_51
timestamp 1644511149
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1644511149
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_57
timestamp 1644511149
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_69
timestamp 1644511149
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_81
timestamp 1644511149
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_93
timestamp 1644511149
transform 1 0 9660 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_111_99
timestamp 1644511149
transform 1 0 10212 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_7
timestamp 1644511149
transform 1 0 1748 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_15
timestamp 1644511149
transform 1 0 2484 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_23
timestamp 1644511149
transform 1 0 3220 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1644511149
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_29
timestamp 1644511149
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_41
timestamp 1644511149
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_53
timestamp 1644511149
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_65
timestamp 1644511149
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_77
timestamp 1644511149
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1644511149
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_85
timestamp 1644511149
transform 1 0 8924 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_112_93
timestamp 1644511149
transform 1 0 9660 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_112_99
timestamp 1644511149
transform 1 0 10212 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_113_7
timestamp 1644511149
transform 1 0 1748 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_113_15
timestamp 1644511149
transform 1 0 2484 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_113_22
timestamp 1644511149
transform 1 0 3128 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_113_32
timestamp 1644511149
transform 1 0 4048 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_44
timestamp 1644511149
transform 1 0 5152 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_57
timestamp 1644511149
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_69
timestamp 1644511149
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_81
timestamp 1644511149
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_93
timestamp 1644511149
transform 1 0 9660 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_113_101
timestamp 1644511149
transform 1 0 10396 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_114_3
timestamp 1644511149
transform 1 0 1380 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_114_17
timestamp 1644511149
transform 1 0 2668 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_114_25
timestamp 1644511149
transform 1 0 3404 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_114_33
timestamp 1644511149
transform 1 0 4140 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_45
timestamp 1644511149
transform 1 0 5244 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_57
timestamp 1644511149
transform 1 0 6348 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_69
timestamp 1644511149
transform 1 0 7452 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_114_81
timestamp 1644511149
transform 1 0 8556 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_114_85
timestamp 1644511149
transform 1 0 8924 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_114_93
timestamp 1644511149
transform 1 0 9660 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_114_99
timestamp 1644511149
transform 1 0 10212 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_11
timestamp 1644511149
transform 1 0 2116 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_22
timestamp 1644511149
transform 1 0 3128 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_115_32
timestamp 1644511149
transform 1 0 4048 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_44
timestamp 1644511149
transform 1 0 5152 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_57
timestamp 1644511149
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_69
timestamp 1644511149
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_81
timestamp 1644511149
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_115_93
timestamp 1644511149
transform 1 0 9660 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_115_99
timestamp 1644511149
transform 1 0 10212 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_6
timestamp 1644511149
transform 1 0 1656 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_116_18
timestamp 1644511149
transform 1 0 2760 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_116_26
timestamp 1644511149
transform 1 0 3496 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_116_33
timestamp 1644511149
transform 1 0 4140 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_45
timestamp 1644511149
transform 1 0 5244 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_57
timestamp 1644511149
transform 1 0 6348 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_69
timestamp 1644511149
transform 1 0 7452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_116_81
timestamp 1644511149
transform 1 0 8556 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_85
timestamp 1644511149
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_97
timestamp 1644511149
transform 1 0 10028 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_3
timestamp 1644511149
transform 1 0 1380 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_12
timestamp 1644511149
transform 1 0 2208 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_117_20
timestamp 1644511149
transform 1 0 2944 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_32
timestamp 1644511149
transform 1 0 4048 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_44
timestamp 1644511149
transform 1 0 5152 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_57
timestamp 1644511149
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_69
timestamp 1644511149
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_81
timestamp 1644511149
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_93
timestamp 1644511149
transform 1 0 9660 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_117_99
timestamp 1644511149
transform 1 0 10212 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_11
timestamp 1644511149
transform 1 0 2116 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_118_19
timestamp 1644511149
transform 1 0 2852 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1644511149
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_29
timestamp 1644511149
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_41
timestamp 1644511149
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_53
timestamp 1644511149
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_65
timestamp 1644511149
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1644511149
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1644511149
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_85
timestamp 1644511149
transform 1 0 8924 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_93
timestamp 1644511149
transform 1 0 9660 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_118_99
timestamp 1644511149
transform 1 0 10212 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_13
timestamp 1644511149
transform 1 0 2300 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_119_20
timestamp 1644511149
transform 1 0 2944 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_32
timestamp 1644511149
transform 1 0 4048 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_44
timestamp 1644511149
transform 1 0 5152 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_57
timestamp 1644511149
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_69
timestamp 1644511149
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_81
timestamp 1644511149
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_93
timestamp 1644511149
transform 1 0 9660 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_99
timestamp 1644511149
transform 1 0 10212 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_120_13
timestamp 1644511149
transform 1 0 2300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_25
timestamp 1644511149
transform 1 0 3404 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_120_29
timestamp 1644511149
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_41
timestamp 1644511149
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_53
timestamp 1644511149
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_65
timestamp 1644511149
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1644511149
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1644511149
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_85
timestamp 1644511149
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_97
timestamp 1644511149
transform 1 0 10028 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_121_13
timestamp 1644511149
transform 1 0 2300 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_25
timestamp 1644511149
transform 1 0 3404 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_37
timestamp 1644511149
transform 1 0 4508 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_49
timestamp 1644511149
transform 1 0 5612 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1644511149
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_57
timestamp 1644511149
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_69
timestamp 1644511149
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_81
timestamp 1644511149
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_121_93
timestamp 1644511149
transform 1 0 9660 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_121_99
timestamp 1644511149
transform 1 0 10212 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_122_6
timestamp 1644511149
transform 1 0 1656 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_12
timestamp 1644511149
transform 1 0 2208 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_122_21
timestamp 1644511149
transform 1 0 3036 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1644511149
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_29
timestamp 1644511149
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_41
timestamp 1644511149
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_53
timestamp 1644511149
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_65
timestamp 1644511149
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1644511149
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1644511149
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_85
timestamp 1644511149
transform 1 0 8924 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_93
timestamp 1644511149
transform 1 0 9660 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_99
timestamp 1644511149
transform 1 0 10212 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_11
timestamp 1644511149
transform 1 0 2116 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_123_18
timestamp 1644511149
transform 1 0 2760 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_30
timestamp 1644511149
transform 1 0 3864 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_42
timestamp 1644511149
transform 1 0 4968 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_54
timestamp 1644511149
transform 1 0 6072 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_57
timestamp 1644511149
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_69
timestamp 1644511149
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_81
timestamp 1644511149
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_93
timestamp 1644511149
transform 1 0 9660 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_123_101
timestamp 1644511149
transform 1 0 10396 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_124_6
timestamp 1644511149
transform 1 0 1656 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_124_13
timestamp 1644511149
transform 1 0 2300 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_124_20
timestamp 1644511149
transform 1 0 2944 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_124_29
timestamp 1644511149
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_41
timestamp 1644511149
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_53
timestamp 1644511149
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_65
timestamp 1644511149
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1644511149
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1644511149
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_85
timestamp 1644511149
transform 1 0 8924 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_124_93
timestamp 1644511149
transform 1 0 9660 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_124_99
timestamp 1644511149
transform 1 0 10212 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_125_11
timestamp 1644511149
transform 1 0 2116 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_125_18
timestamp 1644511149
transform 1 0 2760 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_30
timestamp 1644511149
transform 1 0 3864 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_42
timestamp 1644511149
transform 1 0 4968 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_125_54
timestamp 1644511149
transform 1 0 6072 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_125_57
timestamp 1644511149
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_69
timestamp 1644511149
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_81
timestamp 1644511149
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_125_93
timestamp 1644511149
transform 1 0 9660 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_125_99
timestamp 1644511149
transform 1 0 10212 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_126_6
timestamp 1644511149
transform 1 0 1656 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_18
timestamp 1644511149
transform 1 0 2760 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_126_26
timestamp 1644511149
transform 1 0 3496 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_126_29
timestamp 1644511149
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_41
timestamp 1644511149
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_53
timestamp 1644511149
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_65
timestamp 1644511149
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1644511149
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1644511149
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_85
timestamp 1644511149
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_97
timestamp 1644511149
transform 1 0 10028 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_127_11
timestamp 1644511149
transform 1 0 2116 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_127_23
timestamp 1644511149
transform 1 0 3220 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_35
timestamp 1644511149
transform 1 0 4324 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_47
timestamp 1644511149
transform 1 0 5428 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1644511149
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_57
timestamp 1644511149
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_69
timestamp 1644511149
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_81
timestamp 1644511149
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_93
timestamp 1644511149
transform 1 0 9660 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_127_99
timestamp 1644511149
transform 1 0 10212 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_128_6
timestamp 1644511149
transform 1 0 1656 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_128_13
timestamp 1644511149
transform 1 0 2300 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_128_20
timestamp 1644511149
transform 1 0 2944 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_128_29
timestamp 1644511149
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_41
timestamp 1644511149
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_53
timestamp 1644511149
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_65
timestamp 1644511149
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1644511149
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1644511149
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_85
timestamp 1644511149
transform 1 0 8924 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_128_93
timestamp 1644511149
transform 1 0 9660 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_128_99
timestamp 1644511149
transform 1 0 10212 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_129_11
timestamp 1644511149
transform 1 0 2116 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_129_23
timestamp 1644511149
transform 1 0 3220 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_35
timestamp 1644511149
transform 1 0 4324 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_47
timestamp 1644511149
transform 1 0 5428 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_129_55
timestamp 1644511149
transform 1 0 6164 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_57
timestamp 1644511149
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_69
timestamp 1644511149
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_81
timestamp 1644511149
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_129_93
timestamp 1644511149
transform 1 0 9660 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_129_99
timestamp 1644511149
transform 1 0 10212 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_130_6
timestamp 1644511149
transform 1 0 1656 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_18
timestamp 1644511149
transform 1 0 2760 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_130_26
timestamp 1644511149
transform 1 0 3496 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_130_29
timestamp 1644511149
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_41
timestamp 1644511149
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_53
timestamp 1644511149
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_65
timestamp 1644511149
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1644511149
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1644511149
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_85
timestamp 1644511149
transform 1 0 8924 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_97
timestamp 1644511149
transform 1 0 10028 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_131_6
timestamp 1644511149
transform 1 0 1656 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_131_13
timestamp 1644511149
transform 1 0 2300 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_131_20
timestamp 1644511149
transform 1 0 2944 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_32
timestamp 1644511149
transform 1 0 4048 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_44
timestamp 1644511149
transform 1 0 5152 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_57
timestamp 1644511149
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_69
timestamp 1644511149
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_81
timestamp 1644511149
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_131_93
timestamp 1644511149
transform 1 0 9660 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_131_99
timestamp 1644511149
transform 1 0 10212 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_132_3
timestamp 1644511149
transform 1 0 1380 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_132_17
timestamp 1644511149
transform 1 0 2668 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_132_25
timestamp 1644511149
transform 1 0 3404 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_132_29
timestamp 1644511149
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_41
timestamp 1644511149
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_53
timestamp 1644511149
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_65
timestamp 1644511149
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1644511149
transform 1 0 8188 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1644511149
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_85
timestamp 1644511149
transform 1 0 8924 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_132_93
timestamp 1644511149
transform 1 0 9660 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_132_99
timestamp 1644511149
transform 1 0 10212 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_133_11
timestamp 1644511149
transform 1 0 2116 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_133_18
timestamp 1644511149
transform 1 0 2760 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_30
timestamp 1644511149
transform 1 0 3864 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_42
timestamp 1644511149
transform 1 0 4968 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_133_54
timestamp 1644511149
transform 1 0 6072 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_133_57
timestamp 1644511149
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_69
timestamp 1644511149
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_81
timestamp 1644511149
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_93
timestamp 1644511149
transform 1 0 9660 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_133_101
timestamp 1644511149
transform 1 0 10396 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_134_3
timestamp 1644511149
transform 1 0 1380 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_134_17
timestamp 1644511149
transform 1 0 2668 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_134_25
timestamp 1644511149
transform 1 0 3404 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_134_29
timestamp 1644511149
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_41
timestamp 1644511149
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_53
timestamp 1644511149
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_65
timestamp 1644511149
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1644511149
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1644511149
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_85
timestamp 1644511149
transform 1 0 8924 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_134_93
timestamp 1644511149
transform 1 0 9660 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_134_99
timestamp 1644511149
transform 1 0 10212 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_135_6
timestamp 1644511149
transform 1 0 1656 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_135_22
timestamp 1644511149
transform 1 0 3128 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_29
timestamp 1644511149
transform 1 0 3772 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_41
timestamp 1644511149
transform 1 0 4876 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_135_53
timestamp 1644511149
transform 1 0 5980 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_57
timestamp 1644511149
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_69
timestamp 1644511149
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_81
timestamp 1644511149
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_135_93
timestamp 1644511149
transform 1 0 9660 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_135_99
timestamp 1644511149
transform 1 0 10212 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_136_6
timestamp 1644511149
transform 1 0 1656 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_136_20
timestamp 1644511149
transform 1 0 2944 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_136_32
timestamp 1644511149
transform 1 0 4048 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_44
timestamp 1644511149
transform 1 0 5152 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_56
timestamp 1644511149
transform 1 0 6256 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_68
timestamp 1644511149
transform 1 0 7360 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_80
timestamp 1644511149
transform 1 0 8464 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_136_85
timestamp 1644511149
transform 1 0 8924 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_136_93
timestamp 1644511149
transform 1 0 9660 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_136_99
timestamp 1644511149
transform 1 0 10212 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_11
timestamp 1644511149
transform 1 0 2116 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_18
timestamp 1644511149
transform 1 0 2760 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_25
timestamp 1644511149
transform 1 0 3404 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_32
timestamp 1644511149
transform 1 0 4048 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_137_39
timestamp 1644511149
transform 1 0 4692 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_51
timestamp 1644511149
transform 1 0 5796 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1644511149
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_57
timestamp 1644511149
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_69
timestamp 1644511149
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_81
timestamp 1644511149
transform 1 0 8556 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_87
timestamp 1644511149
transform 1 0 9108 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_137_91
timestamp 1644511149
transform 1 0 9476 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_99
timestamp 1644511149
transform 1 0 10212 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_7
timestamp 1644511149
transform 1 0 1748 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_14
timestamp 1644511149
transform 1 0 2392 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_138_21
timestamp 1644511149
transform 1 0 3036 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 1644511149
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_138_32
timestamp 1644511149
transform 1 0 4048 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_138_39
timestamp 1644511149
transform 1 0 4692 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_138_51
timestamp 1644511149
transform 1 0 5796 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_55
timestamp 1644511149
transform 1 0 6164 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_57
timestamp 1644511149
transform 1 0 6348 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_69
timestamp 1644511149
transform 1 0 7452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1644511149
transform 1 0 8556 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_138_85
timestamp 1644511149
transform 1 0 8924 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_91
timestamp 1644511149
transform 1 0 9476 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_99
timestamp 1644511149
transform 1 0 10212 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 10856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 10856 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 10856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 10856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 10856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 10856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 10856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 10856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 10856 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 10856 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 10856 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 10856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 10856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 10856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 10856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 10856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 10856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 10856 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 10856 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 10856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 10856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 10856 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 10856 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 10856 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 10856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 10856 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 10856 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 10856 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 10856 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 10856 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 10856 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 10856 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 10856 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 10856 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 10856 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 10856 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 10856 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 10856 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 10856 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 10856 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 10856 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 10856 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 10856 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 10856 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 10856 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 10856 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 10856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 10856 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 10856 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 10856 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 10856 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 10856 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1644511149
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1644511149
transform -1 0 10856 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1644511149
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1644511149
transform -1 0 10856 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1644511149
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1644511149
transform -1 0 10856 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1644511149
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1644511149
transform -1 0 10856 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1644511149
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1644511149
transform -1 0 10856 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1644511149
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1644511149
transform -1 0 10856 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1644511149
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1644511149
transform -1 0 10856 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1644511149
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1644511149
transform -1 0 10856 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1644511149
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1644511149
transform -1 0 10856 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1644511149
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1644511149
transform -1 0 10856 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1644511149
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1644511149
transform -1 0 10856 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1644511149
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1644511149
transform -1 0 10856 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1644511149
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1644511149
transform -1 0 10856 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1644511149
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1644511149
transform -1 0 10856 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1644511149
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1644511149
transform -1 0 10856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1644511149
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1644511149
transform -1 0 10856 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1644511149
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1644511149
transform -1 0 10856 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1644511149
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1644511149
transform -1 0 10856 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1644511149
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1644511149
transform -1 0 10856 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1644511149
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1644511149
transform -1 0 10856 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1644511149
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1644511149
transform -1 0 10856 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1644511149
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1644511149
transform -1 0 10856 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1644511149
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1644511149
transform -1 0 10856 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1644511149
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1644511149
transform -1 0 10856 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1644511149
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1644511149
transform -1 0 10856 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1644511149
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1644511149
transform -1 0 10856 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1644511149
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1644511149
transform -1 0 10856 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1644511149
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1644511149
transform -1 0 10856 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1644511149
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1644511149
transform -1 0 10856 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1644511149
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1644511149
transform -1 0 10856 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1644511149
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1644511149
transform -1 0 10856 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1644511149
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1644511149
transform -1 0 10856 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1644511149
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1644511149
transform -1 0 10856 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1644511149
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1644511149
transform -1 0 10856 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1644511149
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1644511149
transform -1 0 10856 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1644511149
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1644511149
transform -1 0 10856 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1644511149
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1644511149
transform -1 0 10856 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1644511149
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1644511149
transform -1 0 10856 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1644511149
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1644511149
transform -1 0 10856 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1644511149
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1644511149
transform -1 0 10856 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1644511149
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1644511149
transform -1 0 10856 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1644511149
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1644511149
transform -1 0 10856 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1644511149
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1644511149
transform -1 0 10856 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1644511149
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1644511149
transform -1 0 10856 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1644511149
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1644511149
transform -1 0 10856 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1644511149
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1644511149
transform -1 0 10856 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1644511149
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1644511149
transform -1 0 10856 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1644511149
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1644511149
transform -1 0 10856 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1644511149
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1644511149
transform -1 0 10856 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1644511149
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1644511149
transform -1 0 10856 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1644511149
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1644511149
transform -1 0 10856 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1644511149
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1644511149
transform -1 0 10856 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__or4bb_1  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _096_
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2392 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _100_
timestamp 1644511149
transform 1 0 2576 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_8  _102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4140 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _106_
timestamp 1644511149
transform 1 0 2668 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1644511149
transform 1 0 2668 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _108_
timestamp 1644511149
transform 1 0 2668 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1644511149
transform 1 0 3496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _110_
timestamp 1644511149
transform 1 0 2668 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1644511149
transform 1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _112_
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1644511149
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _114_
timestamp 1644511149
transform 1 0 1840 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _116_
timestamp 1644511149
transform 1 0 1564 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1644511149
transform 1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _118_
timestamp 1644511149
transform 1 0 2668 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1644511149
transform 1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _120_
timestamp 1644511149
transform 1 0 2668 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1644511149
transform 1 0 1932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _122_
timestamp 1644511149
transform 1 0 2668 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _124_
timestamp 1644511149
transform 1 0 2024 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1644511149
transform 1 0 2668 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _126_
timestamp 1644511149
transform 1 0 1564 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1472 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _128_
timestamp 1644511149
transform 1 0 1840 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1644511149
transform 1 0 1748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _130_
timestamp 1644511149
transform 1 0 1564 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1644511149
transform 1 0 1472 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _132_
timestamp 1644511149
transform 1 0 2392 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _133_
timestamp 1644511149
transform 1 0 1472 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _134_
timestamp 1644511149
transform 1 0 2576 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _135_
timestamp 1644511149
transform 1 0 2208 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1644511149
transform 1 0 2760 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _137_
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _138_
timestamp 1644511149
transform 1 0 2760 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _139_
timestamp 1644511149
transform 1 0 1564 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _140_
timestamp 1644511149
transform 1 0 2392 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _141_
timestamp 1644511149
transform 1 0 2760 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _142_
timestamp 1644511149
transform 1 0 2024 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _143_
timestamp 1644511149
transform 1 0 1564 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _144_
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _145_
timestamp 1644511149
transform 1 0 2392 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _146_
timestamp 1644511149
transform 1 0 1748 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _147_
timestamp 1644511149
transform 1 0 2116 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _148_
timestamp 1644511149
transform 1 0 1840 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _149_
timestamp 1644511149
transform 1 0 2760 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _150_
timestamp 1644511149
transform 1 0 2208 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _151_
timestamp 1644511149
transform 1 0 2392 0 1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _152_
timestamp 1644511149
transform 1 0 2300 0 -1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _153_
timestamp 1644511149
transform 1 0 2484 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2944 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _155_
timestamp 1644511149
transform 1 0 2668 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _156_
timestamp 1644511149
transform 1 0 1472 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _157_
timestamp 1644511149
transform 1 0 1564 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _158_
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _159_
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _160_
timestamp 1644511149
transform 1 0 1472 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _161_
timestamp 1644511149
transform 1 0 2116 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1644511149
transform 1 0 2116 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _163_
timestamp 1644511149
transform 1 0 2392 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1644511149
transform 1 0 2484 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _165_
timestamp 1644511149
transform 1 0 3220 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1644511149
transform 1 0 3588 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _167_
timestamp 1644511149
transform 1 0 2484 0 -1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1644511149
transform 1 0 1380 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2576 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2116 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_4  _171_
timestamp 1644511149
transform 1 0 2576 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 -1 65280
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _174_
timestamp 1644511149
transform 1 0 1380 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _175_
timestamp 1644511149
transform 1 0 1380 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _176_
timestamp 1644511149
transform 1 0 1380 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _177_
timestamp 1644511149
transform 1 0 1380 0 -1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _178_
timestamp 1644511149
transform 1 0 1380 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _179_
timestamp 1644511149
transform 1 0 1380 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _180_
timestamp 1644511149
transform 1 0 1380 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _181_
timestamp 1644511149
transform 1 0 1380 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _182_
timestamp 1644511149
transform 1 0 1380 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _183_
timestamp 1644511149
transform 1 0 2116 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _184_
timestamp 1644511149
transform 1 0 2024 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _185_
timestamp 1644511149
transform 1 0 1932 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _186_
timestamp 1644511149
transform 1 0 1932 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _187_
timestamp 1644511149
transform 1 0 2024 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _188_
timestamp 1644511149
transform 1 0 3496 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _189_
timestamp 1644511149
transform 1 0 3496 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _190_
timestamp 1644511149
transform 1 0 1380 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _191_
timestamp 1644511149
transform 1 0 1472 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _192_
timestamp 1644511149
transform 1 0 1380 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _193_
timestamp 1644511149
transform 1 0 2300 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _194_
timestamp 1644511149
transform 1 0 1380 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _195_
timestamp 1644511149
transform 1 0 1380 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _196_
timestamp 1644511149
transform 1 0 1380 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _197_
timestamp 1644511149
transform 1 0 1380 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _198_
timestamp 1644511149
transform 1 0 2484 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _199_
timestamp 1644511149
transform 1 0 2484 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _200_
timestamp 1644511149
transform 1 0 1932 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _201_
timestamp 1644511149
transform 1 0 1932 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _202_
timestamp 1644511149
transform 1 0 2392 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _203_
timestamp 1644511149
transform 1 0 2208 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _204_
timestamp 1644511149
transform 1 0 1380 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _205_
timestamp 1644511149
transform 1 0 1380 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _206_
timestamp 1644511149
transform 1 0 2852 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _207_
timestamp 1644511149
transform 1 0 1932 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _208_
timestamp 1644511149
transform 1 0 2760 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1644511149
transform 1 0 4324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _210_
timestamp 1644511149
transform 1 0 2668 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 1644511149
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _212_
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _214_
timestamp 1644511149
transform 1 0 3496 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1644511149
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _216_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1644511149
transform 1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _218_
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1644511149
transform 1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _220_
timestamp 1644511149
transform 1 0 2668 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1644511149
transform 1 0 7636 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _222_
timestamp 1644511149
transform 1 0 2760 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1644511149
transform 1 0 3864 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _224_
timestamp 1644511149
transform 1 0 2668 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1644511149
transform 1 0 4508 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _226_
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _228_
timestamp 1644511149
transform 1 0 2668 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1644511149
transform 1 0 4232 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _230_
timestamp 1644511149
transform 1 0 2300 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _232_
timestamp 1644511149
transform 1 0 2668 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _233_
timestamp 1644511149
transform 1 0 4232 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _234_
timestamp 1644511149
transform 1 0 3496 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _235_
timestamp 1644511149
transform 1 0 4508 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _236_
timestamp 1644511149
transform 1 0 2668 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _238_
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _239_
timestamp 1644511149
transform 1 0 4140 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1644511149
transform 1 0 9936 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _241_
timestamp 1644511149
transform 1 0 4508 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1644511149
transform 1 0 9936 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _243_
timestamp 1644511149
transform 1 0 4600 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1644511149
transform 1 0 9200 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _245_
timestamp 1644511149
transform 1 0 3956 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1644511149
transform 1 0 9936 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _247_
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _249_
timestamp 1644511149
transform 1 0 4232 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1644511149
transform 1 0 5336 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _251_
timestamp 1644511149
transform 1 0 4232 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1644511149
transform 1 0 9200 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _253_
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1644511149
transform 1 0 9936 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _255_
timestamp 1644511149
transform 1 0 3864 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1644511149
transform 1 0 9936 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _257_
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _258_
timestamp 1644511149
transform 1 0 9200 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _259_
timestamp 1644511149
transform 1 0 4232 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _261_
timestamp 1644511149
transform 1 0 4324 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1644511149
transform 1 0 5520 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _263_
timestamp 1644511149
transform 1 0 4508 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1644511149
transform 1 0 5612 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _265_
timestamp 1644511149
transform 1 0 4968 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _266_
timestamp 1644511149
transform 1 0 7452 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _267_
timestamp 1644511149
transform 1 0 5060 0 1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp 1644511149
transform 1 0 6808 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _269_
timestamp 1644511149
transform 1 0 4232 0 1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _270_
timestamp 1644511149
transform 1 0 9200 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _271_
timestamp 1644511149
transform 1 0 2760 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 1644511149
transform 1 0 9936 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _273_
timestamp 1644511149
transform 1 0 2852 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1644511149
transform 1 0 9936 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _275_
timestamp 1644511149
transform 1 0 3588 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1644511149
transform 1 0 9200 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _277_
timestamp 1644511149
transform 1 0 3312 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _278_
timestamp 1644511149
transform 1 0 9936 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _279_
timestamp 1644511149
transform 1 0 4048 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp 1644511149
transform 1 0 9936 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _281_
timestamp 1644511149
transform 1 0 3772 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1644511149
transform 1 0 9292 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _283_
timestamp 1644511149
transform 1 0 2852 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 1644511149
transform 1 0 9936 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _285_
timestamp 1644511149
transform 1 0 2024 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _286_
timestamp 1644511149
transform 1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _287_
timestamp 1644511149
transform 1 0 2668 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _289_
timestamp 1644511149
transform 1 0 1656 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _290_
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _291_
timestamp 1644511149
transform 1 0 1840 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _292_
timestamp 1644511149
transform 1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _293_
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _294_
timestamp 1644511149
transform 1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _295_
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _296_
timestamp 1644511149
transform 1 0 2668 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _297__290 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9936 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _298__291
timestamp 1644511149
transform 1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _299__280
timestamp 1644511149
transform 1 0 9936 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _300__281
timestamp 1644511149
transform 1 0 9936 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _301__282
timestamp 1644511149
transform 1 0 9936 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _302__283
timestamp 1644511149
transform 1 0 9936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _303__284
timestamp 1644511149
transform 1 0 9936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _304__285
timestamp 1644511149
transform 1 0 9936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _305__286
timestamp 1644511149
transform 1 0 9936 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _306__287
timestamp 1644511149
transform 1 0 9936 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _307__288
timestamp 1644511149
transform 1 0 9936 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _308__289
timestamp 1644511149
transform 1 0 9936 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1644511149
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1644511149
transform 1 0 2668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1644511149
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp 1644511149
transform 1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 1644511149
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1644511149
transform 1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp 1644511149
transform 1 0 3404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1644511149
transform 1 0 2392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp 1644511149
transform 1 0 3036 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1644511149
transform 1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _321_
timestamp 1644511149
transform 1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1644511149
transform 1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1644511149
transform 1 0 9936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1644511149
transform 1 0 9200 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp 1644511149
transform 1 0 9936 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1644511149
transform 1 0 9200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1644511149
transform 1 0 9844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1644511149
transform 1 0 9200 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _330_
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _331_
timestamp 1644511149
transform 1 0 2668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _332_
timestamp 1644511149
transform 1 0 2668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _333_
timestamp 1644511149
transform 1 0 2668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _334_
timestamp 1644511149
transform 1 0 2300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _335_
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _336_
timestamp 1644511149
transform 1 0 2576 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _337_
timestamp 1644511149
transform 1 0 4140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _338_
timestamp 1644511149
transform 1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _339_
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _340_
timestamp 1644511149
transform 1 0 1656 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _341_
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1644511149
transform 1 0 9844 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 9936 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 9936 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 9936 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 9936 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 9936 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 9936 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 9936 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 9936 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 9936 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 9936 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 9936 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 9936 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 9936 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 9936 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 9936 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 9936 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 9936 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 9936 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 9936 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 9936 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 9936 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 9200 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1644511149
transform 1 0 9292 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 9200 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1644511149
transform 1 0 9844 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1644511149
transform 1 0 9292 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1644511149
transform 1 0 9292 0 -1 58752
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 9936 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 9936 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 9936 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 9936 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 9936 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 2116 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 1380 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 1380 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 1380 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 1380 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 2024 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 2668 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 1380 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 1380 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 2024 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 2668 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 2484 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 2668 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 1380 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 1380 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 3496 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 2484 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 3772 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform 1 0 3128 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform 1 0 2760 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform 1 0 3772 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1644511149
transform 1 0 3772 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform 1 0 4416 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1644511149
transform 1 0 1380 0 -1 67456
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1644511149
transform 1 0 4416 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1644511149
transform 1 0 1380 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1644511149
transform 1 0 1380 0 1 67456
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1644511149
transform 1 0 1380 0 -1 68544
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1644511149
transform 1 0 1380 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1644511149
transform 1 0 2484 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1644511149
transform 1 0 2024 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1644511149
transform 1 0 2668 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1644511149
transform 1 0 2484 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input68
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1644511149
transform 1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1644511149
transform 1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1644511149
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1644511149
transform 1 0 3680 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1644511149
transform 1 0 2668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input89
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1644511149
transform 1 0 3128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input94
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input95
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input96
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1644511149
transform 1 0 2116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1644511149
transform 1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input101
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input102
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input103
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input104
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input105
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input106
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input107
timestamp 1644511149
transform 1 0 2668 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1644511149
transform 1 0 3220 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input110
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input112
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input113
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input114
timestamp 1644511149
transform 1 0 4140 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1644511149
transform 1 0 3496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1644511149
transform 1 0 3496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input117
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input118
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1644511149
transform 1 0 2668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1644511149
transform 1 0 1564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input123
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input124
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1644511149
transform 1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1644511149
transform 1 0 2668 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input128
timestamp 1644511149
transform 1 0 2576 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input129
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input130
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input131
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1644511149
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1644511149
transform 1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input136
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input137
timestamp 1644511149
transform 1 0 5060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1644511149
transform 1 0 9844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1644511149
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1644511149
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1644511149
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1644511149
transform 1 0 9844 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1644511149
transform 1 0 9844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1644511149
transform 1 0 9844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1644511149
transform 1 0 9844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1644511149
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1644511149
transform 1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1644511149
transform 1 0 9844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1644511149
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1644511149
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1644511149
transform 1 0 9844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1644511149
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1644511149
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1644511149
transform 1 0 9844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1644511149
transform 1 0 9844 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1644511149
transform 1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1644511149
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1644511149
transform 1 0 9844 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1644511149
transform 1 0 9844 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1644511149
transform 1 0 9844 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1644511149
transform 1 0 9844 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1644511149
transform 1 0 9844 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1644511149
transform 1 0 9844 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1644511149
transform 1 0 9844 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1644511149
transform 1 0 9844 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1644511149
transform 1 0 9844 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1644511149
transform 1 0 9844 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1644511149
transform 1 0 9844 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1644511149
transform 1 0 9844 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1644511149
transform 1 0 9844 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1644511149
transform 1 0 9844 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1644511149
transform 1 0 9844 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1644511149
transform 1 0 9844 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1644511149
transform 1 0 9844 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1644511149
transform 1 0 9844 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1644511149
transform 1 0 9844 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1644511149
transform 1 0 9844 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1644511149
transform 1 0 9844 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1644511149
transform 1 0 9844 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1644511149
transform 1 0 9844 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1644511149
transform 1 0 9844 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1644511149
transform 1 0 9844 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1644511149
transform 1 0 9844 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1644511149
transform 1 0 9844 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1644511149
transform 1 0 9844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1644511149
transform 1 0 9844 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1644511149
transform 1 0 9844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1644511149
transform 1 0 9844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1644511149
transform 1 0 9844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1644511149
transform 1 0 9844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1644511149
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1644511149
transform 1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1644511149
transform 1 0 9844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1644511149
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1644511149
transform 1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1644511149
transform 1 0 1380 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1644511149
transform 1 0 2116 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1644511149
transform 1 0 2392 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1644511149
transform 1 0 2392 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1644511149
transform 1 0 1380 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1644511149
transform 1 0 1380 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1644511149
transform 1 0 2116 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1644511149
transform 1 0 2852 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1644511149
transform 1 0 1380 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1644511149
transform 1 0 1380 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1644511149
transform 1 0 1380 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1644511149
transform 1 0 1380 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1644511149
transform 1 0 2116 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1644511149
transform 1 0 3312 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1644511149
transform 1 0 3772 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1644511149
transform 1 0 1380 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1644511149
transform -1 0 2852 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1644511149
transform 1 0 2116 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1644511149
transform 1 0 2852 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1644511149
transform 1 0 1380 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1644511149
transform 1 0 2484 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1644511149
transform 1 0 1380 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1644511149
transform 1 0 3496 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1644511149
transform 1 0 1380 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1644511149
transform 1 0 2116 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1644511149
transform 1 0 1380 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1644511149
transform 1 0 2116 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1644511149
transform 1 0 2852 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1644511149
transform 1 0 3772 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1644511149
transform 1 0 2576 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1644511149
transform 1 0 2116 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1644511149
transform 1 0 3772 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1644511149
transform 1 0 2484 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1644511149
transform 1 0 2484 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1644511149
transform 1 0 1380 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1644511149
transform 1 0 2484 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1644511149
transform 1 0 1380 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1644511149
transform 1 0 2116 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1644511149
transform 1 0 2116 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1644511149
transform 1 0 2852 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1644511149
transform 1 0 2668 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1644511149
transform 1 0 3680 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1644511149
transform 1 0 3496 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1644511149
transform 1 0 2116 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1644511149
transform 1 0 3220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1644511149
transform 1 0 3220 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1644511149
transform 1 0 3956 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1644511149
transform 1 0 3680 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1644511149
transform 1 0 3128 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1644511149
transform 1 0 4600 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1644511149
transform 1 0 4416 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1644511149
transform 1 0 3220 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1644511149
transform 1 0 2760 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1644511149
transform 1 0 2116 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1644511149
transform 1 0 3772 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1644511149
transform 1 0 2944 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1644511149
transform 1 0 4600 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1644511149
transform 1 0 2852 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1644511149
transform 1 0 2116 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1644511149
transform 1 0 2852 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1644511149
transform 1 0 2116 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1644511149
transform 1 0 2852 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1644511149
transform 1 0 2392 0 1 34816
box -38 -48 406 592
<< labels >>
rlabel metal4 s 2576 2128 2896 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 5840 2128 6160 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 9104 2128 9424 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 4208 2128 4528 77840 6 vssd1
port 1 nsew ground input
rlabel metal4 s 7472 2128 7792 77840 6 vssd1
port 1 nsew ground input
rlabel metal2 s 5998 0 6054 800 6 wb_clk_i
port 2 nsew signal input
rlabel metal2 s 5998 79200 6054 80000 6 wb_rst_i
port 3 nsew signal input
rlabel metal3 s 11200 79432 12000 79552 6 wbm_a_ack_i
port 4 nsew signal input
rlabel metal3 s 11200 5584 12000 5704 6 wbm_a_adr_o[0]
port 5 nsew signal tristate
rlabel metal3 s 11200 13336 12000 13456 6 wbm_a_adr_o[10]
port 6 nsew signal tristate
rlabel metal3 s 11200 14016 12000 14136 6 wbm_a_adr_o[11]
port 7 nsew signal tristate
rlabel metal3 s 11200 14832 12000 14952 6 wbm_a_adr_o[12]
port 8 nsew signal tristate
rlabel metal3 s 11200 15648 12000 15768 6 wbm_a_adr_o[13]
port 9 nsew signal tristate
rlabel metal3 s 11200 16328 12000 16448 6 wbm_a_adr_o[14]
port 10 nsew signal tristate
rlabel metal3 s 11200 17144 12000 17264 6 wbm_a_adr_o[15]
port 11 nsew signal tristate
rlabel metal3 s 11200 17960 12000 18080 6 wbm_a_adr_o[16]
port 12 nsew signal tristate
rlabel metal3 s 11200 18640 12000 18760 6 wbm_a_adr_o[17]
port 13 nsew signal tristate
rlabel metal3 s 11200 19456 12000 19576 6 wbm_a_adr_o[18]
port 14 nsew signal tristate
rlabel metal3 s 11200 20272 12000 20392 6 wbm_a_adr_o[19]
port 15 nsew signal tristate
rlabel metal3 s 11200 6400 12000 6520 6 wbm_a_adr_o[1]
port 16 nsew signal tristate
rlabel metal3 s 11200 20952 12000 21072 6 wbm_a_adr_o[20]
port 17 nsew signal tristate
rlabel metal3 s 11200 21768 12000 21888 6 wbm_a_adr_o[21]
port 18 nsew signal tristate
rlabel metal3 s 11200 22448 12000 22568 6 wbm_a_adr_o[22]
port 19 nsew signal tristate
rlabel metal3 s 11200 23264 12000 23384 6 wbm_a_adr_o[23]
port 20 nsew signal tristate
rlabel metal3 s 11200 24080 12000 24200 6 wbm_a_adr_o[24]
port 21 nsew signal tristate
rlabel metal3 s 11200 24760 12000 24880 6 wbm_a_adr_o[25]
port 22 nsew signal tristate
rlabel metal3 s 11200 25576 12000 25696 6 wbm_a_adr_o[26]
port 23 nsew signal tristate
rlabel metal3 s 11200 26392 12000 26512 6 wbm_a_adr_o[27]
port 24 nsew signal tristate
rlabel metal3 s 11200 27072 12000 27192 6 wbm_a_adr_o[28]
port 25 nsew signal tristate
rlabel metal3 s 11200 27888 12000 28008 6 wbm_a_adr_o[29]
port 26 nsew signal tristate
rlabel metal3 s 11200 7080 12000 7200 6 wbm_a_adr_o[2]
port 27 nsew signal tristate
rlabel metal3 s 11200 28704 12000 28824 6 wbm_a_adr_o[30]
port 28 nsew signal tristate
rlabel metal3 s 11200 29384 12000 29504 6 wbm_a_adr_o[31]
port 29 nsew signal tristate
rlabel metal3 s 11200 7896 12000 8016 6 wbm_a_adr_o[3]
port 30 nsew signal tristate
rlabel metal3 s 11200 8712 12000 8832 6 wbm_a_adr_o[4]
port 31 nsew signal tristate
rlabel metal3 s 11200 9392 12000 9512 6 wbm_a_adr_o[5]
port 32 nsew signal tristate
rlabel metal3 s 11200 10208 12000 10328 6 wbm_a_adr_o[6]
port 33 nsew signal tristate
rlabel metal3 s 11200 11024 12000 11144 6 wbm_a_adr_o[7]
port 34 nsew signal tristate
rlabel metal3 s 11200 11704 12000 11824 6 wbm_a_adr_o[8]
port 35 nsew signal tristate
rlabel metal3 s 11200 12520 12000 12640 6 wbm_a_adr_o[9]
port 36 nsew signal tristate
rlabel metal3 s 11200 960 12000 1080 6 wbm_a_cyc_o
port 37 nsew signal tristate
rlabel metal3 s 11200 54816 12000 54936 6 wbm_a_dat_i[0]
port 38 nsew signal input
rlabel metal3 s 11200 62432 12000 62552 6 wbm_a_dat_i[10]
port 39 nsew signal input
rlabel metal3 s 11200 63248 12000 63368 6 wbm_a_dat_i[11]
port 40 nsew signal input
rlabel metal3 s 11200 64064 12000 64184 6 wbm_a_dat_i[12]
port 41 nsew signal input
rlabel metal3 s 11200 64744 12000 64864 6 wbm_a_dat_i[13]
port 42 nsew signal input
rlabel metal3 s 11200 65560 12000 65680 6 wbm_a_dat_i[14]
port 43 nsew signal input
rlabel metal3 s 11200 66376 12000 66496 6 wbm_a_dat_i[15]
port 44 nsew signal input
rlabel metal3 s 11200 67056 12000 67176 6 wbm_a_dat_i[16]
port 45 nsew signal input
rlabel metal3 s 11200 67872 12000 67992 6 wbm_a_dat_i[17]
port 46 nsew signal input
rlabel metal3 s 11200 68688 12000 68808 6 wbm_a_dat_i[18]
port 47 nsew signal input
rlabel metal3 s 11200 69368 12000 69488 6 wbm_a_dat_i[19]
port 48 nsew signal input
rlabel metal3 s 11200 55632 12000 55752 6 wbm_a_dat_i[1]
port 49 nsew signal input
rlabel metal3 s 11200 70184 12000 70304 6 wbm_a_dat_i[20]
port 50 nsew signal input
rlabel metal3 s 11200 71000 12000 71120 6 wbm_a_dat_i[21]
port 51 nsew signal input
rlabel metal3 s 11200 71680 12000 71800 6 wbm_a_dat_i[22]
port 52 nsew signal input
rlabel metal3 s 11200 72496 12000 72616 6 wbm_a_dat_i[23]
port 53 nsew signal input
rlabel metal3 s 11200 73312 12000 73432 6 wbm_a_dat_i[24]
port 54 nsew signal input
rlabel metal3 s 11200 73992 12000 74112 6 wbm_a_dat_i[25]
port 55 nsew signal input
rlabel metal3 s 11200 74808 12000 74928 6 wbm_a_dat_i[26]
port 56 nsew signal input
rlabel metal3 s 11200 75624 12000 75744 6 wbm_a_dat_i[27]
port 57 nsew signal input
rlabel metal3 s 11200 76304 12000 76424 6 wbm_a_dat_i[28]
port 58 nsew signal input
rlabel metal3 s 11200 77120 12000 77240 6 wbm_a_dat_i[29]
port 59 nsew signal input
rlabel metal3 s 11200 56312 12000 56432 6 wbm_a_dat_i[2]
port 60 nsew signal input
rlabel metal3 s 11200 77936 12000 78056 6 wbm_a_dat_i[30]
port 61 nsew signal input
rlabel metal3 s 11200 78616 12000 78736 6 wbm_a_dat_i[31]
port 62 nsew signal input
rlabel metal3 s 11200 57128 12000 57248 6 wbm_a_dat_i[3]
port 63 nsew signal input
rlabel metal3 s 11200 57944 12000 58064 6 wbm_a_dat_i[4]
port 64 nsew signal input
rlabel metal3 s 11200 58624 12000 58744 6 wbm_a_dat_i[5]
port 65 nsew signal input
rlabel metal3 s 11200 59440 12000 59560 6 wbm_a_dat_i[6]
port 66 nsew signal input
rlabel metal3 s 11200 60256 12000 60376 6 wbm_a_dat_i[7]
port 67 nsew signal input
rlabel metal3 s 11200 60936 12000 61056 6 wbm_a_dat_i[8]
port 68 nsew signal input
rlabel metal3 s 11200 61752 12000 61872 6 wbm_a_dat_i[9]
port 69 nsew signal input
rlabel metal3 s 11200 30200 12000 30320 6 wbm_a_dat_o[0]
port 70 nsew signal tristate
rlabel metal3 s 11200 37952 12000 38072 6 wbm_a_dat_o[10]
port 71 nsew signal tristate
rlabel metal3 s 11200 38632 12000 38752 6 wbm_a_dat_o[11]
port 72 nsew signal tristate
rlabel metal3 s 11200 39448 12000 39568 6 wbm_a_dat_o[12]
port 73 nsew signal tristate
rlabel metal3 s 11200 40264 12000 40384 6 wbm_a_dat_o[13]
port 74 nsew signal tristate
rlabel metal3 s 11200 40944 12000 41064 6 wbm_a_dat_o[14]
port 75 nsew signal tristate
rlabel metal3 s 11200 41760 12000 41880 6 wbm_a_dat_o[15]
port 76 nsew signal tristate
rlabel metal3 s 11200 42440 12000 42560 6 wbm_a_dat_o[16]
port 77 nsew signal tristate
rlabel metal3 s 11200 43256 12000 43376 6 wbm_a_dat_o[17]
port 78 nsew signal tristate
rlabel metal3 s 11200 44072 12000 44192 6 wbm_a_dat_o[18]
port 79 nsew signal tristate
rlabel metal3 s 11200 44752 12000 44872 6 wbm_a_dat_o[19]
port 80 nsew signal tristate
rlabel metal3 s 11200 31016 12000 31136 6 wbm_a_dat_o[1]
port 81 nsew signal tristate
rlabel metal3 s 11200 45568 12000 45688 6 wbm_a_dat_o[20]
port 82 nsew signal tristate
rlabel metal3 s 11200 46384 12000 46504 6 wbm_a_dat_o[21]
port 83 nsew signal tristate
rlabel metal3 s 11200 47064 12000 47184 6 wbm_a_dat_o[22]
port 84 nsew signal tristate
rlabel metal3 s 11200 47880 12000 48000 6 wbm_a_dat_o[23]
port 85 nsew signal tristate
rlabel metal3 s 11200 48696 12000 48816 6 wbm_a_dat_o[24]
port 86 nsew signal tristate
rlabel metal3 s 11200 49376 12000 49496 6 wbm_a_dat_o[25]
port 87 nsew signal tristate
rlabel metal3 s 11200 50192 12000 50312 6 wbm_a_dat_o[26]
port 88 nsew signal tristate
rlabel metal3 s 11200 51008 12000 51128 6 wbm_a_dat_o[27]
port 89 nsew signal tristate
rlabel metal3 s 11200 51688 12000 51808 6 wbm_a_dat_o[28]
port 90 nsew signal tristate
rlabel metal3 s 11200 52504 12000 52624 6 wbm_a_dat_o[29]
port 91 nsew signal tristate
rlabel metal3 s 11200 31696 12000 31816 6 wbm_a_dat_o[2]
port 92 nsew signal tristate
rlabel metal3 s 11200 53320 12000 53440 6 wbm_a_dat_o[30]
port 93 nsew signal tristate
rlabel metal3 s 11200 54000 12000 54120 6 wbm_a_dat_o[31]
port 94 nsew signal tristate
rlabel metal3 s 11200 32512 12000 32632 6 wbm_a_dat_o[3]
port 95 nsew signal tristate
rlabel metal3 s 11200 33328 12000 33448 6 wbm_a_dat_o[4]
port 96 nsew signal tristate
rlabel metal3 s 11200 34008 12000 34128 6 wbm_a_dat_o[5]
port 97 nsew signal tristate
rlabel metal3 s 11200 34824 12000 34944 6 wbm_a_dat_o[6]
port 98 nsew signal tristate
rlabel metal3 s 11200 35640 12000 35760 6 wbm_a_dat_o[7]
port 99 nsew signal tristate
rlabel metal3 s 11200 36320 12000 36440 6 wbm_a_dat_o[8]
port 100 nsew signal tristate
rlabel metal3 s 11200 37136 12000 37256 6 wbm_a_dat_o[9]
port 101 nsew signal tristate
rlabel metal3 s 11200 2456 12000 2576 6 wbm_a_sel_o[0]
port 102 nsew signal tristate
rlabel metal3 s 11200 3272 12000 3392 6 wbm_a_sel_o[1]
port 103 nsew signal tristate
rlabel metal3 s 11200 4088 12000 4208 6 wbm_a_sel_o[2]
port 104 nsew signal tristate
rlabel metal3 s 11200 4768 12000 4888 6 wbm_a_sel_o[3]
port 105 nsew signal tristate
rlabel metal3 s 11200 280 12000 400 6 wbm_a_stb_o
port 106 nsew signal tristate
rlabel metal3 s 11200 1776 12000 1896 6 wbm_a_we_o
port 107 nsew signal tristate
rlabel metal3 s 0 79568 800 79688 6 wbm_b_ack_i
port 108 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 wbm_b_adr_o[0]
port 109 nsew signal tristate
rlabel metal3 s 0 51824 800 51944 6 wbm_b_adr_o[10]
port 110 nsew signal tristate
rlabel metal3 s 0 48016 800 48136 6 wbm_b_adr_o[1]
port 111 nsew signal tristate
rlabel metal3 s 0 48424 800 48544 6 wbm_b_adr_o[2]
port 112 nsew signal tristate
rlabel metal3 s 0 48832 800 48952 6 wbm_b_adr_o[3]
port 113 nsew signal tristate
rlabel metal3 s 0 49240 800 49360 6 wbm_b_adr_o[4]
port 114 nsew signal tristate
rlabel metal3 s 0 49648 800 49768 6 wbm_b_adr_o[5]
port 115 nsew signal tristate
rlabel metal3 s 0 50056 800 50176 6 wbm_b_adr_o[6]
port 116 nsew signal tristate
rlabel metal3 s 0 50600 800 50720 6 wbm_b_adr_o[7]
port 117 nsew signal tristate
rlabel metal3 s 0 51008 800 51128 6 wbm_b_adr_o[8]
port 118 nsew signal tristate
rlabel metal3 s 0 51416 800 51536 6 wbm_b_adr_o[9]
port 119 nsew signal tristate
rlabel metal3 s 0 45024 800 45144 6 wbm_b_cyc_o
port 120 nsew signal tristate
rlabel metal3 s 0 65968 800 66088 6 wbm_b_dat_i[0]
port 121 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 wbm_b_dat_i[10]
port 122 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 wbm_b_dat_i[11]
port 123 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 wbm_b_dat_i[12]
port 124 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 wbm_b_dat_i[13]
port 125 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 wbm_b_dat_i[14]
port 126 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 wbm_b_dat_i[15]
port 127 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 wbm_b_dat_i[16]
port 128 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 wbm_b_dat_i[17]
port 129 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 wbm_b_dat_i[18]
port 130 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 wbm_b_dat_i[19]
port 131 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 wbm_b_dat_i[1]
port 132 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 wbm_b_dat_i[20]
port 133 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 wbm_b_dat_i[21]
port 134 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 wbm_b_dat_i[22]
port 135 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 wbm_b_dat_i[23]
port 136 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 wbm_b_dat_i[24]
port 137 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 wbm_b_dat_i[25]
port 138 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 wbm_b_dat_i[26]
port 139 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 wbm_b_dat_i[27]
port 140 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 wbm_b_dat_i[28]
port 141 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 wbm_b_dat_i[29]
port 142 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 wbm_b_dat_i[2]
port 143 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 wbm_b_dat_i[30]
port 144 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 wbm_b_dat_i[31]
port 145 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 wbm_b_dat_i[3]
port 146 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 wbm_b_dat_i[4]
port 147 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 wbm_b_dat_i[5]
port 148 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 wbm_b_dat_i[6]
port 149 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 wbm_b_dat_i[7]
port 150 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 wbm_b_dat_i[8]
port 151 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 wbm_b_dat_i[9]
port 152 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 wbm_b_dat_o[0]
port 153 nsew signal tristate
rlabel metal3 s 0 56584 800 56704 6 wbm_b_dat_o[10]
port 154 nsew signal tristate
rlabel metal3 s 0 56992 800 57112 6 wbm_b_dat_o[11]
port 155 nsew signal tristate
rlabel metal3 s 0 57400 800 57520 6 wbm_b_dat_o[12]
port 156 nsew signal tristate
rlabel metal3 s 0 57808 800 57928 6 wbm_b_dat_o[13]
port 157 nsew signal tristate
rlabel metal3 s 0 58216 800 58336 6 wbm_b_dat_o[14]
port 158 nsew signal tristate
rlabel metal3 s 0 58624 800 58744 6 wbm_b_dat_o[15]
port 159 nsew signal tristate
rlabel metal3 s 0 59032 800 59152 6 wbm_b_dat_o[16]
port 160 nsew signal tristate
rlabel metal3 s 0 59576 800 59696 6 wbm_b_dat_o[17]
port 161 nsew signal tristate
rlabel metal3 s 0 59984 800 60104 6 wbm_b_dat_o[18]
port 162 nsew signal tristate
rlabel metal3 s 0 60392 800 60512 6 wbm_b_dat_o[19]
port 163 nsew signal tristate
rlabel metal3 s 0 52640 800 52760 6 wbm_b_dat_o[1]
port 164 nsew signal tristate
rlabel metal3 s 0 60800 800 60920 6 wbm_b_dat_o[20]
port 165 nsew signal tristate
rlabel metal3 s 0 61208 800 61328 6 wbm_b_dat_o[21]
port 166 nsew signal tristate
rlabel metal3 s 0 61616 800 61736 6 wbm_b_dat_o[22]
port 167 nsew signal tristate
rlabel metal3 s 0 62024 800 62144 6 wbm_b_dat_o[23]
port 168 nsew signal tristate
rlabel metal3 s 0 62568 800 62688 6 wbm_b_dat_o[24]
port 169 nsew signal tristate
rlabel metal3 s 0 62976 800 63096 6 wbm_b_dat_o[25]
port 170 nsew signal tristate
rlabel metal3 s 0 63384 800 63504 6 wbm_b_dat_o[26]
port 171 nsew signal tristate
rlabel metal3 s 0 63792 800 63912 6 wbm_b_dat_o[27]
port 172 nsew signal tristate
rlabel metal3 s 0 64200 800 64320 6 wbm_b_dat_o[28]
port 173 nsew signal tristate
rlabel metal3 s 0 64608 800 64728 6 wbm_b_dat_o[29]
port 174 nsew signal tristate
rlabel metal3 s 0 53048 800 53168 6 wbm_b_dat_o[2]
port 175 nsew signal tristate
rlabel metal3 s 0 65016 800 65136 6 wbm_b_dat_o[30]
port 176 nsew signal tristate
rlabel metal3 s 0 65560 800 65680 6 wbm_b_dat_o[31]
port 177 nsew signal tristate
rlabel metal3 s 0 53592 800 53712 6 wbm_b_dat_o[3]
port 178 nsew signal tristate
rlabel metal3 s 0 54000 800 54120 6 wbm_b_dat_o[4]
port 179 nsew signal tristate
rlabel metal3 s 0 54408 800 54528 6 wbm_b_dat_o[5]
port 180 nsew signal tristate
rlabel metal3 s 0 54816 800 54936 6 wbm_b_dat_o[6]
port 181 nsew signal tristate
rlabel metal3 s 0 55224 800 55344 6 wbm_b_dat_o[7]
port 182 nsew signal tristate
rlabel metal3 s 0 55632 800 55752 6 wbm_b_dat_o[8]
port 183 nsew signal tristate
rlabel metal3 s 0 56040 800 56160 6 wbm_b_dat_o[9]
port 184 nsew signal tristate
rlabel metal3 s 0 45840 800 45960 6 wbm_b_sel_o[0]
port 185 nsew signal tristate
rlabel metal3 s 0 46248 800 46368 6 wbm_b_sel_o[1]
port 186 nsew signal tristate
rlabel metal3 s 0 46656 800 46776 6 wbm_b_sel_o[2]
port 187 nsew signal tristate
rlabel metal3 s 0 47064 800 47184 6 wbm_b_sel_o[3]
port 188 nsew signal tristate
rlabel metal3 s 0 44616 800 44736 6 wbm_b_stb_o
port 189 nsew signal tristate
rlabel metal3 s 0 45432 800 45552 6 wbm_b_we_o
port 190 nsew signal tristate
rlabel metal3 s 0 44072 800 44192 6 wbs_ack_o
port 191 nsew signal tristate
rlabel metal3 s 0 3136 800 3256 6 wbs_adr_i[0]
port 192 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 wbs_adr_i[10]
port 193 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 wbs_adr_i[11]
port 194 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 wbs_adr_i[12]
port 195 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 wbs_adr_i[13]
port 196 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 wbs_adr_i[14]
port 197 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wbs_adr_i[15]
port 198 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 wbs_adr_i[16]
port 199 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 wbs_adr_i[17]
port 200 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 wbs_adr_i[18]
port 201 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 wbs_adr_i[19]
port 202 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 wbs_adr_i[1]
port 203 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_adr_i[20]
port 204 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 wbs_adr_i[21]
port 205 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 wbs_adr_i[22]
port 206 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 wbs_adr_i[23]
port 207 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 wbs_adr_i[24]
port 208 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 wbs_adr_i[25]
port 209 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 wbs_adr_i[26]
port 210 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 wbs_adr_i[27]
port 211 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 wbs_adr_i[28]
port 212 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 wbs_adr_i[29]
port 213 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 wbs_adr_i[2]
port 214 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 wbs_adr_i[30]
port 215 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 wbs_adr_i[31]
port 216 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 wbs_adr_i[3]
port 217 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 wbs_adr_i[4]
port 218 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 wbs_adr_i[5]
port 219 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 wbs_adr_i[6]
port 220 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wbs_adr_i[7]
port 221 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 wbs_adr_i[8]
port 222 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 wbs_adr_i[9]
port 223 nsew signal input
rlabel metal3 s 0 552 800 672 6 wbs_cyc_i
port 224 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 wbs_dat_i[0]
port 225 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 wbs_dat_i[10]
port 226 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 wbs_dat_i[11]
port 227 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 wbs_dat_i[12]
port 228 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 wbs_dat_i[13]
port 229 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 wbs_dat_i[14]
port 230 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wbs_dat_i[15]
port 231 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 wbs_dat_i[16]
port 232 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 wbs_dat_i[17]
port 233 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 wbs_dat_i[18]
port 234 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 wbs_dat_i[19]
port 235 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 wbs_dat_i[1]
port 236 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 wbs_dat_i[20]
port 237 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wbs_dat_i[21]
port 238 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 wbs_dat_i[22]
port 239 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 wbs_dat_i[23]
port 240 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 wbs_dat_i[24]
port 241 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 wbs_dat_i[25]
port 242 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 wbs_dat_i[26]
port 243 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 wbs_dat_i[27]
port 244 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 wbs_dat_i[28]
port 245 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 wbs_dat_i[29]
port 246 nsew signal input
rlabel metal3 s 0 17552 800 17672 6 wbs_dat_i[2]
port 247 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 wbs_dat_i[30]
port 248 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 wbs_dat_i[31]
port 249 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wbs_dat_i[3]
port 250 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 wbs_dat_i[4]
port 251 nsew signal input
rlabel metal3 s 0 18912 800 19032 6 wbs_dat_i[5]
port 252 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 wbs_dat_i[6]
port 253 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 wbs_dat_i[7]
port 254 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 wbs_dat_i[8]
port 255 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 wbs_dat_i[9]
port 256 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 wbs_dat_o[0]
port 257 nsew signal tristate
rlabel metal3 s 0 34688 800 34808 6 wbs_dat_o[10]
port 258 nsew signal tristate
rlabel metal3 s 0 35096 800 35216 6 wbs_dat_o[11]
port 259 nsew signal tristate
rlabel metal3 s 0 35504 800 35624 6 wbs_dat_o[12]
port 260 nsew signal tristate
rlabel metal3 s 0 36048 800 36168 6 wbs_dat_o[13]
port 261 nsew signal tristate
rlabel metal3 s 0 36456 800 36576 6 wbs_dat_o[14]
port 262 nsew signal tristate
rlabel metal3 s 0 36864 800 36984 6 wbs_dat_o[15]
port 263 nsew signal tristate
rlabel metal3 s 0 37272 800 37392 6 wbs_dat_o[16]
port 264 nsew signal tristate
rlabel metal3 s 0 37680 800 37800 6 wbs_dat_o[17]
port 265 nsew signal tristate
rlabel metal3 s 0 38088 800 38208 6 wbs_dat_o[18]
port 266 nsew signal tristate
rlabel metal3 s 0 38496 800 38616 6 wbs_dat_o[19]
port 267 nsew signal tristate
rlabel metal3 s 0 30880 800 31000 6 wbs_dat_o[1]
port 268 nsew signal tristate
rlabel metal3 s 0 39040 800 39160 6 wbs_dat_o[20]
port 269 nsew signal tristate
rlabel metal3 s 0 39448 800 39568 6 wbs_dat_o[21]
port 270 nsew signal tristate
rlabel metal3 s 0 39856 800 39976 6 wbs_dat_o[22]
port 271 nsew signal tristate
rlabel metal3 s 0 40264 800 40384 6 wbs_dat_o[23]
port 272 nsew signal tristate
rlabel metal3 s 0 40672 800 40792 6 wbs_dat_o[24]
port 273 nsew signal tristate
rlabel metal3 s 0 41080 800 41200 6 wbs_dat_o[25]
port 274 nsew signal tristate
rlabel metal3 s 0 41624 800 41744 6 wbs_dat_o[26]
port 275 nsew signal tristate
rlabel metal3 s 0 42032 800 42152 6 wbs_dat_o[27]
port 276 nsew signal tristate
rlabel metal3 s 0 42440 800 42560 6 wbs_dat_o[28]
port 277 nsew signal tristate
rlabel metal3 s 0 42848 800 42968 6 wbs_dat_o[29]
port 278 nsew signal tristate
rlabel metal3 s 0 31288 800 31408 6 wbs_dat_o[2]
port 279 nsew signal tristate
rlabel metal3 s 0 43256 800 43376 6 wbs_dat_o[30]
port 280 nsew signal tristate
rlabel metal3 s 0 43664 800 43784 6 wbs_dat_o[31]
port 281 nsew signal tristate
rlabel metal3 s 0 31696 800 31816 6 wbs_dat_o[3]
port 282 nsew signal tristate
rlabel metal3 s 0 32104 800 32224 6 wbs_dat_o[4]
port 283 nsew signal tristate
rlabel metal3 s 0 32512 800 32632 6 wbs_dat_o[5]
port 284 nsew signal tristate
rlabel metal3 s 0 33056 800 33176 6 wbs_dat_o[6]
port 285 nsew signal tristate
rlabel metal3 s 0 33464 800 33584 6 wbs_dat_o[7]
port 286 nsew signal tristate
rlabel metal3 s 0 33872 800 33992 6 wbs_dat_o[8]
port 287 nsew signal tristate
rlabel metal3 s 0 34280 800 34400 6 wbs_dat_o[9]
port 288 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 wbs_sel_i[0]
port 289 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 wbs_sel_i[1]
port 290 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wbs_sel_i[2]
port 291 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 wbs_sel_i[3]
port 292 nsew signal input
rlabel metal3 s 0 144 800 264 6 wbs_stb_i
port 293 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wbs_we_i
port 294 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12000 80000
<< end >>
