magic
tech sky130A
magscale 1 2
timestamp 1647558355
<< viali >>
rect 1409 77537 1443 77571
rect 10149 77537 10183 77571
rect 1685 77469 1719 77503
rect 2881 77469 2915 77503
rect 3985 77469 4019 77503
rect 4629 77469 4663 77503
rect 9413 77469 9447 77503
rect 9965 77469 9999 77503
rect 2697 77333 2731 77367
rect 3801 77333 3835 77367
rect 4445 77333 4479 77367
rect 9229 77333 9263 77367
rect 1409 76993 1443 77027
rect 2329 76993 2363 77027
rect 2973 76993 3007 77027
rect 3617 76993 3651 77027
rect 4261 76993 4295 77027
rect 9413 76993 9447 77027
rect 9873 76993 9907 77027
rect 9229 76857 9263 76891
rect 1593 76789 1627 76823
rect 2145 76789 2179 76823
rect 2789 76789 2823 76823
rect 3433 76789 3467 76823
rect 4077 76789 4111 76823
rect 10057 76789 10091 76823
rect 9965 76585 9999 76619
rect 1961 76517 1995 76551
rect 3065 76517 3099 76551
rect 1409 76381 1443 76415
rect 1593 76381 1627 76415
rect 1829 76381 1863 76415
rect 2513 76381 2547 76415
rect 2886 76381 2920 76415
rect 10149 76381 10183 76415
rect 1685 76313 1719 76347
rect 2697 76313 2731 76347
rect 2789 76313 2823 76347
rect 1409 76041 1443 76075
rect 9965 76041 9999 76075
rect 2605 75973 2639 76007
rect 2898 75973 2932 76007
rect 1593 75905 1627 75939
rect 2329 75905 2363 75939
rect 2513 75905 2547 75939
rect 2702 75905 2736 75939
rect 3617 75905 3651 75939
rect 10149 75905 10183 75939
rect 3433 75701 3467 75735
rect 3065 75497 3099 75531
rect 2513 75429 2547 75463
rect 9965 75429 9999 75463
rect 1961 75293 1995 75327
rect 2237 75293 2271 75327
rect 2357 75293 2391 75327
rect 3249 75293 3283 75327
rect 10149 75293 10183 75327
rect 2145 75225 2179 75259
rect 1593 74885 1627 74919
rect 1685 74885 1719 74919
rect 1409 74817 1443 74851
rect 1829 74817 1863 74851
rect 2697 74817 2731 74851
rect 2513 74681 2547 74715
rect 1961 74613 1995 74647
rect 2513 74341 2547 74375
rect 9965 74341 9999 74375
rect 1961 74205 1995 74239
rect 2381 74205 2415 74239
rect 3249 74205 3283 74239
rect 10149 74205 10183 74239
rect 2145 74137 2179 74171
rect 2237 74137 2271 74171
rect 3065 74069 3099 74103
rect 1593 73729 1627 73763
rect 2237 73729 2271 73763
rect 10149 73729 10183 73763
rect 1409 73593 1443 73627
rect 2053 73525 2087 73559
rect 9965 73525 9999 73559
rect 1409 73117 1443 73151
rect 1593 73117 1627 73151
rect 1829 73117 1863 73151
rect 1685 73049 1719 73083
rect 1978 72981 2012 73015
rect 1593 72641 1627 72675
rect 2237 72641 2271 72675
rect 2881 72641 2915 72675
rect 10149 72641 10183 72675
rect 2053 72505 2087 72539
rect 1409 72437 1443 72471
rect 2697 72437 2731 72471
rect 9965 72437 9999 72471
rect 9965 72233 9999 72267
rect 2605 72165 2639 72199
rect 1593 72029 1627 72063
rect 2053 72029 2087 72063
rect 2237 72029 2271 72063
rect 2329 72029 2363 72063
rect 2473 72029 2507 72063
rect 10149 72029 10183 72063
rect 1409 71893 1443 71927
rect 1685 71621 1719 71655
rect 2789 71621 2823 71655
rect 1409 71553 1443 71587
rect 1593 71553 1627 71587
rect 1829 71553 1863 71587
rect 2513 71553 2547 71587
rect 2697 71553 2731 71587
rect 2886 71553 2920 71587
rect 10149 71553 10183 71587
rect 9965 71417 9999 71451
rect 1961 71349 1995 71383
rect 3065 71349 3099 71383
rect 1409 71077 1443 71111
rect 1593 70941 1627 70975
rect 2237 70941 2271 70975
rect 2053 70805 2087 70839
rect 9965 70601 9999 70635
rect 1685 70533 1719 70567
rect 1409 70465 1443 70499
rect 1593 70465 1627 70499
rect 1829 70465 1863 70499
rect 10149 70465 10183 70499
rect 1961 70261 1995 70295
rect 1593 69853 1627 69887
rect 2237 69853 2271 69887
rect 10149 69853 10183 69887
rect 1409 69717 1443 69751
rect 2053 69717 2087 69751
rect 9965 69717 9999 69751
rect 1593 69377 1627 69411
rect 2237 69377 2271 69411
rect 1409 69173 1443 69207
rect 2053 69173 2087 69207
rect 1961 68969 1995 69003
rect 1409 68765 1443 68799
rect 1685 68765 1719 68799
rect 1829 68765 1863 68799
rect 2697 68765 2731 68799
rect 10149 68765 10183 68799
rect 1593 68697 1627 68731
rect 2513 68629 2547 68663
rect 9965 68629 9999 68663
rect 1593 68357 1627 68391
rect 1685 68357 1719 68391
rect 1409 68289 1443 68323
rect 1829 68289 1863 68323
rect 2697 68289 2731 68323
rect 10149 68289 10183 68323
rect 1961 68153 1995 68187
rect 2513 68085 2547 68119
rect 9965 68085 9999 68119
rect 1409 67813 1443 67847
rect 2789 67813 2823 67847
rect 1593 67677 1627 67711
rect 2237 67677 2271 67711
rect 2513 67677 2547 67711
rect 2657 67677 2691 67711
rect 2421 67609 2455 67643
rect 9965 67337 9999 67371
rect 2881 67269 2915 67303
rect 2697 67201 2731 67235
rect 2973 67201 3007 67235
rect 3117 67201 3151 67235
rect 10149 67201 10183 67235
rect 1409 67133 1443 67167
rect 1685 67133 1719 67167
rect 3249 66997 3283 67031
rect 9965 66793 9999 66827
rect 1685 66657 1719 66691
rect 3065 66657 3099 66691
rect 1409 66589 1443 66623
rect 2789 66589 2823 66623
rect 10149 66589 10183 66623
rect 2881 66181 2915 66215
rect 2973 66181 3007 66215
rect 1685 66113 1719 66147
rect 2697 66113 2731 66147
rect 3117 66113 3151 66147
rect 10149 66113 10183 66147
rect 1409 66045 1443 66079
rect 3249 65909 3283 65943
rect 9965 65909 9999 65943
rect 1409 65569 1443 65603
rect 2973 65569 3007 65603
rect 1685 65501 1719 65535
rect 2697 65501 2731 65535
rect 3801 65501 3835 65535
rect 3985 65365 4019 65399
rect 1409 65025 1443 65059
rect 2145 65025 2179 65059
rect 2881 65025 2915 65059
rect 3617 65025 3651 65059
rect 10149 65025 10183 65059
rect 1593 64889 1627 64923
rect 2329 64889 2363 64923
rect 3065 64889 3099 64923
rect 3801 64889 3835 64923
rect 9965 64889 9999 64923
rect 2513 64549 2547 64583
rect 1961 64413 1995 64447
rect 2237 64413 2271 64447
rect 2381 64413 2415 64447
rect 10149 64413 10183 64447
rect 2145 64345 2179 64379
rect 9965 64277 9999 64311
rect 2234 64005 2268 64039
rect 1961 63937 1995 63971
rect 2145 63937 2179 63971
rect 2381 63937 2415 63971
rect 2513 63733 2547 63767
rect 2513 63461 2547 63495
rect 1961 63325 1995 63359
rect 2237 63325 2271 63359
rect 2381 63325 2415 63359
rect 3801 63325 3835 63359
rect 9321 63325 9355 63359
rect 9597 63325 9631 63359
rect 2145 63257 2179 63291
rect 3985 63189 4019 63223
rect 1685 62917 1719 62951
rect 2789 62917 2823 62951
rect 1409 62849 1443 62883
rect 1593 62849 1627 62883
rect 1829 62849 1863 62883
rect 2513 62849 2547 62883
rect 2697 62849 2731 62883
rect 2881 62849 2915 62883
rect 3525 62849 3559 62883
rect 10149 62849 10183 62883
rect 3709 62713 3743 62747
rect 9965 62713 9999 62747
rect 1961 62645 1995 62679
rect 3065 62645 3099 62679
rect 1409 62237 1443 62271
rect 2145 62237 2179 62271
rect 2881 62237 2915 62271
rect 10149 62237 10183 62271
rect 1593 62101 1627 62135
rect 2329 62101 2363 62135
rect 3065 62101 3099 62135
rect 9965 62101 9999 62135
rect 1409 61761 1443 61795
rect 1593 61761 1627 61795
rect 1685 61761 1719 61795
rect 1829 61761 1863 61795
rect 1961 61557 1995 61591
rect 1409 61149 1443 61183
rect 2145 61149 2179 61183
rect 10149 61149 10183 61183
rect 1593 61013 1627 61047
rect 2329 61013 2363 61047
rect 9965 61013 9999 61047
rect 1593 60741 1627 60775
rect 1409 60673 1443 60707
rect 1685 60673 1719 60707
rect 1782 60673 1816 60707
rect 2513 60673 2547 60707
rect 10149 60673 10183 60707
rect 2697 60537 2731 60571
rect 1961 60469 1995 60503
rect 9965 60469 9999 60503
rect 2881 60265 2915 60299
rect 1409 60061 1443 60095
rect 2145 60061 2179 60095
rect 3065 60061 3099 60095
rect 1593 59925 1627 59959
rect 2329 59925 2363 59959
rect 1409 59585 1443 59619
rect 9597 59585 9631 59619
rect 9321 59517 9355 59551
rect 1593 59381 1627 59415
rect 1409 58973 1443 59007
rect 2145 58973 2179 59007
rect 2881 58973 2915 59007
rect 10149 58973 10183 59007
rect 1593 58837 1627 58871
rect 2329 58837 2363 58871
rect 3065 58837 3099 58871
rect 9965 58837 9999 58871
rect 2145 58565 2179 58599
rect 1869 58497 1903 58531
rect 2053 58497 2087 58531
rect 2289 58497 2323 58531
rect 10149 58497 10183 58531
rect 2421 58293 2455 58327
rect 9965 58293 9999 58327
rect 2881 57953 2915 57987
rect 1409 57885 1443 57919
rect 1685 57885 1719 57919
rect 1829 57885 1863 57919
rect 2697 57885 2731 57919
rect 1593 57817 1627 57851
rect 1969 57749 2003 57783
rect 2329 57545 2363 57579
rect 3617 57545 3651 57579
rect 1409 57409 1443 57443
rect 2145 57409 2179 57443
rect 2881 57409 2915 57443
rect 3801 57409 3835 57443
rect 9321 57341 9355 57375
rect 9597 57341 9631 57375
rect 1593 57205 1627 57239
rect 3065 57205 3099 57239
rect 2973 57001 3007 57035
rect 3801 57001 3835 57035
rect 1961 56933 1995 56967
rect 9597 56865 9631 56899
rect 1409 56797 1443 56831
rect 1829 56797 1863 56831
rect 2697 56797 2731 56831
rect 2789 56797 2823 56831
rect 3985 56797 4019 56831
rect 9321 56797 9355 56831
rect 1593 56729 1627 56763
rect 1685 56729 1719 56763
rect 2145 56457 2179 56491
rect 2881 56389 2915 56423
rect 1961 56321 1995 56355
rect 2605 56321 2639 56355
rect 3709 56321 3743 56355
rect 3893 56321 3927 56355
rect 10149 56321 10183 56355
rect 1777 56253 1811 56287
rect 3525 56253 3559 56287
rect 9965 56117 9999 56151
rect 1593 55913 1627 55947
rect 2789 55913 2823 55947
rect 4813 55845 4847 55879
rect 2421 55777 2455 55811
rect 9597 55777 9631 55811
rect 1409 55709 1443 55743
rect 2605 55709 2639 55743
rect 3893 55709 3927 55743
rect 3985 55709 4019 55743
rect 4629 55709 4663 55743
rect 9321 55709 9355 55743
rect 4169 55573 4203 55607
rect 3433 55369 3467 55403
rect 1593 55301 1627 55335
rect 1409 55233 1443 55267
rect 1682 55233 1716 55267
rect 1782 55233 1816 55267
rect 2513 55233 2547 55267
rect 3249 55233 3283 55267
rect 9321 55233 9355 55267
rect 1961 55029 1995 55063
rect 2697 55029 2731 55063
rect 9551 55029 9585 55063
rect 1409 54621 1443 54655
rect 1685 54621 1719 54655
rect 1777 54621 1811 54655
rect 2421 54621 2455 54655
rect 10149 54621 10183 54655
rect 1593 54553 1627 54587
rect 1961 54485 1995 54519
rect 2605 54485 2639 54519
rect 9965 54485 9999 54519
rect 2881 54281 2915 54315
rect 1409 54145 1443 54179
rect 2145 54145 2179 54179
rect 3065 54145 3099 54179
rect 9873 54145 9907 54179
rect 10057 54009 10091 54043
rect 1593 53941 1627 53975
rect 2329 53941 2363 53975
rect 1409 53533 1443 53567
rect 9873 53533 9907 53567
rect 1593 53397 1627 53431
rect 10057 53397 10091 53431
rect 2513 53193 2547 53227
rect 9229 53193 9263 53227
rect 1409 53057 1443 53091
rect 2329 53057 2363 53091
rect 3249 53057 3283 53091
rect 3433 53057 3467 53091
rect 9413 53057 9447 53091
rect 9873 53057 9907 53091
rect 2145 52989 2179 53023
rect 3065 52989 3099 53023
rect 1593 52853 1627 52887
rect 10057 52853 10091 52887
rect 2329 52581 2363 52615
rect 1409 52445 1443 52479
rect 2145 52445 2179 52479
rect 10149 52445 10183 52479
rect 1593 52309 1627 52343
rect 9965 52309 9999 52343
rect 2237 52105 2271 52139
rect 4077 52105 4111 52139
rect 1409 51969 1443 52003
rect 2421 51969 2455 52003
rect 3065 51969 3099 52003
rect 3893 51969 3927 52003
rect 9873 51969 9907 52003
rect 2881 51901 2915 51935
rect 3709 51901 3743 51935
rect 3249 51833 3283 51867
rect 1593 51765 1627 51799
rect 10057 51765 10091 51799
rect 2789 51561 2823 51595
rect 1409 51357 1443 51391
rect 2513 51357 2547 51391
rect 2605 51357 2639 51391
rect 9873 51357 9907 51391
rect 1593 51221 1627 51255
rect 10057 51221 10091 51255
rect 9965 51017 9999 51051
rect 1409 50881 1443 50915
rect 2145 50881 2179 50915
rect 10149 50881 10183 50915
rect 1593 50745 1627 50779
rect 2329 50745 2363 50779
rect 1409 50269 1443 50303
rect 1593 50269 1627 50303
rect 1777 50269 1811 50303
rect 2421 50269 2455 50303
rect 9873 50269 9907 50303
rect 1685 50201 1719 50235
rect 1961 50133 1995 50167
rect 2605 50133 2639 50167
rect 10057 50133 10091 50167
rect 3157 49929 3191 49963
rect 10057 49929 10091 49963
rect 1685 49861 1719 49895
rect 1409 49793 1443 49827
rect 1593 49793 1627 49827
rect 1777 49793 1811 49827
rect 2421 49793 2455 49827
rect 3341 49793 3375 49827
rect 9873 49793 9907 49827
rect 1961 49589 1995 49623
rect 2605 49589 2639 49623
rect 2789 49385 2823 49419
rect 1409 49181 1443 49215
rect 1593 49181 1627 49215
rect 1777 49181 1811 49215
rect 2421 49181 2455 49215
rect 2605 49181 2639 49215
rect 3801 49181 3835 49215
rect 9873 49181 9907 49215
rect 1685 49113 1719 49147
rect 1961 49045 1995 49079
rect 3985 49045 4019 49079
rect 10057 49045 10091 49079
rect 1961 48841 1995 48875
rect 3157 48841 3191 48875
rect 9965 48841 9999 48875
rect 1409 48705 1443 48739
rect 1593 48705 1627 48739
rect 1685 48705 1719 48739
rect 1777 48705 1811 48739
rect 2789 48705 2823 48739
rect 2973 48705 3007 48739
rect 3617 48705 3651 48739
rect 10149 48705 10183 48739
rect 3801 48501 3835 48535
rect 9229 48229 9263 48263
rect 2697 48161 2731 48195
rect 1409 48093 1443 48127
rect 2421 48093 2455 48127
rect 9413 48093 9447 48127
rect 9873 48093 9907 48127
rect 1593 47957 1627 47991
rect 10057 47957 10091 47991
rect 1409 47617 1443 47651
rect 2881 47617 2915 47651
rect 9873 47617 9907 47651
rect 2605 47549 2639 47583
rect 1593 47413 1627 47447
rect 10057 47413 10091 47447
rect 1961 47209 1995 47243
rect 2789 47209 2823 47243
rect 7757 47209 7791 47243
rect 9965 47209 9999 47243
rect 3985 47141 4019 47175
rect 5549 47073 5583 47107
rect 1685 47005 1719 47039
rect 1777 47005 1811 47039
rect 2513 47005 2547 47039
rect 2605 47005 2639 47039
rect 3801 47005 3835 47039
rect 4537 47005 4571 47039
rect 4721 47005 4755 47039
rect 5733 47005 5767 47039
rect 5917 47005 5951 47039
rect 7941 47005 7975 47039
rect 10149 47005 10183 47039
rect 4905 46937 4939 46971
rect 7849 46665 7883 46699
rect 2237 46529 2271 46563
rect 3249 46529 3283 46563
rect 6561 46529 6595 46563
rect 6745 46529 6779 46563
rect 8033 46529 8067 46563
rect 9873 46529 9907 46563
rect 1961 46461 1995 46495
rect 6377 46461 6411 46495
rect 10057 46393 10091 46427
rect 3433 46325 3467 46359
rect 2421 46121 2455 46155
rect 2053 45917 2087 45951
rect 2237 45917 2271 45951
rect 2881 45917 2915 45951
rect 9873 45917 9907 45951
rect 3065 45781 3099 45815
rect 10057 45781 10091 45815
rect 2329 45577 2363 45611
rect 1409 45441 1443 45475
rect 2145 45441 2179 45475
rect 2881 45441 2915 45475
rect 6561 45441 6595 45475
rect 3065 45305 3099 45339
rect 6377 45305 6411 45339
rect 1593 45237 1627 45271
rect 5365 45033 5399 45067
rect 6653 45033 6687 45067
rect 1777 44897 1811 44931
rect 1501 44829 1535 44863
rect 2789 44829 2823 44863
rect 5089 44829 5123 44863
rect 5181 44829 5215 44863
rect 5825 44829 5859 44863
rect 6009 44829 6043 44863
rect 6193 44829 6227 44863
rect 6837 44829 6871 44863
rect 9873 44829 9907 44863
rect 2973 44693 3007 44727
rect 10057 44693 10091 44727
rect 6377 44489 6411 44523
rect 1685 44353 1719 44387
rect 2973 44353 3007 44387
rect 6561 44353 6595 44387
rect 9873 44353 9907 44387
rect 1961 44285 1995 44319
rect 3157 44149 3191 44183
rect 10057 44149 10091 44183
rect 1869 43945 1903 43979
rect 2697 43945 2731 43979
rect 4905 43945 4939 43979
rect 1501 43809 1535 43843
rect 4537 43809 4571 43843
rect 1685 43741 1719 43775
rect 2329 43741 2363 43775
rect 2513 43741 2547 43775
rect 3801 43741 3835 43775
rect 4721 43741 4755 43775
rect 9873 43741 9907 43775
rect 3985 43605 4019 43639
rect 10057 43605 10091 43639
rect 3341 43401 3375 43435
rect 9965 43401 9999 43435
rect 3065 43333 3099 43367
rect 2789 43265 2823 43299
rect 2973 43265 3007 43299
rect 3157 43265 3191 43299
rect 3801 43265 3835 43299
rect 10149 43265 10183 43299
rect 1501 43197 1535 43231
rect 1777 43197 1811 43231
rect 3985 43129 4019 43163
rect 2145 42857 2179 42891
rect 1777 42721 1811 42755
rect 1961 42653 1995 42687
rect 2605 42653 2639 42687
rect 3801 42653 3835 42687
rect 6469 42653 6503 42687
rect 9873 42653 9907 42687
rect 2789 42517 2823 42551
rect 3985 42517 4019 42551
rect 6285 42517 6319 42551
rect 10057 42517 10091 42551
rect 1409 42177 1443 42211
rect 2145 42177 2179 42211
rect 2881 42177 2915 42211
rect 9873 42177 9907 42211
rect 1593 41973 1627 42007
rect 2329 41973 2363 42007
rect 3065 41973 3099 42007
rect 10057 41973 10091 42007
rect 2651 41769 2685 41803
rect 5089 41769 5123 41803
rect 9965 41769 9999 41803
rect 1961 41701 1995 41735
rect 2421 41633 2455 41667
rect 4721 41565 4755 41599
rect 4905 41565 4939 41599
rect 10149 41565 10183 41599
rect 1777 41497 1811 41531
rect 1961 41225 1995 41259
rect 2881 41225 2915 41259
rect 5365 41225 5399 41259
rect 1777 41089 1811 41123
rect 2697 41089 2731 41123
rect 3341 41089 3375 41123
rect 5181 41089 5215 41123
rect 9873 41089 9907 41123
rect 1593 41021 1627 41055
rect 2513 41021 2547 41055
rect 4997 41021 5031 41055
rect 3525 40953 3559 40987
rect 10057 40953 10091 40987
rect 9229 40681 9263 40715
rect 2421 40545 2455 40579
rect 1409 40477 1443 40511
rect 2145 40477 2179 40511
rect 3801 40477 3835 40511
rect 9413 40477 9447 40511
rect 9873 40477 9907 40511
rect 1593 40341 1627 40375
rect 3985 40341 4019 40375
rect 10057 40341 10091 40375
rect 2421 40137 2455 40171
rect 9229 40137 9263 40171
rect 3157 40069 3191 40103
rect 2237 40001 2271 40035
rect 2881 40001 2915 40035
rect 3801 40001 3835 40035
rect 9413 40001 9447 40035
rect 9873 40001 9907 40035
rect 2053 39933 2087 39967
rect 3985 39797 4019 39831
rect 10057 39797 10091 39831
rect 5641 39593 5675 39627
rect 9873 39593 9907 39627
rect 3157 39525 3191 39559
rect 6653 39525 6687 39559
rect 1409 39389 1443 39423
rect 2881 39389 2915 39423
rect 2973 39389 3007 39423
rect 3801 39389 3835 39423
rect 5273 39389 5307 39423
rect 5457 39389 5491 39423
rect 6837 39389 6871 39423
rect 10057 39389 10091 39423
rect 1593 39253 1627 39287
rect 3985 39253 4019 39287
rect 6745 39049 6779 39083
rect 1777 38913 1811 38947
rect 2789 38913 2823 38947
rect 3525 38913 3559 38947
rect 6561 38913 6595 38947
rect 9873 38913 9907 38947
rect 1501 38845 1535 38879
rect 6377 38845 6411 38879
rect 2973 38709 3007 38743
rect 3709 38709 3743 38743
rect 10057 38709 10091 38743
rect 2973 38505 3007 38539
rect 5273 38505 5307 38539
rect 1777 38369 1811 38403
rect 1501 38301 1535 38335
rect 4997 38301 5031 38335
rect 5089 38301 5123 38335
rect 9873 38301 9907 38335
rect 2881 38233 2915 38267
rect 10057 38165 10091 38199
rect 1869 37961 1903 37995
rect 2697 37961 2731 37995
rect 5089 37961 5123 37995
rect 3433 37893 3467 37927
rect 1501 37825 1535 37859
rect 1685 37825 1719 37859
rect 2329 37825 2363 37859
rect 2513 37825 2547 37859
rect 3249 37825 3283 37859
rect 4905 37825 4939 37859
rect 4721 37757 4755 37791
rect 2329 37281 2363 37315
rect 2513 37213 2547 37247
rect 2697 37213 2731 37247
rect 3801 37213 3835 37247
rect 8401 37213 8435 37247
rect 9873 37213 9907 37247
rect 1685 37145 1719 37179
rect 1777 37077 1811 37111
rect 3985 37077 4019 37111
rect 8217 37077 8251 37111
rect 10057 37077 10091 37111
rect 2421 36873 2455 36907
rect 3065 36873 3099 36907
rect 6377 36873 6411 36907
rect 7021 36873 7055 36907
rect 2237 36737 2271 36771
rect 2881 36737 2915 36771
rect 6561 36737 6595 36771
rect 7205 36737 7239 36771
rect 9873 36737 9907 36771
rect 2053 36669 2087 36703
rect 10057 36533 10091 36567
rect 1961 36329 1995 36363
rect 3985 36329 4019 36363
rect 4537 36329 4571 36363
rect 2513 36125 2547 36159
rect 3801 36125 3835 36159
rect 4721 36125 4755 36159
rect 9873 36125 9907 36159
rect 1869 36057 1903 36091
rect 2697 35989 2731 36023
rect 10057 35989 10091 36023
rect 2973 35785 3007 35819
rect 5457 35785 5491 35819
rect 6745 35785 6779 35819
rect 1409 35649 1443 35683
rect 2789 35649 2823 35683
rect 3985 35649 4019 35683
rect 4353 35649 4387 35683
rect 5273 35649 5307 35683
rect 6561 35649 6595 35683
rect 2605 35581 2639 35615
rect 5089 35581 5123 35615
rect 6377 35581 6411 35615
rect 1593 35445 1627 35479
rect 3801 35241 3835 35275
rect 1409 35037 1443 35071
rect 2145 35037 2179 35071
rect 3985 35037 4019 35071
rect 9873 35037 9907 35071
rect 1593 34901 1627 34935
rect 2329 34901 2363 34935
rect 10057 34901 10091 34935
rect 1593 34697 1627 34731
rect 3801 34697 3835 34731
rect 10057 34697 10091 34731
rect 1409 34561 1443 34595
rect 2145 34561 2179 34595
rect 2881 34561 2915 34595
rect 3985 34561 4019 34595
rect 9873 34561 9907 34595
rect 2329 34357 2363 34391
rect 3065 34357 3099 34391
rect 1961 34153 1995 34187
rect 5365 34153 5399 34187
rect 2789 34085 2823 34119
rect 4997 33949 5031 33983
rect 5181 33949 5215 33983
rect 1869 33881 1903 33915
rect 2605 33881 2639 33915
rect 2145 33609 2179 33643
rect 2973 33609 3007 33643
rect 3801 33609 3835 33643
rect 4261 33609 4295 33643
rect 5733 33609 5767 33643
rect 1869 33473 1903 33507
rect 1961 33473 1995 33507
rect 2789 33473 2823 33507
rect 3617 33473 3651 33507
rect 4445 33473 4479 33507
rect 5457 33473 5491 33507
rect 5549 33473 5583 33507
rect 9873 33473 9907 33507
rect 2605 33405 2639 33439
rect 3433 33405 3467 33439
rect 10057 33337 10091 33371
rect 2237 33065 2271 33099
rect 3157 33065 3191 33099
rect 4721 32997 4755 33031
rect 2789 32861 2823 32895
rect 2973 32861 3007 32895
rect 3801 32861 3835 32895
rect 4353 32861 4387 32895
rect 4537 32861 4571 32895
rect 9873 32861 9907 32895
rect 2145 32793 2179 32827
rect 3985 32725 4019 32759
rect 10057 32725 10091 32759
rect 2605 32521 2639 32555
rect 3249 32521 3283 32555
rect 1593 32385 1627 32419
rect 2421 32385 2455 32419
rect 3157 32385 3191 32419
rect 3801 32385 3835 32419
rect 2237 32317 2271 32351
rect 1777 32249 1811 32283
rect 3985 32181 4019 32215
rect 1777 31977 1811 32011
rect 2973 31977 3007 32011
rect 10057 31909 10091 31943
rect 1409 31841 1443 31875
rect 1593 31773 1627 31807
rect 2605 31773 2639 31807
rect 2789 31773 2823 31807
rect 3801 31773 3835 31807
rect 9873 31773 9907 31807
rect 3985 31637 4019 31671
rect 2237 31365 2271 31399
rect 2053 31297 2087 31331
rect 2697 31297 2731 31331
rect 3433 31297 3467 31331
rect 9873 31297 9907 31331
rect 3617 31161 3651 31195
rect 2881 31093 2915 31127
rect 10057 31093 10091 31127
rect 2513 30889 2547 30923
rect 2145 30753 2179 30787
rect 2329 30685 2363 30719
rect 9873 30685 9907 30719
rect 1501 30617 1535 30651
rect 1685 30617 1719 30651
rect 10057 30549 10091 30583
rect 1869 30209 1903 30243
rect 2513 30209 2547 30243
rect 2053 30141 2087 30175
rect 2697 30073 2731 30107
rect 2881 29801 2915 29835
rect 2053 29733 2087 29767
rect 3065 29597 3099 29631
rect 10149 29597 10183 29631
rect 1869 29529 1903 29563
rect 1961 29257 1995 29291
rect 2789 29189 2823 29223
rect 1869 29121 1903 29155
rect 2605 29121 2639 29155
rect 3341 29121 3375 29155
rect 3525 29053 3559 29087
rect 10149 28985 10183 29019
rect 3801 28713 3835 28747
rect 2421 28509 2455 28543
rect 2605 28509 2639 28543
rect 2789 28509 2823 28543
rect 3985 28509 4019 28543
rect 1777 28441 1811 28475
rect 1961 28441 1995 28475
rect 2145 28169 2179 28203
rect 2881 28101 2915 28135
rect 1961 28033 1995 28067
rect 2697 28033 2731 28067
rect 1777 27965 1811 27999
rect 9965 27965 9999 27999
rect 2973 27557 3007 27591
rect 1685 27489 1719 27523
rect 1409 27421 1443 27455
rect 2789 27353 2823 27387
rect 9965 27285 9999 27319
rect 3249 27013 3283 27047
rect 1501 26945 1535 26979
rect 2329 26945 2363 26979
rect 2513 26945 2547 26979
rect 3065 26945 3099 26979
rect 2145 26877 2179 26911
rect 1685 26809 1719 26843
rect 10149 26741 10183 26775
rect 2053 26537 2087 26571
rect 2789 26469 2823 26503
rect 1685 26333 1719 26367
rect 1869 26333 1903 26367
rect 2605 26265 2639 26299
rect 1961 25993 1995 26027
rect 3433 25993 3467 26027
rect 2789 25925 2823 25959
rect 1869 25857 1903 25891
rect 2605 25857 2639 25891
rect 3341 25857 3375 25891
rect 10149 25653 10183 25687
rect 1961 25449 1995 25483
rect 3985 25449 4019 25483
rect 2789 25381 2823 25415
rect 10149 25245 10183 25279
rect 1869 25177 1903 25211
rect 2605 25177 2639 25211
rect 3893 25177 3927 25211
rect 1777 24769 1811 24803
rect 2605 24769 2639 24803
rect 1961 24701 1995 24735
rect 2421 24701 2455 24735
rect 2789 24565 2823 24599
rect 2053 24293 2087 24327
rect 3801 24225 3835 24259
rect 4077 24225 4111 24259
rect 2697 24157 2731 24191
rect 2789 24157 2823 24191
rect 10149 24157 10183 24191
rect 1869 24089 1903 24123
rect 2973 24021 3007 24055
rect 3065 23817 3099 23851
rect 5089 23817 5123 23851
rect 1685 23681 1719 23715
rect 2881 23681 2915 23715
rect 3801 23681 3835 23715
rect 5273 23681 5307 23715
rect 1409 23613 1443 23647
rect 2697 23613 2731 23647
rect 4077 23613 4111 23647
rect 10149 23477 10183 23511
rect 4353 23273 4387 23307
rect 5089 23273 5123 23307
rect 1685 23137 1719 23171
rect 1409 23069 1443 23103
rect 2697 23069 2731 23103
rect 2881 23069 2915 23103
rect 4997 23069 5031 23103
rect 3065 23001 3099 23035
rect 4261 23001 4295 23035
rect 3617 22729 3651 22763
rect 2973 22661 3007 22695
rect 1869 22593 1903 22627
rect 2789 22593 2823 22627
rect 3525 22593 3559 22627
rect 1685 22525 1719 22559
rect 2605 22525 2639 22559
rect 2053 22457 2087 22491
rect 10149 22457 10183 22491
rect 10149 22117 10183 22151
rect 1685 22049 1719 22083
rect 2973 22049 3007 22083
rect 1409 21981 1443 22015
rect 2789 21981 2823 22015
rect 2881 21641 2915 21675
rect 3709 21573 3743 21607
rect 2789 21505 2823 21539
rect 3525 21505 3559 21539
rect 1409 21437 1443 21471
rect 1685 21437 1719 21471
rect 10149 21301 10183 21335
rect 3065 21097 3099 21131
rect 1409 20961 1443 20995
rect 1685 20961 1719 20995
rect 2697 20893 2731 20927
rect 2881 20893 2915 20927
rect 1685 20417 1719 20451
rect 2697 20417 2731 20451
rect 2973 20417 3007 20451
rect 9873 20417 9907 20451
rect 1409 20349 1443 20383
rect 10057 20281 10091 20315
rect 3065 20009 3099 20043
rect 1685 19873 1719 19907
rect 2697 19873 2731 19907
rect 1409 19805 1443 19839
rect 2881 19805 2915 19839
rect 9873 19805 9907 19839
rect 10057 19669 10091 19703
rect 9229 19465 9263 19499
rect 1685 19329 1719 19363
rect 2789 19329 2823 19363
rect 9413 19329 9447 19363
rect 10057 19329 10091 19363
rect 1409 19261 1443 19295
rect 2973 19193 3007 19227
rect 9873 19125 9907 19159
rect 3801 18921 3835 18955
rect 1409 18785 1443 18819
rect 1685 18785 1719 18819
rect 2973 18785 3007 18819
rect 2697 18717 2731 18751
rect 3985 18717 4019 18751
rect 9873 18717 9907 18751
rect 10057 18581 10091 18615
rect 2053 18377 2087 18411
rect 3525 18377 3559 18411
rect 2881 18309 2915 18343
rect 1777 18241 1811 18275
rect 1869 18241 1903 18275
rect 3709 18241 3743 18275
rect 9873 18241 9907 18275
rect 2513 18105 2547 18139
rect 2881 18037 2915 18071
rect 3065 18037 3099 18071
rect 10057 18037 10091 18071
rect 1409 17833 1443 17867
rect 3985 17833 4019 17867
rect 2421 17765 2455 17799
rect 4169 17765 4203 17799
rect 1593 17629 1627 17663
rect 2329 17629 2363 17663
rect 2881 17629 2915 17663
rect 3157 17629 3191 17663
rect 9873 17629 9907 17663
rect 3801 17561 3835 17595
rect 4001 17493 4035 17527
rect 10057 17493 10091 17527
rect 1961 17289 1995 17323
rect 9965 17289 9999 17323
rect 1869 17221 1903 17255
rect 2973 17153 3007 17187
rect 10149 17153 10183 17187
rect 3249 17085 3283 17119
rect 1593 16541 1627 16575
rect 2421 16541 2455 16575
rect 3065 16541 3099 16575
rect 3985 16541 4019 16575
rect 9873 16541 9907 16575
rect 1409 16405 1443 16439
rect 2237 16405 2271 16439
rect 2881 16405 2915 16439
rect 3801 16405 3835 16439
rect 10057 16405 10091 16439
rect 9229 16201 9263 16235
rect 1593 16065 1627 16099
rect 2237 16065 2271 16099
rect 2881 16065 2915 16099
rect 9413 16065 9447 16099
rect 9873 16065 9907 16099
rect 1409 15861 1443 15895
rect 2053 15861 2087 15895
rect 2697 15861 2731 15895
rect 10057 15861 10091 15895
rect 1961 15657 1995 15691
rect 9965 15657 9999 15691
rect 2881 15589 2915 15623
rect 1501 15521 1535 15555
rect 1593 15453 1627 15487
rect 1961 15453 1995 15487
rect 10149 15453 10183 15487
rect 2697 15385 2731 15419
rect 2145 15317 2179 15351
rect 2053 15113 2087 15147
rect 1961 15045 1995 15079
rect 2789 14977 2823 15011
rect 9873 14977 9907 15011
rect 10057 14841 10091 14875
rect 2605 14773 2639 14807
rect 1685 14569 1719 14603
rect 1869 14569 1903 14603
rect 2329 14569 2363 14603
rect 2697 14569 2731 14603
rect 1501 14433 1535 14467
rect 2421 14433 2455 14467
rect 1685 14365 1719 14399
rect 2329 14365 2363 14399
rect 3985 14365 4019 14399
rect 9873 14365 9907 14399
rect 1409 14297 1443 14331
rect 3801 14229 3835 14263
rect 10057 14229 10091 14263
rect 2605 14025 2639 14059
rect 9229 14025 9263 14059
rect 10057 14025 10091 14059
rect 1593 13889 1627 13923
rect 2789 13889 2823 13923
rect 3433 13889 3467 13923
rect 9413 13889 9447 13923
rect 9873 13889 9907 13923
rect 3249 13753 3283 13787
rect 1409 13685 1443 13719
rect 3065 13481 3099 13515
rect 9321 13481 9355 13515
rect 9965 13481 9999 13515
rect 2513 13413 2547 13447
rect 1593 13277 1627 13311
rect 2789 13277 2823 13311
rect 2881 13277 2915 13311
rect 3985 13277 4019 13311
rect 9505 13277 9539 13311
rect 10149 13277 10183 13311
rect 1409 13141 1443 13175
rect 2697 13141 2731 13175
rect 3801 13141 3835 13175
rect 1869 12937 1903 12971
rect 2907 12937 2941 12971
rect 3525 12937 3559 12971
rect 1409 12869 1443 12903
rect 2697 12869 2731 12903
rect 1685 12801 1719 12835
rect 3709 12801 3743 12835
rect 9873 12801 9907 12835
rect 1593 12733 1627 12767
rect 3065 12665 3099 12699
rect 1685 12597 1719 12631
rect 2881 12597 2915 12631
rect 10057 12597 10091 12631
rect 1685 12257 1719 12291
rect 1409 12189 1443 12223
rect 2881 12189 2915 12223
rect 9873 12189 9907 12223
rect 2697 12053 2731 12087
rect 10057 12053 10091 12087
rect 3065 11849 3099 11883
rect 9965 11849 9999 11883
rect 1685 11713 1719 11747
rect 2881 11713 2915 11747
rect 3709 11713 3743 11747
rect 10149 11713 10183 11747
rect 1409 11645 1443 11679
rect 2697 11645 2731 11679
rect 3525 11577 3559 11611
rect 3065 11305 3099 11339
rect 10057 11237 10091 11271
rect 1685 11169 1719 11203
rect 1409 11101 1443 11135
rect 2789 11101 2823 11135
rect 2881 11101 2915 11135
rect 9873 11101 9907 11135
rect 3433 10761 3467 10795
rect 1685 10625 1719 10659
rect 2697 10625 2731 10659
rect 3617 10625 3651 10659
rect 9873 10625 9907 10659
rect 1409 10557 1443 10591
rect 2881 10489 2915 10523
rect 10057 10421 10091 10455
rect 3985 10217 4019 10251
rect 2881 10149 2915 10183
rect 1685 10081 1719 10115
rect 1409 10013 1443 10047
rect 2697 10013 2731 10047
rect 3801 10013 3835 10047
rect 1685 9537 1719 9571
rect 2697 9537 2731 9571
rect 3617 9537 3651 9571
rect 4261 9537 4295 9571
rect 9873 9537 9907 9571
rect 1409 9469 1443 9503
rect 3433 9401 3467 9435
rect 4077 9401 4111 9435
rect 10057 9401 10091 9435
rect 2881 9333 2915 9367
rect 1685 8993 1719 9027
rect 1409 8925 1443 8959
rect 3249 8925 3283 8959
rect 3985 8925 4019 8959
rect 9873 8925 9907 8959
rect 3065 8789 3099 8823
rect 3801 8789 3835 8823
rect 10057 8789 10091 8823
rect 2881 8585 2915 8619
rect 1685 8449 1719 8483
rect 2697 8449 2731 8483
rect 9873 8449 9907 8483
rect 1409 8381 1443 8415
rect 10057 8313 10091 8347
rect 2881 8041 2915 8075
rect 1685 7905 1719 7939
rect 1409 7837 1443 7871
rect 2697 7837 2731 7871
rect 3985 7837 4019 7871
rect 3801 7701 3835 7735
rect 2973 7497 3007 7531
rect 3709 7497 3743 7531
rect 2053 7361 2087 7395
rect 2145 7361 2179 7395
rect 2881 7361 2915 7395
rect 3617 7361 3651 7395
rect 4445 7361 4479 7395
rect 9873 7361 9907 7395
rect 2329 7157 2363 7191
rect 4261 7157 4295 7191
rect 10057 7157 10091 7191
rect 2973 6817 3007 6851
rect 4445 6817 4479 6851
rect 1777 6749 1811 6783
rect 1961 6749 1995 6783
rect 2605 6749 2639 6783
rect 2789 6749 2823 6783
rect 9873 6749 9907 6783
rect 4261 6681 4295 6715
rect 2145 6613 2179 6647
rect 10057 6613 10091 6647
rect 1869 6409 1903 6443
rect 2605 6409 2639 6443
rect 1685 6273 1719 6307
rect 2421 6273 2455 6307
rect 3341 6273 3375 6307
rect 3525 6273 3559 6307
rect 3709 6069 3743 6103
rect 2881 5865 2915 5899
rect 4445 5865 4479 5899
rect 3801 5797 3835 5831
rect 1685 5729 1719 5763
rect 1409 5661 1443 5695
rect 2697 5661 2731 5695
rect 3985 5661 4019 5695
rect 4629 5661 4663 5695
rect 9873 5661 9907 5695
rect 10057 5525 10091 5559
rect 2881 5321 2915 5355
rect 3433 5321 3467 5355
rect 1409 5185 1443 5219
rect 2697 5185 2731 5219
rect 3617 5185 3651 5219
rect 4537 5185 4571 5219
rect 9413 5185 9447 5219
rect 9873 5185 9907 5219
rect 1685 5117 1719 5151
rect 9229 5049 9263 5083
rect 4353 4981 4387 5015
rect 10057 4981 10091 5015
rect 1961 4777 1995 4811
rect 2789 4777 2823 4811
rect 3801 4641 3835 4675
rect 1685 4573 1719 4607
rect 1777 4573 1811 4607
rect 2513 4573 2547 4607
rect 2605 4573 2639 4607
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 9873 4573 9907 4607
rect 4169 4505 4203 4539
rect 4629 4437 4663 4471
rect 10057 4437 10091 4471
rect 4629 4233 4663 4267
rect 1409 4097 1443 4131
rect 2789 4097 2823 4131
rect 2973 4097 3007 4131
rect 3617 4097 3651 4131
rect 4445 4097 4479 4131
rect 5273 4097 5307 4131
rect 2605 4029 2639 4063
rect 3433 4029 3467 4063
rect 4261 4029 4295 4063
rect 1593 3961 1627 3995
rect 3801 3893 3835 3927
rect 5089 3893 5123 3927
rect 1409 3689 1443 3723
rect 3801 3621 3835 3655
rect 1593 3485 1627 3519
rect 2513 3485 2547 3519
rect 3985 3485 4019 3519
rect 4629 3485 4663 3519
rect 9873 3485 9907 3519
rect 2329 3349 2363 3383
rect 4445 3349 4479 3383
rect 10057 3349 10091 3383
rect 1409 3145 1443 3179
rect 2053 3145 2087 3179
rect 2697 3145 2731 3179
rect 3341 3145 3375 3179
rect 1593 3009 1627 3043
rect 2237 3009 2271 3043
rect 2881 3009 2915 3043
rect 3525 3009 3559 3043
rect 9137 3009 9171 3043
rect 9873 3009 9907 3043
rect 9321 2805 9355 2839
rect 10057 2805 10091 2839
rect 2053 2601 2087 2635
rect 3801 2601 3835 2635
rect 1409 2533 1443 2567
rect 2697 2533 2731 2567
rect 1593 2397 1627 2431
rect 2237 2397 2271 2431
rect 2881 2397 2915 2431
rect 3985 2397 4019 2431
rect 4629 2397 4663 2431
rect 9137 2397 9171 2431
rect 9873 2397 9907 2431
rect 4445 2261 4479 2295
rect 9321 2261 9355 2295
rect 10057 2261 10091 2295
<< metal1 >>
rect 1104 77818 10856 77840
rect 1104 77766 2582 77818
rect 2634 77766 2646 77818
rect 2698 77766 2710 77818
rect 2762 77766 2774 77818
rect 2826 77766 2838 77818
rect 2890 77766 5846 77818
rect 5898 77766 5910 77818
rect 5962 77766 5974 77818
rect 6026 77766 6038 77818
rect 6090 77766 6102 77818
rect 6154 77766 9110 77818
rect 9162 77766 9174 77818
rect 9226 77766 9238 77818
rect 9290 77766 9302 77818
rect 9354 77766 9366 77818
rect 9418 77766 10856 77818
rect 1104 77744 10856 77766
rect 1394 77568 1400 77580
rect 1355 77540 1400 77568
rect 1394 77528 1400 77540
rect 1452 77528 1458 77580
rect 3786 77528 3792 77580
rect 3844 77568 3850 77580
rect 10137 77571 10195 77577
rect 10137 77568 10149 77571
rect 3844 77540 10149 77568
rect 3844 77528 3850 77540
rect 10137 77537 10149 77540
rect 10183 77537 10195 77571
rect 10137 77531 10195 77537
rect 1673 77503 1731 77509
rect 1673 77469 1685 77503
rect 1719 77500 1731 77503
rect 1762 77500 1768 77512
rect 1719 77472 1768 77500
rect 1719 77469 1731 77472
rect 1673 77463 1731 77469
rect 1762 77460 1768 77472
rect 1820 77460 1826 77512
rect 2866 77500 2872 77512
rect 2827 77472 2872 77500
rect 2866 77460 2872 77472
rect 2924 77460 2930 77512
rect 3970 77500 3976 77512
rect 3931 77472 3976 77500
rect 3970 77460 3976 77472
rect 4028 77460 4034 77512
rect 4062 77460 4068 77512
rect 4120 77500 4126 77512
rect 4617 77503 4675 77509
rect 4617 77500 4629 77503
rect 4120 77472 4629 77500
rect 4120 77460 4126 77472
rect 4617 77469 4629 77472
rect 4663 77469 4675 77503
rect 9398 77500 9404 77512
rect 9359 77472 9404 77500
rect 4617 77463 4675 77469
rect 9398 77460 9404 77472
rect 9456 77460 9462 77512
rect 9950 77500 9956 77512
rect 9911 77472 9956 77500
rect 9950 77460 9956 77472
rect 10008 77460 10014 77512
rect 2222 77324 2228 77376
rect 2280 77364 2286 77376
rect 2685 77367 2743 77373
rect 2685 77364 2697 77367
rect 2280 77336 2697 77364
rect 2280 77324 2286 77336
rect 2685 77333 2697 77336
rect 2731 77333 2743 77367
rect 2685 77327 2743 77333
rect 3050 77324 3056 77376
rect 3108 77364 3114 77376
rect 3789 77367 3847 77373
rect 3789 77364 3801 77367
rect 3108 77336 3801 77364
rect 3108 77324 3114 77336
rect 3789 77333 3801 77336
rect 3835 77333 3847 77367
rect 3789 77327 3847 77333
rect 4062 77324 4068 77376
rect 4120 77364 4126 77376
rect 4433 77367 4491 77373
rect 4433 77364 4445 77367
rect 4120 77336 4445 77364
rect 4120 77324 4126 77336
rect 4433 77333 4445 77336
rect 4479 77333 4491 77367
rect 4433 77327 4491 77333
rect 8294 77324 8300 77376
rect 8352 77364 8358 77376
rect 9217 77367 9275 77373
rect 9217 77364 9229 77367
rect 8352 77336 9229 77364
rect 8352 77324 8358 77336
rect 9217 77333 9229 77336
rect 9263 77333 9275 77367
rect 9217 77327 9275 77333
rect 1104 77274 10856 77296
rect 1104 77222 4214 77274
rect 4266 77222 4278 77274
rect 4330 77222 4342 77274
rect 4394 77222 4406 77274
rect 4458 77222 4470 77274
rect 4522 77222 7478 77274
rect 7530 77222 7542 77274
rect 7594 77222 7606 77274
rect 7658 77222 7670 77274
rect 7722 77222 7734 77274
rect 7786 77222 10856 77274
rect 1104 77200 10856 77222
rect 1302 76984 1308 77036
rect 1360 77024 1366 77036
rect 1397 77027 1455 77033
rect 1397 77024 1409 77027
rect 1360 76996 1409 77024
rect 1360 76984 1366 76996
rect 1397 76993 1409 76996
rect 1443 76993 1455 77027
rect 1397 76987 1455 76993
rect 1486 76984 1492 77036
rect 1544 77024 1550 77036
rect 2317 77027 2375 77033
rect 2317 77024 2329 77027
rect 1544 76996 2329 77024
rect 1544 76984 1550 76996
rect 2317 76993 2329 76996
rect 2363 76993 2375 77027
rect 2958 77024 2964 77036
rect 2919 76996 2964 77024
rect 2317 76987 2375 76993
rect 2958 76984 2964 76996
rect 3016 76984 3022 77036
rect 3602 77024 3608 77036
rect 3563 76996 3608 77024
rect 3602 76984 3608 76996
rect 3660 76984 3666 77036
rect 3878 76984 3884 77036
rect 3936 77024 3942 77036
rect 4249 77027 4307 77033
rect 4249 77024 4261 77027
rect 3936 76996 4261 77024
rect 3936 76984 3942 76996
rect 4249 76993 4261 76996
rect 4295 76993 4307 77027
rect 4249 76987 4307 76993
rect 9401 77027 9459 77033
rect 9401 76993 9413 77027
rect 9447 77024 9459 77027
rect 9490 77024 9496 77036
rect 9447 76996 9496 77024
rect 9447 76993 9459 76996
rect 9401 76987 9459 76993
rect 9490 76984 9496 76996
rect 9548 76984 9554 77036
rect 9582 76984 9588 77036
rect 9640 77024 9646 77036
rect 9861 77027 9919 77033
rect 9861 77024 9873 77027
rect 9640 76996 9873 77024
rect 9640 76984 9646 76996
rect 9861 76993 9873 76996
rect 9907 76993 9919 77027
rect 9861 76987 9919 76993
rect 2498 76848 2504 76900
rect 2556 76888 2562 76900
rect 9217 76891 9275 76897
rect 9217 76888 9229 76891
rect 2556 76860 9229 76888
rect 2556 76848 2562 76860
rect 9217 76857 9229 76860
rect 9263 76857 9275 76891
rect 9217 76851 9275 76857
rect 1394 76780 1400 76832
rect 1452 76820 1458 76832
rect 1581 76823 1639 76829
rect 1581 76820 1593 76823
rect 1452 76792 1593 76820
rect 1452 76780 1458 76792
rect 1581 76789 1593 76792
rect 1627 76789 1639 76823
rect 1581 76783 1639 76789
rect 2133 76823 2191 76829
rect 2133 76789 2145 76823
rect 2179 76820 2191 76823
rect 2314 76820 2320 76832
rect 2179 76792 2320 76820
rect 2179 76789 2191 76792
rect 2133 76783 2191 76789
rect 2314 76780 2320 76792
rect 2372 76780 2378 76832
rect 2777 76823 2835 76829
rect 2777 76789 2789 76823
rect 2823 76820 2835 76823
rect 3142 76820 3148 76832
rect 2823 76792 3148 76820
rect 2823 76789 2835 76792
rect 2777 76783 2835 76789
rect 3142 76780 3148 76792
rect 3200 76780 3206 76832
rect 3418 76820 3424 76832
rect 3379 76792 3424 76820
rect 3418 76780 3424 76792
rect 3476 76780 3482 76832
rect 4062 76820 4068 76832
rect 4023 76792 4068 76820
rect 4062 76780 4068 76792
rect 4120 76780 4126 76832
rect 9766 76780 9772 76832
rect 9824 76820 9830 76832
rect 10045 76823 10103 76829
rect 10045 76820 10057 76823
rect 9824 76792 10057 76820
rect 9824 76780 9830 76792
rect 10045 76789 10057 76792
rect 10091 76789 10103 76823
rect 10045 76783 10103 76789
rect 1104 76730 10856 76752
rect 1104 76678 2582 76730
rect 2634 76678 2646 76730
rect 2698 76678 2710 76730
rect 2762 76678 2774 76730
rect 2826 76678 2838 76730
rect 2890 76678 5846 76730
rect 5898 76678 5910 76730
rect 5962 76678 5974 76730
rect 6026 76678 6038 76730
rect 6090 76678 6102 76730
rect 6154 76678 9110 76730
rect 9162 76678 9174 76730
rect 9226 76678 9238 76730
rect 9290 76678 9302 76730
rect 9354 76678 9366 76730
rect 9418 76678 10856 76730
rect 1104 76656 10856 76678
rect 9953 76619 10011 76625
rect 9953 76616 9965 76619
rect 1504 76588 9965 76616
rect 1397 76415 1455 76421
rect 1397 76381 1409 76415
rect 1443 76412 1455 76415
rect 1504 76412 1532 76588
rect 9953 76585 9965 76588
rect 9999 76585 10011 76619
rect 9953 76579 10011 76585
rect 1946 76548 1952 76560
rect 1907 76520 1952 76548
rect 1946 76508 1952 76520
rect 2004 76508 2010 76560
rect 3053 76551 3111 76557
rect 3053 76517 3065 76551
rect 3099 76548 3111 76551
rect 3786 76548 3792 76560
rect 3099 76520 3792 76548
rect 3099 76517 3111 76520
rect 3053 76511 3111 76517
rect 3786 76508 3792 76520
rect 3844 76508 3850 76560
rect 2130 76480 2136 76492
rect 1596 76452 2136 76480
rect 1596 76421 1624 76452
rect 2130 76440 2136 76452
rect 2188 76440 2194 76492
rect 2424 76452 2917 76480
rect 1443 76384 1532 76412
rect 1581 76415 1639 76421
rect 1443 76381 1455 76384
rect 1397 76375 1455 76381
rect 1581 76381 1593 76415
rect 1627 76381 1639 76415
rect 1581 76375 1639 76381
rect 1817 76415 1875 76421
rect 1817 76381 1829 76415
rect 1863 76412 1875 76415
rect 2038 76412 2044 76424
rect 1863 76384 2044 76412
rect 1863 76381 1875 76384
rect 1817 76375 1875 76381
rect 2038 76372 2044 76384
rect 2096 76412 2102 76424
rect 2424 76412 2452 76452
rect 2096 76384 2452 76412
rect 2096 76372 2102 76384
rect 2498 76372 2504 76424
rect 2556 76412 2562 76424
rect 2889 76421 2917 76452
rect 2874 76415 2932 76421
rect 2556 76384 2601 76412
rect 2556 76372 2562 76384
rect 2874 76381 2886 76415
rect 2920 76381 2932 76415
rect 10134 76412 10140 76424
rect 10095 76384 10140 76412
rect 2874 76375 2932 76381
rect 10134 76372 10140 76384
rect 10192 76372 10198 76424
rect 1673 76347 1731 76353
rect 1673 76313 1685 76347
rect 1719 76313 1731 76347
rect 1673 76307 1731 76313
rect 1688 76276 1716 76307
rect 2130 76304 2136 76356
rect 2188 76344 2194 76356
rect 2685 76347 2743 76353
rect 2685 76344 2697 76347
rect 2188 76316 2697 76344
rect 2188 76304 2194 76316
rect 2685 76313 2697 76316
rect 2731 76313 2743 76347
rect 2685 76307 2743 76313
rect 2777 76347 2835 76353
rect 2777 76313 2789 76347
rect 2823 76344 2835 76347
rect 4062 76344 4068 76356
rect 2823 76316 4068 76344
rect 2823 76313 2835 76316
rect 2777 76307 2835 76313
rect 4062 76304 4068 76316
rect 4120 76304 4126 76356
rect 3418 76276 3424 76288
rect 1688 76248 3424 76276
rect 3418 76236 3424 76248
rect 3476 76236 3482 76288
rect 1104 76186 10856 76208
rect 1104 76134 4214 76186
rect 4266 76134 4278 76186
rect 4330 76134 4342 76186
rect 4394 76134 4406 76186
rect 4458 76134 4470 76186
rect 4522 76134 7478 76186
rect 7530 76134 7542 76186
rect 7594 76134 7606 76186
rect 7658 76134 7670 76186
rect 7722 76134 7734 76186
rect 7786 76134 10856 76186
rect 1104 76112 10856 76134
rect 1397 76075 1455 76081
rect 1397 76041 1409 76075
rect 1443 76072 1455 76075
rect 1670 76072 1676 76084
rect 1443 76044 1676 76072
rect 1443 76041 1455 76044
rect 1397 76035 1455 76041
rect 1670 76032 1676 76044
rect 1728 76032 1734 76084
rect 9953 76075 10011 76081
rect 9953 76072 9965 76075
rect 2332 76044 9965 76072
rect 1578 75936 1584 75948
rect 1539 75908 1584 75936
rect 1578 75896 1584 75908
rect 1636 75896 1642 75948
rect 2332 75945 2360 76044
rect 9953 76041 9965 76044
rect 9999 76041 10011 76075
rect 9953 76035 10011 76041
rect 2590 76004 2596 76016
rect 2551 75976 2596 76004
rect 2590 75964 2596 75976
rect 2648 75964 2654 76016
rect 2886 76007 2944 76013
rect 2886 75973 2898 76007
rect 2932 76004 2944 76007
rect 3510 76004 3516 76016
rect 2932 75976 3516 76004
rect 2932 75973 2944 75976
rect 2886 75967 2944 75973
rect 3510 75964 3516 75976
rect 3568 75964 3574 76016
rect 2317 75939 2375 75945
rect 2317 75905 2329 75939
rect 2363 75905 2375 75939
rect 2498 75936 2504 75948
rect 2459 75908 2504 75936
rect 2317 75899 2375 75905
rect 2498 75896 2504 75908
rect 2556 75896 2562 75948
rect 2690 75939 2748 75945
rect 2690 75905 2702 75939
rect 2736 75905 2748 75939
rect 3602 75936 3608 75948
rect 3563 75908 3608 75936
rect 2690 75899 2748 75905
rect 2038 75828 2044 75880
rect 2096 75868 2102 75880
rect 2700 75868 2728 75899
rect 3602 75896 3608 75908
rect 3660 75896 3666 75948
rect 10134 75936 10140 75948
rect 10095 75908 10140 75936
rect 10134 75896 10140 75908
rect 10192 75896 10198 75948
rect 2096 75840 2728 75868
rect 2096 75828 2102 75840
rect 2130 75760 2136 75812
rect 2188 75800 2194 75812
rect 2498 75800 2504 75812
rect 2188 75772 2504 75800
rect 2188 75760 2194 75772
rect 2498 75760 2504 75772
rect 2556 75760 2562 75812
rect 3418 75732 3424 75744
rect 3379 75704 3424 75732
rect 3418 75692 3424 75704
rect 3476 75692 3482 75744
rect 1104 75642 10856 75664
rect 1104 75590 2582 75642
rect 2634 75590 2646 75642
rect 2698 75590 2710 75642
rect 2762 75590 2774 75642
rect 2826 75590 2838 75642
rect 2890 75590 5846 75642
rect 5898 75590 5910 75642
rect 5962 75590 5974 75642
rect 6026 75590 6038 75642
rect 6090 75590 6102 75642
rect 6154 75590 9110 75642
rect 9162 75590 9174 75642
rect 9226 75590 9238 75642
rect 9290 75590 9302 75642
rect 9354 75590 9366 75642
rect 9418 75590 10856 75642
rect 1104 75568 10856 75590
rect 1854 75488 1860 75540
rect 1912 75528 1918 75540
rect 3053 75531 3111 75537
rect 3053 75528 3065 75531
rect 1912 75500 3065 75528
rect 1912 75488 1918 75500
rect 3053 75497 3065 75500
rect 3099 75497 3111 75531
rect 3053 75491 3111 75497
rect 2498 75460 2504 75472
rect 2459 75432 2504 75460
rect 2498 75420 2504 75432
rect 2556 75420 2562 75472
rect 9953 75463 10011 75469
rect 9953 75460 9965 75463
rect 2746 75432 9965 75460
rect 2746 75392 2774 75432
rect 9953 75429 9965 75432
rect 9999 75429 10011 75463
rect 9953 75423 10011 75429
rect 1964 75364 2774 75392
rect 1964 75333 1992 75364
rect 1949 75327 2007 75333
rect 1949 75293 1961 75327
rect 1995 75293 2007 75327
rect 2222 75324 2228 75336
rect 2183 75296 2228 75324
rect 1949 75287 2007 75293
rect 2222 75284 2228 75296
rect 2280 75284 2286 75336
rect 2345 75327 2403 75333
rect 2345 75324 2357 75327
rect 2332 75293 2357 75324
rect 2391 75293 2403 75327
rect 3234 75324 3240 75336
rect 3195 75296 3240 75324
rect 2332 75287 2403 75293
rect 2130 75256 2136 75268
rect 2091 75228 2136 75256
rect 2130 75216 2136 75228
rect 2188 75216 2194 75268
rect 2038 75148 2044 75200
rect 2096 75188 2102 75200
rect 2332 75188 2360 75287
rect 3234 75284 3240 75296
rect 3292 75284 3298 75336
rect 10134 75324 10140 75336
rect 10095 75296 10140 75324
rect 10134 75284 10140 75296
rect 10192 75284 10198 75336
rect 2096 75160 2360 75188
rect 2096 75148 2102 75160
rect 1104 75098 10856 75120
rect 1104 75046 4214 75098
rect 4266 75046 4278 75098
rect 4330 75046 4342 75098
rect 4394 75046 4406 75098
rect 4458 75046 4470 75098
rect 4522 75046 7478 75098
rect 7530 75046 7542 75098
rect 7594 75046 7606 75098
rect 7658 75046 7670 75098
rect 7722 75046 7734 75098
rect 7786 75046 10856 75098
rect 1104 75024 10856 75046
rect 2130 74984 2136 74996
rect 1596 74956 2136 74984
rect 1596 74925 1624 74956
rect 2130 74944 2136 74956
rect 2188 74944 2194 74996
rect 1581 74919 1639 74925
rect 1581 74885 1593 74919
rect 1627 74885 1639 74919
rect 1581 74879 1639 74885
rect 1673 74919 1731 74925
rect 1673 74885 1685 74919
rect 1719 74916 1731 74919
rect 3970 74916 3976 74928
rect 1719 74888 3976 74916
rect 1719 74885 1731 74888
rect 1673 74879 1731 74885
rect 3970 74876 3976 74888
rect 4028 74876 4034 74928
rect 1397 74851 1455 74857
rect 1397 74817 1409 74851
rect 1443 74817 1455 74851
rect 1397 74811 1455 74817
rect 1817 74851 1875 74857
rect 1817 74817 1829 74851
rect 1863 74848 1875 74851
rect 2038 74848 2044 74860
rect 1863 74820 2044 74848
rect 1863 74817 1875 74820
rect 1817 74811 1875 74817
rect 1412 74780 1440 74811
rect 2038 74808 2044 74820
rect 2096 74808 2102 74860
rect 2685 74851 2743 74857
rect 2685 74817 2697 74851
rect 2731 74848 2743 74851
rect 2958 74848 2964 74860
rect 2731 74820 2964 74848
rect 2731 74817 2743 74820
rect 2685 74811 2743 74817
rect 2958 74808 2964 74820
rect 3016 74808 3022 74860
rect 8294 74780 8300 74792
rect 1412 74752 8300 74780
rect 8294 74740 8300 74752
rect 8352 74740 8358 74792
rect 1486 74672 1492 74724
rect 1544 74712 1550 74724
rect 2501 74715 2559 74721
rect 2501 74712 2513 74715
rect 1544 74684 2513 74712
rect 1544 74672 1550 74684
rect 2501 74681 2513 74684
rect 2547 74681 2559 74715
rect 2501 74675 2559 74681
rect 1946 74644 1952 74656
rect 1907 74616 1952 74644
rect 1946 74604 1952 74616
rect 2004 74604 2010 74656
rect 1104 74554 10856 74576
rect 1104 74502 2582 74554
rect 2634 74502 2646 74554
rect 2698 74502 2710 74554
rect 2762 74502 2774 74554
rect 2826 74502 2838 74554
rect 2890 74502 5846 74554
rect 5898 74502 5910 74554
rect 5962 74502 5974 74554
rect 6026 74502 6038 74554
rect 6090 74502 6102 74554
rect 6154 74502 9110 74554
rect 9162 74502 9174 74554
rect 9226 74502 9238 74554
rect 9290 74502 9302 74554
rect 9354 74502 9366 74554
rect 9418 74502 10856 74554
rect 1104 74480 10856 74502
rect 2406 74332 2412 74384
rect 2464 74372 2470 74384
rect 2501 74375 2559 74381
rect 2501 74372 2513 74375
rect 2464 74344 2513 74372
rect 2464 74332 2470 74344
rect 2501 74341 2513 74344
rect 2547 74341 2559 74375
rect 9953 74375 10011 74381
rect 9953 74372 9965 74375
rect 2501 74335 2559 74341
rect 2746 74344 9965 74372
rect 2746 74304 2774 74344
rect 9953 74341 9965 74344
rect 9999 74341 10011 74375
rect 9953 74335 10011 74341
rect 1964 74276 2774 74304
rect 1964 74245 1992 74276
rect 1949 74239 2007 74245
rect 1949 74205 1961 74239
rect 1995 74205 2007 74239
rect 1949 74199 2007 74205
rect 2038 74196 2044 74248
rect 2096 74236 2102 74248
rect 2369 74239 2427 74245
rect 2369 74236 2381 74239
rect 2096 74208 2381 74236
rect 2096 74196 2102 74208
rect 2369 74205 2381 74208
rect 2415 74236 2427 74239
rect 2866 74236 2872 74248
rect 2415 74208 2872 74236
rect 2415 74205 2427 74208
rect 2369 74199 2427 74205
rect 2866 74196 2872 74208
rect 2924 74196 2930 74248
rect 3234 74236 3240 74248
rect 3195 74208 3240 74236
rect 3234 74196 3240 74208
rect 3292 74196 3298 74248
rect 10134 74236 10140 74248
rect 10095 74208 10140 74236
rect 10134 74196 10140 74208
rect 10192 74196 10198 74248
rect 2130 74168 2136 74180
rect 2091 74140 2136 74168
rect 2130 74128 2136 74140
rect 2188 74128 2194 74180
rect 2225 74171 2283 74177
rect 2225 74137 2237 74171
rect 2271 74168 2283 74171
rect 3142 74168 3148 74180
rect 2271 74140 3148 74168
rect 2271 74137 2283 74140
rect 2225 74131 2283 74137
rect 3142 74128 3148 74140
rect 3200 74128 3206 74180
rect 3053 74103 3111 74109
rect 3053 74069 3065 74103
rect 3099 74100 3111 74103
rect 3234 74100 3240 74112
rect 3099 74072 3240 74100
rect 3099 74069 3111 74072
rect 3053 74063 3111 74069
rect 3234 74060 3240 74072
rect 3292 74060 3298 74112
rect 1104 74010 10856 74032
rect 1104 73958 4214 74010
rect 4266 73958 4278 74010
rect 4330 73958 4342 74010
rect 4394 73958 4406 74010
rect 4458 73958 4470 74010
rect 4522 73958 7478 74010
rect 7530 73958 7542 74010
rect 7594 73958 7606 74010
rect 7658 73958 7670 74010
rect 7722 73958 7734 74010
rect 7786 73958 10856 74010
rect 1104 73936 10856 73958
rect 1578 73760 1584 73772
rect 1539 73732 1584 73760
rect 1578 73720 1584 73732
rect 1636 73720 1642 73772
rect 2222 73760 2228 73772
rect 2183 73732 2228 73760
rect 2222 73720 2228 73732
rect 2280 73720 2286 73772
rect 10134 73760 10140 73772
rect 10095 73732 10140 73760
rect 10134 73720 10140 73732
rect 10192 73720 10198 73772
rect 1210 73652 1216 73704
rect 1268 73692 1274 73704
rect 1268 73664 9674 73692
rect 1268 73652 1274 73664
rect 1397 73627 1455 73633
rect 1397 73593 1409 73627
rect 1443 73624 1455 73627
rect 3142 73624 3148 73636
rect 1443 73596 3148 73624
rect 1443 73593 1455 73596
rect 1397 73587 1455 73593
rect 3142 73584 3148 73596
rect 3200 73584 3206 73636
rect 2038 73556 2044 73568
rect 1999 73528 2044 73556
rect 2038 73516 2044 73528
rect 2096 73516 2102 73568
rect 9646 73556 9674 73664
rect 9953 73559 10011 73565
rect 9953 73556 9965 73559
rect 9646 73528 9965 73556
rect 9953 73525 9965 73528
rect 9999 73525 10011 73559
rect 9953 73519 10011 73525
rect 1104 73466 10856 73488
rect 1104 73414 2582 73466
rect 2634 73414 2646 73466
rect 2698 73414 2710 73466
rect 2762 73414 2774 73466
rect 2826 73414 2838 73466
rect 2890 73414 5846 73466
rect 5898 73414 5910 73466
rect 5962 73414 5974 73466
rect 6026 73414 6038 73466
rect 6090 73414 6102 73466
rect 6154 73414 9110 73466
rect 9162 73414 9174 73466
rect 9226 73414 9238 73466
rect 9290 73414 9302 73466
rect 9354 73414 9366 73466
rect 9418 73414 10856 73466
rect 1104 73392 10856 73414
rect 1504 73256 9674 73284
rect 1397 73151 1455 73157
rect 1397 73117 1409 73151
rect 1443 73148 1455 73151
rect 1504 73148 1532 73256
rect 2130 73216 2136 73228
rect 1596 73188 2136 73216
rect 1596 73157 1624 73188
rect 2130 73176 2136 73188
rect 2188 73176 2194 73228
rect 1443 73120 1532 73148
rect 1581 73151 1639 73157
rect 1443 73117 1455 73120
rect 1397 73111 1455 73117
rect 1581 73117 1593 73151
rect 1627 73117 1639 73151
rect 1581 73111 1639 73117
rect 1817 73151 1875 73157
rect 1817 73117 1829 73151
rect 1863 73148 1875 73151
rect 2958 73148 2964 73160
rect 1863 73120 2964 73148
rect 1863 73117 1875 73120
rect 1817 73111 1875 73117
rect 2958 73108 2964 73120
rect 3016 73108 3022 73160
rect 9646 73148 9674 73256
rect 9950 73148 9956 73160
rect 9646 73120 9956 73148
rect 9950 73108 9956 73120
rect 10008 73108 10014 73160
rect 1673 73083 1731 73089
rect 1673 73049 1685 73083
rect 1719 73049 1731 73083
rect 1673 73043 1731 73049
rect 1688 73012 1716 73043
rect 1854 73012 1860 73024
rect 1688 72984 1860 73012
rect 1854 72972 1860 72984
rect 1912 72972 1918 73024
rect 1966 73015 2024 73021
rect 1966 72981 1978 73015
rect 2012 73012 2024 73015
rect 4706 73012 4712 73024
rect 2012 72984 4712 73012
rect 2012 72981 2024 72984
rect 1966 72975 2024 72981
rect 4706 72972 4712 72984
rect 4764 72972 4770 73024
rect 1104 72922 10856 72944
rect 1104 72870 4214 72922
rect 4266 72870 4278 72922
rect 4330 72870 4342 72922
rect 4394 72870 4406 72922
rect 4458 72870 4470 72922
rect 4522 72870 7478 72922
rect 7530 72870 7542 72922
rect 7594 72870 7606 72922
rect 7658 72870 7670 72922
rect 7722 72870 7734 72922
rect 7786 72870 10856 72922
rect 1104 72848 10856 72870
rect 1394 72632 1400 72684
rect 1452 72672 1458 72684
rect 1581 72675 1639 72681
rect 1581 72672 1593 72675
rect 1452 72644 1593 72672
rect 1452 72632 1458 72644
rect 1581 72641 1593 72644
rect 1627 72641 1639 72675
rect 2222 72672 2228 72684
rect 2183 72644 2228 72672
rect 1581 72635 1639 72641
rect 2222 72632 2228 72644
rect 2280 72632 2286 72684
rect 2866 72672 2872 72684
rect 2827 72644 2872 72672
rect 2866 72632 2872 72644
rect 2924 72632 2930 72684
rect 10134 72672 10140 72684
rect 10095 72644 10140 72672
rect 10134 72632 10140 72644
rect 10192 72632 10198 72684
rect 2041 72539 2099 72545
rect 2041 72505 2053 72539
rect 2087 72536 2099 72539
rect 3326 72536 3332 72548
rect 2087 72508 3332 72536
rect 2087 72505 2099 72508
rect 2041 72499 2099 72505
rect 3326 72496 3332 72508
rect 3384 72496 3390 72548
rect 1397 72471 1455 72477
rect 1397 72437 1409 72471
rect 1443 72468 1455 72471
rect 1486 72468 1492 72480
rect 1443 72440 1492 72468
rect 1443 72437 1455 72440
rect 1397 72431 1455 72437
rect 1486 72428 1492 72440
rect 1544 72428 1550 72480
rect 2498 72428 2504 72480
rect 2556 72468 2562 72480
rect 2685 72471 2743 72477
rect 2685 72468 2697 72471
rect 2556 72440 2697 72468
rect 2556 72428 2562 72440
rect 2685 72437 2697 72440
rect 2731 72437 2743 72471
rect 2685 72431 2743 72437
rect 8294 72428 8300 72480
rect 8352 72468 8358 72480
rect 9953 72471 10011 72477
rect 9953 72468 9965 72471
rect 8352 72440 9965 72468
rect 8352 72428 8358 72440
rect 9953 72437 9965 72440
rect 9999 72437 10011 72471
rect 9953 72431 10011 72437
rect 1104 72378 10856 72400
rect 1104 72326 2582 72378
rect 2634 72326 2646 72378
rect 2698 72326 2710 72378
rect 2762 72326 2774 72378
rect 2826 72326 2838 72378
rect 2890 72326 5846 72378
rect 5898 72326 5910 72378
rect 5962 72326 5974 72378
rect 6026 72326 6038 72378
rect 6090 72326 6102 72378
rect 6154 72326 9110 72378
rect 9162 72326 9174 72378
rect 9226 72326 9238 72378
rect 9290 72326 9302 72378
rect 9354 72326 9366 72378
rect 9418 72326 10856 72378
rect 1104 72304 10856 72326
rect 9950 72264 9956 72276
rect 9911 72236 9956 72264
rect 9950 72224 9956 72236
rect 10008 72224 10014 72276
rect 658 72156 664 72208
rect 716 72196 722 72208
rect 2593 72199 2651 72205
rect 2593 72196 2605 72199
rect 716 72168 2605 72196
rect 716 72156 722 72168
rect 2593 72165 2605 72168
rect 2639 72165 2651 72199
rect 2593 72159 2651 72165
rect 1210 72088 1216 72140
rect 1268 72128 1274 72140
rect 1268 72100 2084 72128
rect 1268 72088 1274 72100
rect 1578 72060 1584 72072
rect 1539 72032 1584 72060
rect 1578 72020 1584 72032
rect 1636 72020 1642 72072
rect 2056 72069 2084 72100
rect 2130 72088 2136 72140
rect 2188 72128 2194 72140
rect 2188 72100 2268 72128
rect 2188 72088 2194 72100
rect 2240 72069 2268 72100
rect 2041 72063 2099 72069
rect 2041 72029 2053 72063
rect 2087 72029 2099 72063
rect 2041 72023 2099 72029
rect 2225 72063 2283 72069
rect 2225 72029 2237 72063
rect 2271 72029 2283 72063
rect 2225 72023 2283 72029
rect 2314 72020 2320 72072
rect 2372 72060 2378 72072
rect 2461 72063 2519 72069
rect 2372 72032 2417 72060
rect 2372 72020 2378 72032
rect 2461 72029 2473 72063
rect 2507 72060 2519 72063
rect 2866 72060 2872 72072
rect 2507 72032 2872 72060
rect 2507 72029 2519 72032
rect 2461 72023 2519 72029
rect 2866 72020 2872 72032
rect 2924 72020 2930 72072
rect 10134 72060 10140 72072
rect 10095 72032 10140 72060
rect 10134 72020 10140 72032
rect 10192 72020 10198 72072
rect 1397 71927 1455 71933
rect 1397 71893 1409 71927
rect 1443 71924 1455 71927
rect 1854 71924 1860 71936
rect 1443 71896 1860 71924
rect 1443 71893 1455 71896
rect 1397 71887 1455 71893
rect 1854 71884 1860 71896
rect 1912 71884 1918 71936
rect 1104 71834 10856 71856
rect 1104 71782 4214 71834
rect 4266 71782 4278 71834
rect 4330 71782 4342 71834
rect 4394 71782 4406 71834
rect 4458 71782 4470 71834
rect 4522 71782 7478 71834
rect 7530 71782 7542 71834
rect 7594 71782 7606 71834
rect 7658 71782 7670 71834
rect 7722 71782 7734 71834
rect 7786 71782 10856 71834
rect 1104 71760 10856 71782
rect 2222 71720 2228 71732
rect 1981 71692 2228 71720
rect 1670 71652 1676 71664
rect 1631 71624 1676 71652
rect 1670 71612 1676 71624
rect 1728 71612 1734 71664
rect 1397 71587 1455 71593
rect 1397 71553 1409 71587
rect 1443 71553 1455 71587
rect 1397 71547 1455 71553
rect 1581 71587 1639 71593
rect 1581 71553 1593 71587
rect 1627 71553 1639 71587
rect 1581 71547 1639 71553
rect 1817 71587 1875 71593
rect 1817 71553 1829 71587
rect 1863 71584 1875 71587
rect 1981 71584 2009 71692
rect 2222 71680 2228 71692
rect 2280 71720 2286 71732
rect 2866 71720 2872 71732
rect 2280 71692 2872 71720
rect 2280 71680 2286 71692
rect 2866 71680 2872 71692
rect 2924 71680 2930 71732
rect 2130 71652 2136 71664
rect 1863 71556 2009 71584
rect 2056 71624 2136 71652
rect 1863 71553 1875 71556
rect 1817 71547 1875 71553
rect 1412 71516 1440 71547
rect 1596 71516 1624 71547
rect 1670 71516 1676 71528
rect 1412 71488 1532 71516
rect 1596 71488 1676 71516
rect 1504 71380 1532 71488
rect 1670 71476 1676 71488
rect 1728 71516 1734 71528
rect 2056 71516 2084 71624
rect 2130 71612 2136 71624
rect 2188 71652 2194 71664
rect 2777 71655 2835 71661
rect 2188 71624 2728 71652
rect 2188 71612 2194 71624
rect 2700 71593 2728 71624
rect 2777 71621 2789 71655
rect 2823 71652 2835 71655
rect 3418 71652 3424 71664
rect 2823 71624 3424 71652
rect 2823 71621 2835 71624
rect 2777 71615 2835 71621
rect 3418 71612 3424 71624
rect 3476 71612 3482 71664
rect 2501 71587 2559 71593
rect 2501 71553 2513 71587
rect 2547 71553 2559 71587
rect 2501 71547 2559 71553
rect 2685 71587 2743 71593
rect 2685 71553 2697 71587
rect 2731 71553 2743 71587
rect 2685 71547 2743 71553
rect 1728 71488 2084 71516
rect 2516 71516 2544 71547
rect 2866 71544 2872 71596
rect 2924 71593 2930 71596
rect 2924 71584 2932 71593
rect 10134 71584 10140 71596
rect 2924 71556 2969 71584
rect 10095 71556 10140 71584
rect 2924 71547 2932 71556
rect 2924 71544 2930 71547
rect 10134 71544 10140 71556
rect 10192 71544 10198 71596
rect 8294 71516 8300 71528
rect 2516 71488 8300 71516
rect 1728 71476 1734 71488
rect 8294 71476 8300 71488
rect 8352 71476 8358 71528
rect 9953 71451 10011 71457
rect 9953 71448 9965 71451
rect 1785 71420 9965 71448
rect 1785 71380 1813 71420
rect 9953 71417 9965 71420
rect 9999 71417 10011 71451
rect 9953 71411 10011 71417
rect 1504 71352 1813 71380
rect 1949 71383 2007 71389
rect 1949 71349 1961 71383
rect 1995 71380 2007 71383
rect 2958 71380 2964 71392
rect 1995 71352 2964 71380
rect 1995 71349 2007 71352
rect 1949 71343 2007 71349
rect 2958 71340 2964 71352
rect 3016 71340 3022 71392
rect 3053 71383 3111 71389
rect 3053 71349 3065 71383
rect 3099 71380 3111 71383
rect 3970 71380 3976 71392
rect 3099 71352 3976 71380
rect 3099 71349 3111 71352
rect 3053 71343 3111 71349
rect 3970 71340 3976 71352
rect 4028 71340 4034 71392
rect 1104 71290 10856 71312
rect 1104 71238 2582 71290
rect 2634 71238 2646 71290
rect 2698 71238 2710 71290
rect 2762 71238 2774 71290
rect 2826 71238 2838 71290
rect 2890 71238 5846 71290
rect 5898 71238 5910 71290
rect 5962 71238 5974 71290
rect 6026 71238 6038 71290
rect 6090 71238 6102 71290
rect 6154 71238 9110 71290
rect 9162 71238 9174 71290
rect 9226 71238 9238 71290
rect 9290 71238 9302 71290
rect 9354 71238 9366 71290
rect 9418 71238 10856 71290
rect 1104 71216 10856 71238
rect 1397 71111 1455 71117
rect 1397 71077 1409 71111
rect 1443 71108 1455 71111
rect 2682 71108 2688 71120
rect 1443 71080 2688 71108
rect 1443 71077 1455 71080
rect 1397 71071 1455 71077
rect 2682 71068 2688 71080
rect 2740 71068 2746 71120
rect 934 70932 940 70984
rect 992 70972 998 70984
rect 1581 70975 1639 70981
rect 1581 70972 1593 70975
rect 992 70944 1593 70972
rect 992 70932 998 70944
rect 1581 70941 1593 70944
rect 1627 70941 1639 70975
rect 2222 70972 2228 70984
rect 2183 70944 2228 70972
rect 1581 70935 1639 70941
rect 2222 70932 2228 70944
rect 2280 70932 2286 70984
rect 2958 70864 2964 70916
rect 3016 70904 3022 70916
rect 3602 70904 3608 70916
rect 3016 70876 3608 70904
rect 3016 70864 3022 70876
rect 3602 70864 3608 70876
rect 3660 70864 3666 70916
rect 1118 70796 1124 70848
rect 1176 70836 1182 70848
rect 1486 70836 1492 70848
rect 1176 70808 1492 70836
rect 1176 70796 1182 70808
rect 1486 70796 1492 70808
rect 1544 70796 1550 70848
rect 2041 70839 2099 70845
rect 2041 70805 2053 70839
rect 2087 70836 2099 70839
rect 2314 70836 2320 70848
rect 2087 70808 2320 70836
rect 2087 70805 2099 70808
rect 2041 70799 2099 70805
rect 2314 70796 2320 70808
rect 2372 70796 2378 70848
rect 1104 70746 10856 70768
rect 1104 70694 4214 70746
rect 4266 70694 4278 70746
rect 4330 70694 4342 70746
rect 4394 70694 4406 70746
rect 4458 70694 4470 70746
rect 4522 70694 7478 70746
rect 7530 70694 7542 70746
rect 7594 70694 7606 70746
rect 7658 70694 7670 70746
rect 7722 70694 7734 70746
rect 7786 70694 10856 70746
rect 1104 70672 10856 70694
rect 9953 70635 10011 70641
rect 9953 70632 9965 70635
rect 1412 70604 9965 70632
rect 1412 70505 1440 70604
rect 9953 70601 9965 70604
rect 9999 70601 10011 70635
rect 9953 70595 10011 70601
rect 1673 70567 1731 70573
rect 1673 70533 1685 70567
rect 1719 70564 1731 70567
rect 3234 70564 3240 70576
rect 1719 70536 3240 70564
rect 1719 70533 1731 70536
rect 1673 70527 1731 70533
rect 3234 70524 3240 70536
rect 3292 70524 3298 70576
rect 1397 70499 1455 70505
rect 1397 70465 1409 70499
rect 1443 70465 1455 70499
rect 1578 70496 1584 70508
rect 1539 70468 1584 70496
rect 1397 70459 1455 70465
rect 1578 70456 1584 70468
rect 1636 70456 1642 70508
rect 1817 70499 1875 70505
rect 1817 70465 1829 70499
rect 1863 70496 1875 70499
rect 2130 70496 2136 70508
rect 1863 70468 2136 70496
rect 1863 70465 1875 70468
rect 1817 70459 1875 70465
rect 2130 70456 2136 70468
rect 2188 70496 2194 70508
rect 10134 70496 10140 70508
rect 2188 70468 3280 70496
rect 10095 70468 10140 70496
rect 2188 70456 2194 70468
rect 3252 70440 3280 70468
rect 10134 70456 10140 70468
rect 10192 70456 10198 70508
rect 1210 70388 1216 70440
rect 1268 70428 1274 70440
rect 1268 70400 1440 70428
rect 1268 70388 1274 70400
rect 1412 70360 1440 70400
rect 3234 70388 3240 70440
rect 3292 70388 3298 70440
rect 1412 70332 1992 70360
rect 1964 70301 1992 70332
rect 1949 70295 2007 70301
rect 1949 70261 1961 70295
rect 1995 70261 2007 70295
rect 1949 70255 2007 70261
rect 1104 70202 10856 70224
rect 1104 70150 2582 70202
rect 2634 70150 2646 70202
rect 2698 70150 2710 70202
rect 2762 70150 2774 70202
rect 2826 70150 2838 70202
rect 2890 70150 5846 70202
rect 5898 70150 5910 70202
rect 5962 70150 5974 70202
rect 6026 70150 6038 70202
rect 6090 70150 6102 70202
rect 6154 70150 9110 70202
rect 9162 70150 9174 70202
rect 9226 70150 9238 70202
rect 9290 70150 9302 70202
rect 9354 70150 9366 70202
rect 9418 70150 10856 70202
rect 1104 70128 10856 70150
rect 1302 70048 1308 70100
rect 1360 70088 1366 70100
rect 1578 70088 1584 70100
rect 1360 70060 1584 70088
rect 1360 70048 1366 70060
rect 1578 70048 1584 70060
rect 1636 70048 1642 70100
rect 1578 69884 1584 69896
rect 1539 69856 1584 69884
rect 1578 69844 1584 69856
rect 1636 69844 1642 69896
rect 1670 69844 1676 69896
rect 1728 69884 1734 69896
rect 2225 69887 2283 69893
rect 2225 69884 2237 69887
rect 1728 69856 2237 69884
rect 1728 69844 1734 69856
rect 2225 69853 2237 69856
rect 2271 69853 2283 69887
rect 10134 69884 10140 69896
rect 10095 69856 10140 69884
rect 2225 69847 2283 69853
rect 10134 69844 10140 69856
rect 10192 69844 10198 69896
rect 1394 69748 1400 69760
rect 1355 69720 1400 69748
rect 1394 69708 1400 69720
rect 1452 69708 1458 69760
rect 1762 69708 1768 69760
rect 1820 69748 1826 69760
rect 2041 69751 2099 69757
rect 2041 69748 2053 69751
rect 1820 69720 2053 69748
rect 1820 69708 1826 69720
rect 2041 69717 2053 69720
rect 2087 69717 2099 69751
rect 9950 69748 9956 69760
rect 9911 69720 9956 69748
rect 2041 69711 2099 69717
rect 9950 69708 9956 69720
rect 10008 69708 10014 69760
rect 1104 69658 10856 69680
rect 1104 69606 4214 69658
rect 4266 69606 4278 69658
rect 4330 69606 4342 69658
rect 4394 69606 4406 69658
rect 4458 69606 4470 69658
rect 4522 69606 7478 69658
rect 7530 69606 7542 69658
rect 7594 69606 7606 69658
rect 7658 69606 7670 69658
rect 7722 69606 7734 69658
rect 7786 69606 10856 69658
rect 1104 69584 10856 69606
rect 566 69436 572 69488
rect 624 69476 630 69488
rect 1854 69476 1860 69488
rect 624 69448 1860 69476
rect 624 69436 630 69448
rect 1854 69436 1860 69448
rect 1912 69436 1918 69488
rect 1578 69408 1584 69420
rect 1539 69380 1584 69408
rect 1578 69368 1584 69380
rect 1636 69368 1642 69420
rect 2222 69408 2228 69420
rect 2183 69380 2228 69408
rect 2222 69368 2228 69380
rect 2280 69368 2286 69420
rect 1394 69300 1400 69352
rect 1452 69340 1458 69352
rect 1670 69340 1676 69352
rect 1452 69312 1676 69340
rect 1452 69300 1458 69312
rect 1670 69300 1676 69312
rect 1728 69300 1734 69352
rect 1394 69204 1400 69216
rect 1355 69176 1400 69204
rect 1394 69164 1400 69176
rect 1452 69164 1458 69216
rect 1854 69164 1860 69216
rect 1912 69204 1918 69216
rect 2041 69207 2099 69213
rect 2041 69204 2053 69207
rect 1912 69176 2053 69204
rect 1912 69164 1918 69176
rect 2041 69173 2053 69176
rect 2087 69173 2099 69207
rect 2041 69167 2099 69173
rect 1104 69114 10856 69136
rect 1104 69062 2582 69114
rect 2634 69062 2646 69114
rect 2698 69062 2710 69114
rect 2762 69062 2774 69114
rect 2826 69062 2838 69114
rect 2890 69062 5846 69114
rect 5898 69062 5910 69114
rect 5962 69062 5974 69114
rect 6026 69062 6038 69114
rect 6090 69062 6102 69114
rect 6154 69062 9110 69114
rect 9162 69062 9174 69114
rect 9226 69062 9238 69114
rect 9290 69062 9302 69114
rect 9354 69062 9366 69114
rect 9418 69062 10856 69114
rect 1104 69040 10856 69062
rect 1949 69003 2007 69009
rect 1949 68969 1961 69003
rect 1995 69000 2007 69003
rect 4890 69000 4896 69012
rect 1995 68972 4896 69000
rect 1995 68969 2007 68972
rect 1949 68963 2007 68969
rect 4890 68960 4896 68972
rect 4948 68960 4954 69012
rect 9950 68864 9956 68876
rect 1412 68836 9956 68864
rect 1412 68805 1440 68836
rect 9950 68824 9956 68836
rect 10008 68824 10014 68876
rect 1397 68799 1455 68805
rect 1397 68765 1409 68799
rect 1443 68765 1455 68799
rect 1397 68759 1455 68765
rect 1486 68756 1492 68808
rect 1544 68796 1550 68808
rect 1673 68799 1731 68805
rect 1673 68796 1685 68799
rect 1544 68768 1685 68796
rect 1544 68756 1550 68768
rect 1673 68765 1685 68768
rect 1719 68765 1731 68799
rect 1673 68759 1731 68765
rect 1817 68799 1875 68805
rect 1817 68765 1829 68799
rect 1863 68765 1875 68799
rect 1817 68759 1875 68765
rect 1302 68688 1308 68740
rect 1360 68728 1366 68740
rect 1581 68731 1639 68737
rect 1581 68728 1593 68731
rect 1360 68700 1593 68728
rect 1360 68688 1366 68700
rect 1581 68697 1593 68700
rect 1627 68697 1639 68731
rect 1832 68728 1860 68759
rect 1946 68756 1952 68808
rect 2004 68796 2010 68808
rect 2222 68796 2228 68808
rect 2004 68768 2228 68796
rect 2004 68756 2010 68768
rect 2222 68756 2228 68768
rect 2280 68756 2286 68808
rect 2685 68799 2743 68805
rect 2685 68765 2697 68799
rect 2731 68796 2743 68799
rect 2774 68796 2780 68808
rect 2731 68768 2780 68796
rect 2731 68765 2743 68768
rect 2685 68759 2743 68765
rect 2774 68756 2780 68768
rect 2832 68756 2838 68808
rect 10134 68796 10140 68808
rect 10095 68768 10140 68796
rect 10134 68756 10140 68768
rect 10192 68756 10198 68808
rect 2590 68728 2596 68740
rect 1832 68700 2596 68728
rect 1581 68691 1639 68697
rect 2590 68688 2596 68700
rect 2648 68688 2654 68740
rect 1486 68620 1492 68672
rect 1544 68660 1550 68672
rect 2501 68663 2559 68669
rect 2501 68660 2513 68663
rect 1544 68632 2513 68660
rect 1544 68620 1550 68632
rect 2501 68629 2513 68632
rect 2547 68629 2559 68663
rect 9950 68660 9956 68672
rect 9911 68632 9956 68660
rect 2501 68623 2559 68629
rect 9950 68620 9956 68632
rect 10008 68620 10014 68672
rect 1104 68570 10856 68592
rect 1104 68518 4214 68570
rect 4266 68518 4278 68570
rect 4330 68518 4342 68570
rect 4394 68518 4406 68570
rect 4458 68518 4470 68570
rect 4522 68518 7478 68570
rect 7530 68518 7542 68570
rect 7594 68518 7606 68570
rect 7658 68518 7670 68570
rect 7722 68518 7734 68570
rect 7786 68518 10856 68570
rect 1104 68496 10856 68518
rect 2038 68456 2044 68468
rect 1688 68428 2044 68456
rect 1302 68348 1308 68400
rect 1360 68388 1366 68400
rect 1688 68397 1716 68428
rect 2038 68416 2044 68428
rect 2096 68416 2102 68468
rect 1581 68391 1639 68397
rect 1581 68388 1593 68391
rect 1360 68360 1593 68388
rect 1360 68348 1366 68360
rect 1581 68357 1593 68360
rect 1627 68357 1639 68391
rect 1581 68351 1639 68357
rect 1673 68391 1731 68397
rect 1673 68357 1685 68391
rect 1719 68357 1731 68391
rect 2590 68388 2596 68400
rect 1673 68351 1731 68357
rect 1832 68360 2596 68388
rect 1832 68329 1860 68360
rect 2590 68348 2596 68360
rect 2648 68388 2654 68400
rect 3234 68388 3240 68400
rect 2648 68360 3240 68388
rect 2648 68348 2654 68360
rect 3234 68348 3240 68360
rect 3292 68348 3298 68400
rect 1397 68323 1455 68329
rect 1397 68289 1409 68323
rect 1443 68289 1455 68323
rect 1397 68283 1455 68289
rect 1817 68323 1875 68329
rect 1817 68289 1829 68323
rect 1863 68289 1875 68323
rect 1817 68283 1875 68289
rect 1412 68252 1440 68283
rect 1946 68280 1952 68332
rect 2004 68320 2010 68332
rect 2406 68320 2412 68332
rect 2004 68292 2412 68320
rect 2004 68280 2010 68292
rect 2406 68280 2412 68292
rect 2464 68280 2470 68332
rect 2685 68323 2743 68329
rect 2685 68289 2697 68323
rect 2731 68320 2743 68323
rect 2958 68320 2964 68332
rect 2731 68292 2964 68320
rect 2731 68289 2743 68292
rect 2685 68283 2743 68289
rect 2958 68280 2964 68292
rect 3016 68280 3022 68332
rect 10134 68320 10140 68332
rect 10095 68292 10140 68320
rect 10134 68280 10140 68292
rect 10192 68280 10198 68332
rect 9950 68252 9956 68264
rect 1412 68224 9956 68252
rect 9950 68212 9956 68224
rect 10008 68212 10014 68264
rect 1949 68187 2007 68193
rect 1949 68153 1961 68187
rect 1995 68184 2007 68187
rect 4614 68184 4620 68196
rect 1995 68156 4620 68184
rect 1995 68153 2007 68156
rect 1949 68147 2007 68153
rect 4614 68144 4620 68156
rect 4672 68144 4678 68196
rect 2406 68076 2412 68128
rect 2464 68116 2470 68128
rect 2501 68119 2559 68125
rect 2501 68116 2513 68119
rect 2464 68088 2513 68116
rect 2464 68076 2470 68088
rect 2501 68085 2513 68088
rect 2547 68085 2559 68119
rect 2501 68079 2559 68085
rect 9858 68076 9864 68128
rect 9916 68116 9922 68128
rect 9953 68119 10011 68125
rect 9953 68116 9965 68119
rect 9916 68088 9965 68116
rect 9916 68076 9922 68088
rect 9953 68085 9965 68088
rect 9999 68085 10011 68119
rect 9953 68079 10011 68085
rect 1104 68026 10856 68048
rect 1104 67974 2582 68026
rect 2634 67974 2646 68026
rect 2698 67974 2710 68026
rect 2762 67974 2774 68026
rect 2826 67974 2838 68026
rect 2890 67974 5846 68026
rect 5898 67974 5910 68026
rect 5962 67974 5974 68026
rect 6026 67974 6038 68026
rect 6090 67974 6102 68026
rect 6154 67974 9110 68026
rect 9162 67974 9174 68026
rect 9226 67974 9238 68026
rect 9290 67974 9302 68026
rect 9354 67974 9366 68026
rect 9418 67974 10856 68026
rect 1104 67952 10856 67974
rect 1397 67847 1455 67853
rect 1397 67813 1409 67847
rect 1443 67844 1455 67847
rect 2038 67844 2044 67856
rect 1443 67816 2044 67844
rect 1443 67813 1455 67816
rect 1397 67807 1455 67813
rect 2038 67804 2044 67816
rect 2096 67804 2102 67856
rect 2777 67847 2835 67853
rect 2777 67813 2789 67847
rect 2823 67844 2835 67847
rect 3694 67844 3700 67856
rect 2823 67816 3700 67844
rect 2823 67813 2835 67816
rect 2777 67807 2835 67813
rect 3694 67804 3700 67816
rect 3752 67804 3758 67856
rect 1302 67736 1308 67788
rect 1360 67776 1366 67788
rect 9950 67776 9956 67788
rect 1360 67748 1716 67776
rect 1360 67736 1366 67748
rect 1578 67708 1584 67720
rect 1539 67680 1584 67708
rect 1578 67668 1584 67680
rect 1636 67668 1642 67720
rect 934 67600 940 67652
rect 992 67640 998 67652
rect 1486 67640 1492 67652
rect 992 67612 1492 67640
rect 992 67600 998 67612
rect 1486 67600 1492 67612
rect 1544 67600 1550 67652
rect 1688 67640 1716 67748
rect 2240 67748 9956 67776
rect 2240 67717 2268 67748
rect 9950 67736 9956 67748
rect 10008 67736 10014 67788
rect 2225 67711 2283 67717
rect 2225 67677 2237 67711
rect 2271 67677 2283 67711
rect 2498 67708 2504 67720
rect 2459 67680 2504 67708
rect 2225 67671 2283 67677
rect 2498 67668 2504 67680
rect 2556 67668 2562 67720
rect 2645 67711 2703 67717
rect 2645 67677 2657 67711
rect 2691 67708 2703 67711
rect 3234 67708 3240 67720
rect 2691 67680 3240 67708
rect 2691 67677 2703 67680
rect 2645 67671 2703 67677
rect 3234 67668 3240 67680
rect 3292 67668 3298 67720
rect 2409 67643 2467 67649
rect 2409 67640 2421 67643
rect 1688 67612 2421 67640
rect 2409 67609 2421 67612
rect 2455 67640 2467 67643
rect 2866 67640 2872 67652
rect 2455 67612 2872 67640
rect 2455 67609 2467 67612
rect 2409 67603 2467 67609
rect 2866 67600 2872 67612
rect 2924 67600 2930 67652
rect 1104 67482 10856 67504
rect 1104 67430 4214 67482
rect 4266 67430 4278 67482
rect 4330 67430 4342 67482
rect 4394 67430 4406 67482
rect 4458 67430 4470 67482
rect 4522 67430 7478 67482
rect 7530 67430 7542 67482
rect 7594 67430 7606 67482
rect 7658 67430 7670 67482
rect 7722 67430 7734 67482
rect 7786 67430 10856 67482
rect 1104 67408 10856 67430
rect 9674 67368 9680 67380
rect 2746 67340 9680 67368
rect 2746 67300 2774 67340
rect 9674 67328 9680 67340
rect 9732 67328 9738 67380
rect 9950 67368 9956 67380
rect 9911 67340 9956 67368
rect 9950 67328 9956 67340
rect 10008 67328 10014 67380
rect 2866 67300 2872 67312
rect 2700 67272 2774 67300
rect 2827 67272 2872 67300
rect 2700 67241 2728 67272
rect 2866 67260 2872 67272
rect 2924 67260 2930 67312
rect 2685 67235 2743 67241
rect 2685 67201 2697 67235
rect 2731 67201 2743 67235
rect 2685 67195 2743 67201
rect 2774 67192 2780 67244
rect 2832 67232 2838 67244
rect 2961 67235 3019 67241
rect 2961 67232 2973 67235
rect 2832 67204 2973 67232
rect 2832 67192 2838 67204
rect 2961 67201 2973 67204
rect 3007 67201 3019 67235
rect 2961 67195 3019 67201
rect 3105 67235 3163 67241
rect 3105 67201 3117 67235
rect 3151 67232 3163 67235
rect 3234 67232 3240 67244
rect 3151 67204 3240 67232
rect 3151 67201 3163 67204
rect 3105 67195 3163 67201
rect 3234 67192 3240 67204
rect 3292 67192 3298 67244
rect 10134 67232 10140 67244
rect 10095 67204 10140 67232
rect 10134 67192 10140 67204
rect 10192 67192 10198 67244
rect 1394 67164 1400 67176
rect 1355 67136 1400 67164
rect 1394 67124 1400 67136
rect 1452 67124 1458 67176
rect 1670 67164 1676 67176
rect 1631 67136 1676 67164
rect 1670 67124 1676 67136
rect 1728 67124 1734 67176
rect 3237 67031 3295 67037
rect 3237 66997 3249 67031
rect 3283 67028 3295 67031
rect 8478 67028 8484 67040
rect 3283 67000 8484 67028
rect 3283 66997 3295 67000
rect 3237 66991 3295 66997
rect 8478 66988 8484 67000
rect 8536 66988 8542 67040
rect 1104 66938 10856 66960
rect 1104 66886 2582 66938
rect 2634 66886 2646 66938
rect 2698 66886 2710 66938
rect 2762 66886 2774 66938
rect 2826 66886 2838 66938
rect 2890 66886 5846 66938
rect 5898 66886 5910 66938
rect 5962 66886 5974 66938
rect 6026 66886 6038 66938
rect 6090 66886 6102 66938
rect 6154 66886 9110 66938
rect 9162 66886 9174 66938
rect 9226 66886 9238 66938
rect 9290 66886 9302 66938
rect 9354 66886 9366 66938
rect 9418 66886 10856 66938
rect 1104 66864 10856 66886
rect 9674 66784 9680 66836
rect 9732 66824 9738 66836
rect 9953 66827 10011 66833
rect 9953 66824 9965 66827
rect 9732 66796 9965 66824
rect 9732 66784 9738 66796
rect 9953 66793 9965 66796
rect 9999 66793 10011 66827
rect 9953 66787 10011 66793
rect 2958 66716 2964 66768
rect 3016 66716 3022 66768
rect 842 66648 848 66700
rect 900 66688 906 66700
rect 1673 66691 1731 66697
rect 1673 66688 1685 66691
rect 900 66660 1685 66688
rect 900 66648 906 66660
rect 1673 66657 1685 66660
rect 1719 66657 1731 66691
rect 2976 66688 3004 66716
rect 3053 66691 3111 66697
rect 3053 66688 3065 66691
rect 2976 66660 3065 66688
rect 1673 66651 1731 66657
rect 3053 66657 3065 66660
rect 3099 66657 3111 66691
rect 3053 66651 3111 66657
rect 1394 66620 1400 66632
rect 1355 66592 1400 66620
rect 1394 66580 1400 66592
rect 1452 66580 1458 66632
rect 2774 66620 2780 66632
rect 2735 66592 2780 66620
rect 2774 66580 2780 66592
rect 2832 66580 2838 66632
rect 10134 66620 10140 66632
rect 10095 66592 10140 66620
rect 10134 66580 10140 66592
rect 10192 66580 10198 66632
rect 1104 66394 10856 66416
rect 1104 66342 4214 66394
rect 4266 66342 4278 66394
rect 4330 66342 4342 66394
rect 4394 66342 4406 66394
rect 4458 66342 4470 66394
rect 4522 66342 7478 66394
rect 7530 66342 7542 66394
rect 7594 66342 7606 66394
rect 7658 66342 7670 66394
rect 7722 66342 7734 66394
rect 7786 66342 10856 66394
rect 1104 66320 10856 66342
rect 3142 66240 3148 66292
rect 3200 66240 3206 66292
rect 2866 66212 2872 66224
rect 2827 66184 2872 66212
rect 2866 66172 2872 66184
rect 2924 66172 2930 66224
rect 2961 66215 3019 66221
rect 2961 66181 2973 66215
rect 3007 66212 3019 66215
rect 3160 66212 3188 66240
rect 3007 66184 3188 66212
rect 3007 66181 3019 66184
rect 2961 66175 3019 66181
rect 198 66104 204 66156
rect 256 66144 262 66156
rect 1673 66147 1731 66153
rect 1673 66144 1685 66147
rect 256 66116 1685 66144
rect 256 66104 262 66116
rect 1673 66113 1685 66116
rect 1719 66113 1731 66147
rect 1673 66107 1731 66113
rect 2685 66147 2743 66153
rect 2685 66113 2697 66147
rect 2731 66113 2743 66147
rect 2685 66107 2743 66113
rect 3105 66147 3163 66153
rect 3105 66113 3117 66147
rect 3151 66144 3163 66147
rect 3234 66144 3240 66156
rect 3151 66116 3240 66144
rect 3151 66113 3163 66116
rect 3105 66107 3163 66113
rect 1394 66076 1400 66088
rect 1355 66048 1400 66076
rect 1394 66036 1400 66048
rect 1452 66036 1458 66088
rect 2700 66076 2728 66107
rect 3234 66104 3240 66116
rect 3292 66104 3298 66156
rect 10134 66144 10140 66156
rect 10095 66116 10140 66144
rect 10134 66104 10140 66116
rect 10192 66104 10198 66156
rect 9858 66076 9864 66088
rect 2700 66048 9864 66076
rect 9858 66036 9864 66048
rect 9916 66036 9922 66088
rect 3234 65940 3240 65952
rect 3195 65912 3240 65940
rect 3234 65900 3240 65912
rect 3292 65900 3298 65952
rect 8294 65900 8300 65952
rect 8352 65940 8358 65952
rect 9953 65943 10011 65949
rect 9953 65940 9965 65943
rect 8352 65912 9965 65940
rect 8352 65900 8358 65912
rect 9953 65909 9965 65912
rect 9999 65909 10011 65943
rect 9953 65903 10011 65909
rect 1104 65850 10856 65872
rect 1104 65798 2582 65850
rect 2634 65798 2646 65850
rect 2698 65798 2710 65850
rect 2762 65798 2774 65850
rect 2826 65798 2838 65850
rect 2890 65798 5846 65850
rect 5898 65798 5910 65850
rect 5962 65798 5974 65850
rect 6026 65798 6038 65850
rect 6090 65798 6102 65850
rect 6154 65798 9110 65850
rect 9162 65798 9174 65850
rect 9226 65798 9238 65850
rect 9290 65798 9302 65850
rect 9354 65798 9366 65850
rect 9418 65798 10856 65850
rect 1104 65776 10856 65798
rect 3878 65628 3884 65680
rect 3936 65668 3942 65680
rect 4982 65668 4988 65680
rect 3936 65640 4988 65668
rect 3936 65628 3942 65640
rect 4982 65628 4988 65640
rect 5040 65628 5046 65680
rect 658 65560 664 65612
rect 716 65600 722 65612
rect 1118 65600 1124 65612
rect 716 65572 1124 65600
rect 716 65560 722 65572
rect 1118 65560 1124 65572
rect 1176 65560 1182 65612
rect 1302 65560 1308 65612
rect 1360 65600 1366 65612
rect 1397 65603 1455 65609
rect 1397 65600 1409 65603
rect 1360 65572 1409 65600
rect 1360 65560 1366 65572
rect 1397 65569 1409 65572
rect 1443 65569 1455 65603
rect 1397 65563 1455 65569
rect 2961 65603 3019 65609
rect 2961 65569 2973 65603
rect 3007 65600 3019 65603
rect 3142 65600 3148 65612
rect 3007 65572 3148 65600
rect 3007 65569 3019 65572
rect 2961 65563 3019 65569
rect 3142 65560 3148 65572
rect 3200 65560 3206 65612
rect 474 65492 480 65544
rect 532 65532 538 65544
rect 1210 65532 1216 65544
rect 532 65504 1216 65532
rect 532 65492 538 65504
rect 1210 65492 1216 65504
rect 1268 65492 1274 65544
rect 1670 65532 1676 65544
rect 1631 65504 1676 65532
rect 1670 65492 1676 65504
rect 1728 65492 1734 65544
rect 2498 65492 2504 65544
rect 2556 65532 2562 65544
rect 2685 65535 2743 65541
rect 2685 65532 2697 65535
rect 2556 65504 2697 65532
rect 2556 65492 2562 65504
rect 2685 65501 2697 65504
rect 2731 65501 2743 65535
rect 2685 65495 2743 65501
rect 3789 65535 3847 65541
rect 3789 65501 3801 65535
rect 3835 65532 3847 65535
rect 4062 65532 4068 65544
rect 3835 65504 4068 65532
rect 3835 65501 3847 65504
rect 3789 65495 3847 65501
rect 4062 65492 4068 65504
rect 4120 65492 4126 65544
rect 3970 65396 3976 65408
rect 3931 65368 3976 65396
rect 3970 65356 3976 65368
rect 4028 65356 4034 65408
rect 1104 65306 10856 65328
rect 1104 65254 4214 65306
rect 4266 65254 4278 65306
rect 4330 65254 4342 65306
rect 4394 65254 4406 65306
rect 4458 65254 4470 65306
rect 4522 65254 7478 65306
rect 7530 65254 7542 65306
rect 7594 65254 7606 65306
rect 7658 65254 7670 65306
rect 7722 65254 7734 65306
rect 7786 65254 10856 65306
rect 1104 65232 10856 65254
rect 1210 65152 1216 65204
rect 1268 65192 1274 65204
rect 2038 65192 2044 65204
rect 1268 65164 2044 65192
rect 1268 65152 1274 65164
rect 2038 65152 2044 65164
rect 2096 65152 2102 65204
rect 3694 65084 3700 65136
rect 3752 65124 3758 65136
rect 3970 65124 3976 65136
rect 3752 65096 3976 65124
rect 3752 65084 3758 65096
rect 3970 65084 3976 65096
rect 4028 65084 4034 65136
rect 1397 65059 1455 65065
rect 1397 65025 1409 65059
rect 1443 65025 1455 65059
rect 1397 65019 1455 65025
rect 1412 64988 1440 65019
rect 2038 65016 2044 65068
rect 2096 65056 2102 65068
rect 2133 65059 2191 65065
rect 2133 65056 2145 65059
rect 2096 65028 2145 65056
rect 2096 65016 2102 65028
rect 2133 65025 2145 65028
rect 2179 65025 2191 65059
rect 2133 65019 2191 65025
rect 2869 65059 2927 65065
rect 2869 65025 2881 65059
rect 2915 65056 2927 65059
rect 2915 65028 3280 65056
rect 2915 65025 2927 65028
rect 2869 65019 2927 65025
rect 3142 64988 3148 65000
rect 1412 64960 1716 64988
rect 1578 64920 1584 64932
rect 1539 64892 1584 64920
rect 1578 64880 1584 64892
rect 1636 64880 1642 64932
rect 1688 64864 1716 64960
rect 2746 64960 3148 64988
rect 2317 64923 2375 64929
rect 2317 64889 2329 64923
rect 2363 64920 2375 64923
rect 2746 64920 2774 64960
rect 3142 64948 3148 64960
rect 3200 64948 3206 65000
rect 3252 64988 3280 65028
rect 3418 65016 3424 65068
rect 3476 65056 3482 65068
rect 3605 65059 3663 65065
rect 3605 65056 3617 65059
rect 3476 65028 3617 65056
rect 3476 65016 3482 65028
rect 3605 65025 3617 65028
rect 3651 65025 3663 65059
rect 10134 65056 10140 65068
rect 10095 65028 10140 65056
rect 3605 65019 3663 65025
rect 10134 65016 10140 65028
rect 10192 65016 10198 65068
rect 3694 64988 3700 65000
rect 3252 64960 3700 64988
rect 3694 64948 3700 64960
rect 3752 64948 3758 65000
rect 3050 64920 3056 64932
rect 2363 64892 2774 64920
rect 3011 64892 3056 64920
rect 2363 64889 2375 64892
rect 2317 64883 2375 64889
rect 3050 64880 3056 64892
rect 3108 64880 3114 64932
rect 3789 64923 3847 64929
rect 3789 64920 3801 64923
rect 3344 64892 3801 64920
rect 3344 64864 3372 64892
rect 3789 64889 3801 64892
rect 3835 64889 3847 64923
rect 3789 64883 3847 64889
rect 8386 64880 8392 64932
rect 8444 64920 8450 64932
rect 9953 64923 10011 64929
rect 9953 64920 9965 64923
rect 8444 64892 9965 64920
rect 8444 64880 8450 64892
rect 9953 64889 9965 64892
rect 9999 64889 10011 64923
rect 9953 64883 10011 64889
rect 1670 64812 1676 64864
rect 1728 64812 1734 64864
rect 3326 64812 3332 64864
rect 3384 64812 3390 64864
rect 1104 64762 10856 64784
rect 1104 64710 2582 64762
rect 2634 64710 2646 64762
rect 2698 64710 2710 64762
rect 2762 64710 2774 64762
rect 2826 64710 2838 64762
rect 2890 64710 5846 64762
rect 5898 64710 5910 64762
rect 5962 64710 5974 64762
rect 6026 64710 6038 64762
rect 6090 64710 6102 64762
rect 6154 64710 9110 64762
rect 9162 64710 9174 64762
rect 9226 64710 9238 64762
rect 9290 64710 9302 64762
rect 9354 64710 9366 64762
rect 9418 64710 10856 64762
rect 1104 64688 10856 64710
rect 8294 64648 8300 64660
rect 1964 64620 8300 64648
rect 1964 64453 1992 64620
rect 8294 64608 8300 64620
rect 8352 64608 8358 64660
rect 2501 64583 2559 64589
rect 2501 64549 2513 64583
rect 2547 64580 2559 64583
rect 4798 64580 4804 64592
rect 2547 64552 4804 64580
rect 2547 64549 2559 64552
rect 2501 64543 2559 64549
rect 4798 64540 4804 64552
rect 4856 64540 4862 64592
rect 1949 64447 2007 64453
rect 1949 64413 1961 64447
rect 1995 64413 2007 64447
rect 2225 64447 2283 64453
rect 2225 64444 2237 64447
rect 1949 64407 2007 64413
rect 2056 64416 2237 64444
rect 1026 64336 1032 64388
rect 1084 64376 1090 64388
rect 2056 64376 2084 64416
rect 2225 64413 2237 64416
rect 2271 64413 2283 64447
rect 2225 64407 2283 64413
rect 2369 64447 2427 64453
rect 2369 64413 2381 64447
rect 2415 64444 2427 64447
rect 10134 64444 10140 64456
rect 2415 64416 3096 64444
rect 10095 64416 10140 64444
rect 2415 64413 2427 64416
rect 2369 64407 2427 64413
rect 1084 64348 2084 64376
rect 2133 64379 2191 64385
rect 1084 64336 1090 64348
rect 2133 64345 2145 64379
rect 2179 64376 2191 64379
rect 2958 64376 2964 64388
rect 2179 64348 2964 64376
rect 2179 64345 2191 64348
rect 2133 64339 2191 64345
rect 2958 64336 2964 64348
rect 3016 64336 3022 64388
rect 3068 64320 3096 64416
rect 10134 64404 10140 64416
rect 10192 64404 10198 64456
rect 3050 64268 3056 64320
rect 3108 64268 3114 64320
rect 8294 64268 8300 64320
rect 8352 64308 8358 64320
rect 9953 64311 10011 64317
rect 9953 64308 9965 64311
rect 8352 64280 9965 64308
rect 8352 64268 8358 64280
rect 9953 64277 9965 64280
rect 9999 64277 10011 64311
rect 9953 64271 10011 64277
rect 1104 64218 10856 64240
rect 1104 64166 4214 64218
rect 4266 64166 4278 64218
rect 4330 64166 4342 64218
rect 4394 64166 4406 64218
rect 4458 64166 4470 64218
rect 4522 64166 7478 64218
rect 7530 64166 7542 64218
rect 7594 64166 7606 64218
rect 7658 64166 7670 64218
rect 7722 64166 7734 64218
rect 7786 64166 10856 64218
rect 1104 64144 10856 64166
rect 2314 64104 2320 64116
rect 2148 64076 2320 64104
rect 2148 64036 2176 64076
rect 2314 64064 2320 64076
rect 2372 64064 2378 64116
rect 2222 64039 2280 64045
rect 2222 64036 2234 64039
rect 2148 64008 2234 64036
rect 2222 64005 2234 64008
rect 2268 64005 2280 64039
rect 2222 63999 2280 64005
rect 1949 63971 2007 63977
rect 1949 63937 1961 63971
rect 1995 63937 2007 63971
rect 1949 63931 2007 63937
rect 2133 63971 2191 63977
rect 2133 63937 2145 63971
rect 2179 63937 2191 63971
rect 2133 63931 2191 63937
rect 2369 63971 2427 63977
rect 2369 63937 2381 63971
rect 2415 63968 2427 63971
rect 3050 63968 3056 63980
rect 2415 63940 3056 63968
rect 2415 63937 2427 63940
rect 2369 63931 2427 63937
rect 1964 63764 1992 63931
rect 2148 63900 2176 63931
rect 3050 63928 3056 63940
rect 3108 63928 3114 63980
rect 2222 63900 2228 63912
rect 2148 63872 2228 63900
rect 2222 63860 2228 63872
rect 2280 63860 2286 63912
rect 8386 63900 8392 63912
rect 2332 63872 8392 63900
rect 2332 63764 2360 63872
rect 8386 63860 8392 63872
rect 8444 63860 8450 63912
rect 1964 63736 2360 63764
rect 2501 63767 2559 63773
rect 2501 63733 2513 63767
rect 2547 63764 2559 63767
rect 5166 63764 5172 63776
rect 2547 63736 5172 63764
rect 2547 63733 2559 63736
rect 2501 63727 2559 63733
rect 5166 63724 5172 63736
rect 5224 63724 5230 63776
rect 1104 63674 10856 63696
rect 1104 63622 2582 63674
rect 2634 63622 2646 63674
rect 2698 63622 2710 63674
rect 2762 63622 2774 63674
rect 2826 63622 2838 63674
rect 2890 63622 5846 63674
rect 5898 63622 5910 63674
rect 5962 63622 5974 63674
rect 6026 63622 6038 63674
rect 6090 63622 6102 63674
rect 6154 63622 9110 63674
rect 9162 63622 9174 63674
rect 9226 63622 9238 63674
rect 9290 63622 9302 63674
rect 9354 63622 9366 63674
rect 9418 63622 10856 63674
rect 1104 63600 10856 63622
rect 2222 63492 2228 63504
rect 1872 63464 2228 63492
rect 1578 63248 1584 63300
rect 1636 63288 1642 63300
rect 1872 63288 1900 63464
rect 2222 63452 2228 63464
rect 2280 63452 2286 63504
rect 2501 63495 2559 63501
rect 2501 63461 2513 63495
rect 2547 63492 2559 63495
rect 3050 63492 3056 63504
rect 2547 63464 3056 63492
rect 2547 63461 2559 63464
rect 2501 63455 2559 63461
rect 3050 63452 3056 63464
rect 3108 63452 3114 63504
rect 3142 63452 3148 63504
rect 3200 63492 3206 63504
rect 3418 63492 3424 63504
rect 3200 63464 3424 63492
rect 3200 63452 3206 63464
rect 3418 63452 3424 63464
rect 3476 63452 3482 63504
rect 8294 63492 8300 63504
rect 6380 63464 8300 63492
rect 6380 63424 6408 63464
rect 8294 63452 8300 63464
rect 8352 63452 8358 63504
rect 1964 63396 6408 63424
rect 1964 63365 1992 63396
rect 1949 63359 2007 63365
rect 1949 63325 1961 63359
rect 1995 63325 2007 63359
rect 2222 63356 2228 63368
rect 2183 63328 2228 63356
rect 1949 63319 2007 63325
rect 2222 63316 2228 63328
rect 2280 63316 2286 63368
rect 2406 63365 2412 63368
rect 2369 63359 2412 63365
rect 2369 63325 2381 63359
rect 2464 63356 2470 63368
rect 2866 63356 2872 63368
rect 2464 63328 2872 63356
rect 2369 63319 2412 63325
rect 2406 63316 2412 63319
rect 2464 63316 2470 63328
rect 2866 63316 2872 63328
rect 2924 63316 2930 63368
rect 3418 63316 3424 63368
rect 3476 63356 3482 63368
rect 3789 63359 3847 63365
rect 3789 63356 3801 63359
rect 3476 63328 3801 63356
rect 3476 63316 3482 63328
rect 3789 63325 3801 63328
rect 3835 63325 3847 63359
rect 9306 63356 9312 63368
rect 9267 63328 9312 63356
rect 3789 63319 3847 63325
rect 9306 63316 9312 63328
rect 9364 63316 9370 63368
rect 9582 63356 9588 63368
rect 9543 63328 9588 63356
rect 9582 63316 9588 63328
rect 9640 63316 9646 63368
rect 2133 63291 2191 63297
rect 2133 63288 2145 63291
rect 1636 63260 2145 63288
rect 1636 63248 1642 63260
rect 2133 63257 2145 63260
rect 2179 63288 2191 63291
rect 2682 63288 2688 63300
rect 2179 63260 2688 63288
rect 2179 63257 2191 63260
rect 2133 63251 2191 63257
rect 2682 63248 2688 63260
rect 2740 63288 2746 63300
rect 2958 63288 2964 63300
rect 2740 63260 2964 63288
rect 2740 63248 2746 63260
rect 2958 63248 2964 63260
rect 3016 63248 3022 63300
rect 3326 63180 3332 63232
rect 3384 63220 3390 63232
rect 3973 63223 4031 63229
rect 3973 63220 3985 63223
rect 3384 63192 3985 63220
rect 3384 63180 3390 63192
rect 3973 63189 3985 63192
rect 4019 63189 4031 63223
rect 3973 63183 4031 63189
rect 1104 63130 10856 63152
rect 1104 63078 4214 63130
rect 4266 63078 4278 63130
rect 4330 63078 4342 63130
rect 4394 63078 4406 63130
rect 4458 63078 4470 63130
rect 4522 63078 7478 63130
rect 7530 63078 7542 63130
rect 7594 63078 7606 63130
rect 7658 63078 7670 63130
rect 7722 63078 7734 63130
rect 7786 63078 10856 63130
rect 1104 63056 10856 63078
rect 1394 62976 1400 63028
rect 1452 62976 1458 63028
rect 4982 63016 4988 63028
rect 2516 62988 4988 63016
rect 1412 62948 1440 62976
rect 1673 62951 1731 62957
rect 1673 62948 1685 62951
rect 1412 62920 1685 62948
rect 1673 62917 1685 62920
rect 1719 62917 1731 62951
rect 1673 62911 1731 62917
rect 1397 62883 1455 62889
rect 1397 62849 1409 62883
rect 1443 62849 1455 62883
rect 1578 62880 1584 62892
rect 1539 62852 1584 62880
rect 1397 62843 1455 62849
rect 1412 62812 1440 62843
rect 1578 62840 1584 62852
rect 1636 62840 1642 62892
rect 1817 62883 1875 62889
rect 1817 62849 1829 62883
rect 1863 62880 1875 62883
rect 2406 62880 2412 62892
rect 1863 62852 2412 62880
rect 1863 62849 1875 62852
rect 1817 62843 1875 62849
rect 2406 62840 2412 62852
rect 2464 62840 2470 62892
rect 2516 62889 2544 62988
rect 4982 62976 4988 62988
rect 5040 62976 5046 63028
rect 2590 62908 2596 62960
rect 2648 62948 2654 62960
rect 2777 62951 2835 62957
rect 2777 62948 2789 62951
rect 2648 62920 2789 62948
rect 2648 62908 2654 62920
rect 2777 62917 2789 62920
rect 2823 62917 2835 62951
rect 2777 62911 2835 62917
rect 3326 62908 3332 62960
rect 3384 62948 3390 62960
rect 3694 62948 3700 62960
rect 3384 62920 3700 62948
rect 3384 62908 3390 62920
rect 3694 62908 3700 62920
rect 3752 62908 3758 62960
rect 2501 62883 2559 62889
rect 2501 62849 2513 62883
rect 2547 62849 2559 62883
rect 2682 62880 2688 62892
rect 2643 62852 2688 62880
rect 2501 62843 2559 62849
rect 2682 62840 2688 62852
rect 2740 62840 2746 62892
rect 2866 62880 2872 62892
rect 2827 62852 2872 62880
rect 2866 62840 2872 62852
rect 2924 62840 2930 62892
rect 3513 62883 3571 62889
rect 3513 62849 3525 62883
rect 3559 62880 3571 62883
rect 5350 62880 5356 62892
rect 3559 62852 5356 62880
rect 3559 62849 3571 62852
rect 3513 62843 3571 62849
rect 5350 62840 5356 62852
rect 5408 62840 5414 62892
rect 10134 62880 10140 62892
rect 10095 62852 10140 62880
rect 10134 62840 10140 62852
rect 10192 62840 10198 62892
rect 1412 62784 9996 62812
rect 1394 62704 1400 62756
rect 1452 62744 1458 62756
rect 1578 62744 1584 62756
rect 1452 62716 1584 62744
rect 1452 62704 1458 62716
rect 1578 62704 1584 62716
rect 1636 62704 1642 62756
rect 3694 62744 3700 62756
rect 3655 62716 3700 62744
rect 3694 62704 3700 62716
rect 3752 62704 3758 62756
rect 9968 62753 9996 62784
rect 9953 62747 10011 62753
rect 9953 62713 9965 62747
rect 9999 62713 10011 62747
rect 9953 62707 10011 62713
rect 1946 62676 1952 62688
rect 1907 62648 1952 62676
rect 1946 62636 1952 62648
rect 2004 62636 2010 62688
rect 3053 62679 3111 62685
rect 3053 62645 3065 62679
rect 3099 62676 3111 62679
rect 5258 62676 5264 62688
rect 3099 62648 5264 62676
rect 3099 62645 3111 62648
rect 3053 62639 3111 62645
rect 5258 62636 5264 62648
rect 5316 62636 5322 62688
rect 1104 62586 10856 62608
rect 1104 62534 2582 62586
rect 2634 62534 2646 62586
rect 2698 62534 2710 62586
rect 2762 62534 2774 62586
rect 2826 62534 2838 62586
rect 2890 62534 5846 62586
rect 5898 62534 5910 62586
rect 5962 62534 5974 62586
rect 6026 62534 6038 62586
rect 6090 62534 6102 62586
rect 6154 62534 9110 62586
rect 9162 62534 9174 62586
rect 9226 62534 9238 62586
rect 9290 62534 9302 62586
rect 9354 62534 9366 62586
rect 9418 62534 10856 62586
rect 1104 62512 10856 62534
rect 1946 62432 1952 62484
rect 2004 62472 2010 62484
rect 3970 62472 3976 62484
rect 2004 62444 3976 62472
rect 2004 62432 2010 62444
rect 3970 62432 3976 62444
rect 4028 62432 4034 62484
rect 2406 62364 2412 62416
rect 2464 62404 2470 62416
rect 2590 62404 2596 62416
rect 2464 62376 2596 62404
rect 2464 62364 2470 62376
rect 2590 62364 2596 62376
rect 2648 62364 2654 62416
rect 1946 62296 1952 62348
rect 2004 62336 2010 62348
rect 2314 62336 2320 62348
rect 2004 62308 2320 62336
rect 2004 62296 2010 62308
rect 2314 62296 2320 62308
rect 2372 62296 2378 62348
rect 14 62228 20 62280
rect 72 62268 78 62280
rect 1397 62271 1455 62277
rect 1397 62268 1409 62271
rect 72 62240 1409 62268
rect 72 62228 78 62240
rect 1397 62237 1409 62240
rect 1443 62237 1455 62271
rect 1397 62231 1455 62237
rect 2133 62271 2191 62277
rect 2133 62237 2145 62271
rect 2179 62237 2191 62271
rect 2133 62231 2191 62237
rect 566 62160 572 62212
rect 624 62200 630 62212
rect 2148 62200 2176 62231
rect 2406 62228 2412 62280
rect 2464 62268 2470 62280
rect 2869 62271 2927 62277
rect 2869 62268 2881 62271
rect 2464 62240 2881 62268
rect 2464 62228 2470 62240
rect 2869 62237 2881 62240
rect 2915 62237 2927 62271
rect 10134 62268 10140 62280
rect 10095 62240 10140 62268
rect 2869 62231 2927 62237
rect 10134 62228 10140 62240
rect 10192 62228 10198 62280
rect 624 62172 2176 62200
rect 624 62160 630 62172
rect 1578 62132 1584 62144
rect 1539 62104 1584 62132
rect 1578 62092 1584 62104
rect 1636 62092 1642 62144
rect 2314 62132 2320 62144
rect 2275 62104 2320 62132
rect 2314 62092 2320 62104
rect 2372 62092 2378 62144
rect 2774 62092 2780 62144
rect 2832 62132 2838 62144
rect 3053 62135 3111 62141
rect 3053 62132 3065 62135
rect 2832 62104 3065 62132
rect 2832 62092 2838 62104
rect 3053 62101 3065 62104
rect 3099 62101 3111 62135
rect 3053 62095 3111 62101
rect 8294 62092 8300 62144
rect 8352 62132 8358 62144
rect 9953 62135 10011 62141
rect 9953 62132 9965 62135
rect 8352 62104 9965 62132
rect 8352 62092 8358 62104
rect 9953 62101 9965 62104
rect 9999 62101 10011 62135
rect 9953 62095 10011 62101
rect 1104 62042 10856 62064
rect 1104 61990 4214 62042
rect 4266 61990 4278 62042
rect 4330 61990 4342 62042
rect 4394 61990 4406 62042
rect 4458 61990 4470 62042
rect 4522 61990 7478 62042
rect 7530 61990 7542 62042
rect 7594 61990 7606 62042
rect 7658 61990 7670 62042
rect 7722 61990 7734 62042
rect 7786 61990 10856 62042
rect 1104 61968 10856 61990
rect 8294 61860 8300 61872
rect 1412 61832 8300 61860
rect 1412 61801 1440 61832
rect 8294 61820 8300 61832
rect 8352 61820 8358 61872
rect 1397 61795 1455 61801
rect 1397 61761 1409 61795
rect 1443 61761 1455 61795
rect 1397 61755 1455 61761
rect 1581 61795 1639 61801
rect 1581 61761 1593 61795
rect 1627 61761 1639 61795
rect 1581 61755 1639 61761
rect 1394 61616 1400 61668
rect 1452 61656 1458 61668
rect 1596 61656 1624 61755
rect 1670 61752 1676 61804
rect 1728 61792 1734 61804
rect 1817 61795 1875 61801
rect 1728 61764 1773 61792
rect 1728 61752 1734 61764
rect 1817 61761 1829 61795
rect 1863 61792 1875 61795
rect 2590 61792 2596 61804
rect 1863 61764 2596 61792
rect 1863 61761 1875 61764
rect 1817 61755 1875 61761
rect 2590 61752 2596 61764
rect 2648 61752 2654 61804
rect 1452 61628 1624 61656
rect 1452 61616 1458 61628
rect 934 61548 940 61600
rect 992 61588 998 61600
rect 1670 61588 1676 61600
rect 992 61560 1676 61588
rect 992 61548 998 61560
rect 1670 61548 1676 61560
rect 1728 61548 1734 61600
rect 1949 61591 2007 61597
rect 1949 61557 1961 61591
rect 1995 61588 2007 61591
rect 2038 61588 2044 61600
rect 1995 61560 2044 61588
rect 1995 61557 2007 61560
rect 1949 61551 2007 61557
rect 2038 61548 2044 61560
rect 2096 61548 2102 61600
rect 1104 61498 10856 61520
rect 1104 61446 2582 61498
rect 2634 61446 2646 61498
rect 2698 61446 2710 61498
rect 2762 61446 2774 61498
rect 2826 61446 2838 61498
rect 2890 61446 5846 61498
rect 5898 61446 5910 61498
rect 5962 61446 5974 61498
rect 6026 61446 6038 61498
rect 6090 61446 6102 61498
rect 6154 61446 9110 61498
rect 9162 61446 9174 61498
rect 9226 61446 9238 61498
rect 9290 61446 9302 61498
rect 9354 61446 9366 61498
rect 9418 61446 10856 61498
rect 1104 61424 10856 61446
rect 1210 61344 1216 61396
rect 1268 61384 1274 61396
rect 1762 61384 1768 61396
rect 1268 61356 1768 61384
rect 1268 61344 1274 61356
rect 1762 61344 1768 61356
rect 1820 61344 1826 61396
rect 1026 61140 1032 61192
rect 1084 61180 1090 61192
rect 1397 61183 1455 61189
rect 1397 61180 1409 61183
rect 1084 61152 1409 61180
rect 1084 61140 1090 61152
rect 1397 61149 1409 61152
rect 1443 61149 1455 61183
rect 1397 61143 1455 61149
rect 2133 61183 2191 61189
rect 2133 61149 2145 61183
rect 2179 61149 2191 61183
rect 10134 61180 10140 61192
rect 10095 61152 10140 61180
rect 2133 61143 2191 61149
rect 934 61072 940 61124
rect 992 61112 998 61124
rect 2148 61112 2176 61143
rect 10134 61140 10140 61152
rect 10192 61140 10198 61192
rect 992 61084 2176 61112
rect 992 61072 998 61084
rect 1578 61044 1584 61056
rect 1539 61016 1584 61044
rect 1578 61004 1584 61016
rect 1636 61004 1642 61056
rect 1946 61004 1952 61056
rect 2004 61044 2010 61056
rect 2130 61044 2136 61056
rect 2004 61016 2136 61044
rect 2004 61004 2010 61016
rect 2130 61004 2136 61016
rect 2188 61004 2194 61056
rect 2314 61044 2320 61056
rect 2275 61016 2320 61044
rect 2314 61004 2320 61016
rect 2372 61004 2378 61056
rect 2774 61004 2780 61056
rect 2832 61044 2838 61056
rect 9953 61047 10011 61053
rect 9953 61044 9965 61047
rect 2832 61016 9965 61044
rect 2832 61004 2838 61016
rect 9953 61013 9965 61016
rect 9999 61013 10011 61047
rect 9953 61007 10011 61013
rect 1104 60954 10856 60976
rect 1104 60902 4214 60954
rect 4266 60902 4278 60954
rect 4330 60902 4342 60954
rect 4394 60902 4406 60954
rect 4458 60902 4470 60954
rect 4522 60902 7478 60954
rect 7530 60902 7542 60954
rect 7594 60902 7606 60954
rect 7658 60902 7670 60954
rect 7722 60902 7734 60954
rect 7786 60902 10856 60954
rect 1104 60880 10856 60902
rect 2774 60840 2780 60852
rect 1504 60812 2780 60840
rect 1397 60707 1455 60713
rect 1397 60673 1409 60707
rect 1443 60704 1455 60707
rect 1504 60704 1532 60812
rect 2774 60800 2780 60812
rect 2832 60800 2838 60852
rect 1581 60775 1639 60781
rect 1581 60741 1593 60775
rect 1627 60741 1639 60775
rect 2314 60772 2320 60784
rect 1581 60735 1639 60741
rect 1872 60744 2320 60772
rect 1443 60676 1532 60704
rect 1443 60673 1455 60676
rect 1397 60667 1455 60673
rect 1596 60636 1624 60735
rect 1673 60707 1731 60713
rect 1673 60673 1685 60707
rect 1719 60673 1731 60707
rect 1673 60667 1731 60673
rect 1770 60707 1828 60713
rect 1770 60673 1782 60707
rect 1816 60704 1828 60707
rect 1872 60704 1900 60744
rect 2314 60732 2320 60744
rect 2372 60732 2378 60784
rect 1816 60676 1900 60704
rect 2501 60707 2559 60713
rect 1816 60673 1828 60676
rect 1770 60667 1828 60673
rect 2501 60673 2513 60707
rect 2547 60704 2559 60707
rect 2547 60676 3004 60704
rect 2547 60673 2559 60676
rect 2501 60667 2559 60673
rect 1412 60608 1624 60636
rect 1688 60636 1716 60667
rect 2976 60648 3004 60676
rect 3050 60664 3056 60716
rect 3108 60704 3114 60716
rect 3970 60704 3976 60716
rect 3108 60676 3976 60704
rect 3108 60664 3114 60676
rect 3970 60664 3976 60676
rect 4028 60664 4034 60716
rect 10134 60704 10140 60716
rect 10095 60676 10140 60704
rect 10134 60664 10140 60676
rect 10192 60664 10198 60716
rect 1854 60636 1860 60648
rect 1688 60608 1860 60636
rect 1412 60580 1440 60608
rect 1854 60596 1860 60608
rect 1912 60596 1918 60648
rect 2958 60596 2964 60648
rect 3016 60596 3022 60648
rect 1394 60528 1400 60580
rect 1452 60528 1458 60580
rect 2685 60571 2743 60577
rect 2685 60537 2697 60571
rect 2731 60568 2743 60571
rect 2774 60568 2780 60580
rect 2731 60540 2780 60568
rect 2731 60537 2743 60540
rect 2685 60531 2743 60537
rect 2774 60528 2780 60540
rect 2832 60528 2838 60580
rect 1854 60460 1860 60512
rect 1912 60500 1918 60512
rect 1949 60503 2007 60509
rect 1949 60500 1961 60503
rect 1912 60472 1961 60500
rect 1912 60460 1918 60472
rect 1949 60469 1961 60472
rect 1995 60469 2007 60503
rect 1949 60463 2007 60469
rect 6914 60460 6920 60512
rect 6972 60500 6978 60512
rect 9953 60503 10011 60509
rect 9953 60500 9965 60503
rect 6972 60472 9965 60500
rect 6972 60460 6978 60472
rect 9953 60469 9965 60472
rect 9999 60469 10011 60503
rect 9953 60463 10011 60469
rect 1104 60410 10856 60432
rect 1104 60358 2582 60410
rect 2634 60358 2646 60410
rect 2698 60358 2710 60410
rect 2762 60358 2774 60410
rect 2826 60358 2838 60410
rect 2890 60358 5846 60410
rect 5898 60358 5910 60410
rect 5962 60358 5974 60410
rect 6026 60358 6038 60410
rect 6090 60358 6102 60410
rect 6154 60358 9110 60410
rect 9162 60358 9174 60410
rect 9226 60358 9238 60410
rect 9290 60358 9302 60410
rect 9354 60358 9366 60410
rect 9418 60358 10856 60410
rect 1104 60336 10856 60358
rect 2869 60299 2927 60305
rect 2869 60265 2881 60299
rect 2915 60296 2927 60299
rect 3142 60296 3148 60308
rect 2915 60268 3148 60296
rect 2915 60265 2927 60268
rect 2869 60259 2927 60265
rect 3142 60256 3148 60268
rect 3200 60256 3206 60308
rect 2958 60188 2964 60240
rect 3016 60228 3022 60240
rect 3016 60200 3188 60228
rect 3016 60188 3022 60200
rect 3160 60172 3188 60200
rect 3142 60120 3148 60172
rect 3200 60120 3206 60172
rect 750 60052 756 60104
rect 808 60092 814 60104
rect 1397 60095 1455 60101
rect 1397 60092 1409 60095
rect 808 60064 1409 60092
rect 808 60052 814 60064
rect 1397 60061 1409 60064
rect 1443 60061 1455 60095
rect 1397 60055 1455 60061
rect 2133 60095 2191 60101
rect 2133 60061 2145 60095
rect 2179 60061 2191 60095
rect 2133 60055 2191 60061
rect 106 59984 112 60036
rect 164 60024 170 60036
rect 2148 60024 2176 60055
rect 2958 60052 2964 60104
rect 3016 60092 3022 60104
rect 3053 60095 3111 60101
rect 3053 60092 3065 60095
rect 3016 60064 3065 60092
rect 3016 60052 3022 60064
rect 3053 60061 3065 60064
rect 3099 60061 3111 60095
rect 3053 60055 3111 60061
rect 164 59996 2176 60024
rect 164 59984 170 59996
rect 1578 59956 1584 59968
rect 1539 59928 1584 59956
rect 1578 59916 1584 59928
rect 1636 59916 1642 59968
rect 2314 59956 2320 59968
rect 2275 59928 2320 59956
rect 2314 59916 2320 59928
rect 2372 59916 2378 59968
rect 1104 59866 10856 59888
rect 1104 59814 4214 59866
rect 4266 59814 4278 59866
rect 4330 59814 4342 59866
rect 4394 59814 4406 59866
rect 4458 59814 4470 59866
rect 4522 59814 7478 59866
rect 7530 59814 7542 59866
rect 7594 59814 7606 59866
rect 7658 59814 7670 59866
rect 7722 59814 7734 59866
rect 7786 59814 10856 59866
rect 1104 59792 10856 59814
rect 382 59576 388 59628
rect 440 59616 446 59628
rect 1397 59619 1455 59625
rect 1397 59616 1409 59619
rect 440 59588 1409 59616
rect 440 59576 446 59588
rect 1397 59585 1409 59588
rect 1443 59585 1455 59619
rect 1397 59579 1455 59585
rect 8294 59576 8300 59628
rect 8352 59616 8358 59628
rect 9585 59619 9643 59625
rect 9585 59616 9597 59619
rect 8352 59588 9597 59616
rect 8352 59576 8358 59588
rect 9585 59585 9597 59588
rect 9631 59585 9643 59619
rect 9585 59579 9643 59585
rect 9306 59548 9312 59560
rect 9267 59520 9312 59548
rect 9306 59508 9312 59520
rect 9364 59508 9370 59560
rect 1394 59372 1400 59424
rect 1452 59412 1458 59424
rect 1581 59415 1639 59421
rect 1581 59412 1593 59415
rect 1452 59384 1593 59412
rect 1452 59372 1458 59384
rect 1581 59381 1593 59384
rect 1627 59381 1639 59415
rect 1581 59375 1639 59381
rect 1104 59322 10856 59344
rect 1104 59270 2582 59322
rect 2634 59270 2646 59322
rect 2698 59270 2710 59322
rect 2762 59270 2774 59322
rect 2826 59270 2838 59322
rect 2890 59270 5846 59322
rect 5898 59270 5910 59322
rect 5962 59270 5974 59322
rect 6026 59270 6038 59322
rect 6090 59270 6102 59322
rect 6154 59270 9110 59322
rect 9162 59270 9174 59322
rect 9226 59270 9238 59322
rect 9290 59270 9302 59322
rect 9354 59270 9366 59322
rect 9418 59270 10856 59322
rect 1104 59248 10856 59270
rect 474 58964 480 59016
rect 532 59004 538 59016
rect 1397 59007 1455 59013
rect 1397 59004 1409 59007
rect 532 58976 1409 59004
rect 532 58964 538 58976
rect 1397 58973 1409 58976
rect 1443 58973 1455 59007
rect 1397 58967 1455 58973
rect 2133 59007 2191 59013
rect 2133 58973 2145 59007
rect 2179 59004 2191 59007
rect 2774 59004 2780 59016
rect 2179 58976 2780 59004
rect 2179 58973 2191 58976
rect 2133 58967 2191 58973
rect 2774 58964 2780 58976
rect 2832 58964 2838 59016
rect 2869 59007 2927 59013
rect 2869 58973 2881 59007
rect 2915 59004 2927 59007
rect 5074 59004 5080 59016
rect 2915 58976 5080 59004
rect 2915 58973 2927 58976
rect 2869 58967 2927 58973
rect 5074 58964 5080 58976
rect 5132 58964 5138 59016
rect 10134 59004 10140 59016
rect 10095 58976 10140 59004
rect 10134 58964 10140 58976
rect 10192 58964 10198 59016
rect 1578 58868 1584 58880
rect 1539 58840 1584 58868
rect 1578 58828 1584 58840
rect 1636 58828 1642 58880
rect 2314 58868 2320 58880
rect 2275 58840 2320 58868
rect 2314 58828 2320 58840
rect 2372 58828 2378 58880
rect 3050 58868 3056 58880
rect 3011 58840 3056 58868
rect 3050 58828 3056 58840
rect 3108 58828 3114 58880
rect 9950 58868 9956 58880
rect 9911 58840 9956 58868
rect 9950 58828 9956 58840
rect 10008 58828 10014 58880
rect 1104 58778 10856 58800
rect 1104 58726 4214 58778
rect 4266 58726 4278 58778
rect 4330 58726 4342 58778
rect 4394 58726 4406 58778
rect 4458 58726 4470 58778
rect 4522 58726 7478 58778
rect 7530 58726 7542 58778
rect 7594 58726 7606 58778
rect 7658 58726 7670 58778
rect 7722 58726 7734 58778
rect 7786 58726 10856 58778
rect 1104 58704 10856 58726
rect 2682 58664 2688 58676
rect 2148 58636 2688 58664
rect 1486 58556 1492 58608
rect 1544 58596 1550 58608
rect 2148 58605 2176 58636
rect 2682 58624 2688 58636
rect 2740 58624 2746 58676
rect 2774 58624 2780 58676
rect 2832 58664 2838 58676
rect 3050 58664 3056 58676
rect 2832 58636 3056 58664
rect 2832 58624 2838 58636
rect 3050 58624 3056 58636
rect 3108 58624 3114 58676
rect 2133 58599 2191 58605
rect 1544 58568 1992 58596
rect 1544 58556 1550 58568
rect 1857 58531 1915 58537
rect 1857 58528 1869 58531
rect 1780 58500 1869 58528
rect 1780 58392 1808 58500
rect 1857 58497 1869 58500
rect 1903 58497 1915 58531
rect 1964 58528 1992 58568
rect 2133 58565 2145 58599
rect 2179 58565 2191 58599
rect 2133 58559 2191 58565
rect 2041 58531 2099 58537
rect 2041 58528 2053 58531
rect 1964 58500 2053 58528
rect 1857 58491 1915 58497
rect 2041 58497 2053 58500
rect 2087 58497 2099 58531
rect 2041 58491 2099 58497
rect 2277 58531 2335 58537
rect 2277 58497 2289 58531
rect 2323 58528 2335 58531
rect 2682 58528 2688 58540
rect 2323 58500 2688 58528
rect 2323 58497 2335 58500
rect 2277 58491 2335 58497
rect 2682 58488 2688 58500
rect 2740 58488 2746 58540
rect 10134 58528 10140 58540
rect 10095 58500 10140 58528
rect 10134 58488 10140 58500
rect 10192 58488 10198 58540
rect 9582 58392 9588 58404
rect 1780 58364 9588 58392
rect 9582 58352 9588 58364
rect 9640 58352 9646 58404
rect 1118 58284 1124 58336
rect 1176 58324 1182 58336
rect 2409 58327 2467 58333
rect 2409 58324 2421 58327
rect 1176 58296 2421 58324
rect 1176 58284 1182 58296
rect 2409 58293 2421 58296
rect 2455 58293 2467 58327
rect 2409 58287 2467 58293
rect 9674 58284 9680 58336
rect 9732 58324 9738 58336
rect 9953 58327 10011 58333
rect 9953 58324 9965 58327
rect 9732 58296 9965 58324
rect 9732 58284 9738 58296
rect 9953 58293 9965 58296
rect 9999 58293 10011 58327
rect 9953 58287 10011 58293
rect 1104 58234 10856 58256
rect 1104 58182 2582 58234
rect 2634 58182 2646 58234
rect 2698 58182 2710 58234
rect 2762 58182 2774 58234
rect 2826 58182 2838 58234
rect 2890 58182 5846 58234
rect 5898 58182 5910 58234
rect 5962 58182 5974 58234
rect 6026 58182 6038 58234
rect 6090 58182 6102 58234
rect 6154 58182 9110 58234
rect 9162 58182 9174 58234
rect 9226 58182 9238 58234
rect 9290 58182 9302 58234
rect 9354 58182 9366 58234
rect 9418 58182 10856 58234
rect 1104 58160 10856 58182
rect 2314 58052 2320 58064
rect 2056 58024 2320 58052
rect 1486 57944 1492 57996
rect 1544 57944 1550 57996
rect 1397 57919 1455 57925
rect 1397 57885 1409 57919
rect 1443 57885 1455 57919
rect 1397 57879 1455 57885
rect 1412 57780 1440 57879
rect 1504 57848 1532 57944
rect 1670 57916 1676 57928
rect 1631 57888 1676 57916
rect 1670 57876 1676 57888
rect 1728 57876 1734 57928
rect 1817 57919 1875 57925
rect 1817 57885 1829 57919
rect 1863 57916 1875 57919
rect 2056 57916 2084 58024
rect 2314 58012 2320 58024
rect 2372 58052 2378 58064
rect 2682 58052 2688 58064
rect 2372 58024 2688 58052
rect 2372 58012 2378 58024
rect 2682 58012 2688 58024
rect 2740 58012 2746 58064
rect 2869 57987 2927 57993
rect 2869 57984 2881 57987
rect 1863 57888 2084 57916
rect 2332 57956 2881 57984
rect 1863 57885 1875 57888
rect 1817 57879 1875 57885
rect 1581 57851 1639 57857
rect 1581 57848 1593 57851
rect 1504 57820 1593 57848
rect 1581 57817 1593 57820
rect 1627 57848 1639 57851
rect 2332 57848 2360 57956
rect 2869 57953 2881 57956
rect 2915 57953 2927 57987
rect 2869 57947 2927 57953
rect 2590 57876 2596 57928
rect 2648 57876 2654 57928
rect 2685 57919 2743 57925
rect 2685 57885 2697 57919
rect 2731 57916 2743 57919
rect 2774 57916 2780 57928
rect 2731 57888 2780 57916
rect 2731 57885 2743 57888
rect 2685 57879 2743 57885
rect 2774 57876 2780 57888
rect 2832 57876 2838 57928
rect 1627 57820 2360 57848
rect 1627 57817 1639 57820
rect 1581 57811 1639 57817
rect 1486 57780 1492 57792
rect 1412 57752 1492 57780
rect 1486 57740 1492 57752
rect 1544 57740 1550 57792
rect 1596 57780 1624 57811
rect 2608 57792 2636 57876
rect 1670 57780 1676 57792
rect 1596 57752 1676 57780
rect 1670 57740 1676 57752
rect 1728 57740 1734 57792
rect 1854 57740 1860 57792
rect 1912 57780 1918 57792
rect 1957 57783 2015 57789
rect 1957 57780 1969 57783
rect 1912 57752 1969 57780
rect 1912 57740 1918 57752
rect 1957 57749 1969 57752
rect 2003 57749 2015 57783
rect 1957 57743 2015 57749
rect 2590 57740 2596 57792
rect 2648 57740 2654 57792
rect 1104 57690 10856 57712
rect 1104 57638 4214 57690
rect 4266 57638 4278 57690
rect 4330 57638 4342 57690
rect 4394 57638 4406 57690
rect 4458 57638 4470 57690
rect 4522 57638 7478 57690
rect 7530 57638 7542 57690
rect 7594 57638 7606 57690
rect 7658 57638 7670 57690
rect 7722 57638 7734 57690
rect 7786 57638 10856 57690
rect 1104 57616 10856 57638
rect 2317 57579 2375 57585
rect 2317 57545 2329 57579
rect 2363 57576 2375 57579
rect 2406 57576 2412 57588
rect 2363 57548 2412 57576
rect 2363 57545 2375 57548
rect 2317 57539 2375 57545
rect 2406 57536 2412 57548
rect 2464 57536 2470 57588
rect 3326 57536 3332 57588
rect 3384 57576 3390 57588
rect 3605 57579 3663 57585
rect 3605 57576 3617 57579
rect 3384 57548 3617 57576
rect 3384 57536 3390 57548
rect 3605 57545 3617 57548
rect 3651 57545 3663 57579
rect 3605 57539 3663 57545
rect 290 57400 296 57452
rect 348 57440 354 57452
rect 1397 57443 1455 57449
rect 1397 57440 1409 57443
rect 348 57412 1409 57440
rect 348 57400 354 57412
rect 1397 57409 1409 57412
rect 1443 57409 1455 57443
rect 2133 57443 2191 57449
rect 2133 57440 2145 57443
rect 1397 57403 1455 57409
rect 1504 57412 2145 57440
rect 1302 57332 1308 57384
rect 1360 57372 1366 57384
rect 1504 57372 1532 57412
rect 2133 57409 2145 57412
rect 2179 57409 2191 57443
rect 2133 57403 2191 57409
rect 2869 57443 2927 57449
rect 2869 57409 2881 57443
rect 2915 57440 2927 57443
rect 3050 57440 3056 57452
rect 2915 57412 3056 57440
rect 2915 57409 2927 57412
rect 2869 57403 2927 57409
rect 3050 57400 3056 57412
rect 3108 57400 3114 57452
rect 3142 57400 3148 57452
rect 3200 57440 3206 57452
rect 3789 57443 3847 57449
rect 3789 57440 3801 57443
rect 3200 57412 3801 57440
rect 3200 57400 3206 57412
rect 3789 57409 3801 57412
rect 3835 57409 3847 57443
rect 3789 57403 3847 57409
rect 1360 57344 1532 57372
rect 9309 57375 9367 57381
rect 1360 57332 1366 57344
rect 9309 57341 9321 57375
rect 9355 57372 9367 57375
rect 9490 57372 9496 57384
rect 9355 57344 9496 57372
rect 9355 57341 9367 57344
rect 9309 57335 9367 57341
rect 9490 57332 9496 57344
rect 9548 57332 9554 57384
rect 9585 57375 9643 57381
rect 9585 57341 9597 57375
rect 9631 57341 9643 57375
rect 9585 57335 9643 57341
rect 2498 57264 2504 57316
rect 2556 57264 2562 57316
rect 2774 57264 2780 57316
rect 2832 57304 2838 57316
rect 3326 57304 3332 57316
rect 2832 57276 3332 57304
rect 2832 57264 2838 57276
rect 3326 57264 3332 57276
rect 3384 57264 3390 57316
rect 6270 57264 6276 57316
rect 6328 57304 6334 57316
rect 9600 57304 9628 57335
rect 6328 57276 9628 57304
rect 6328 57264 6334 57276
rect 1486 57196 1492 57248
rect 1544 57236 1550 57248
rect 1581 57239 1639 57245
rect 1581 57236 1593 57239
rect 1544 57208 1593 57236
rect 1544 57196 1550 57208
rect 1581 57205 1593 57208
rect 1627 57205 1639 57239
rect 1581 57199 1639 57205
rect 2406 57196 2412 57248
rect 2464 57236 2470 57248
rect 2516 57236 2544 57264
rect 3050 57236 3056 57248
rect 2464 57208 2544 57236
rect 3011 57208 3056 57236
rect 2464 57196 2470 57208
rect 3050 57196 3056 57208
rect 3108 57196 3114 57248
rect 1104 57146 10856 57168
rect 1104 57094 2582 57146
rect 2634 57094 2646 57146
rect 2698 57094 2710 57146
rect 2762 57094 2774 57146
rect 2826 57094 2838 57146
rect 2890 57094 5846 57146
rect 5898 57094 5910 57146
rect 5962 57094 5974 57146
rect 6026 57094 6038 57146
rect 6090 57094 6102 57146
rect 6154 57094 9110 57146
rect 9162 57094 9174 57146
rect 9226 57094 9238 57146
rect 9290 57094 9302 57146
rect 9354 57094 9366 57146
rect 9418 57094 10856 57146
rect 1104 57072 10856 57094
rect 2958 57032 2964 57044
rect 1412 57004 2636 57032
rect 2919 57004 2964 57032
rect 1412 56837 1440 57004
rect 1486 56924 1492 56976
rect 1544 56964 1550 56976
rect 1949 56967 2007 56973
rect 1949 56964 1961 56967
rect 1544 56936 1961 56964
rect 1544 56924 1550 56936
rect 1949 56933 1961 56936
rect 1995 56933 2007 56967
rect 2608 56964 2636 57004
rect 2958 56992 2964 57004
rect 3016 56992 3022 57044
rect 3789 57035 3847 57041
rect 3789 57001 3801 57035
rect 3835 57032 3847 57035
rect 4062 57032 4068 57044
rect 3835 57004 4068 57032
rect 3835 57001 3847 57004
rect 3789 56995 3847 57001
rect 4062 56992 4068 57004
rect 4120 56992 4126 57044
rect 9950 56964 9956 56976
rect 2608 56936 9956 56964
rect 1949 56927 2007 56933
rect 9950 56924 9956 56936
rect 10008 56924 10014 56976
rect 2590 56896 2596 56908
rect 1832 56868 2596 56896
rect 1832 56837 1860 56868
rect 2590 56856 2596 56868
rect 2648 56856 2654 56908
rect 6454 56856 6460 56908
rect 6512 56896 6518 56908
rect 9585 56899 9643 56905
rect 9585 56896 9597 56899
rect 6512 56868 9597 56896
rect 6512 56856 6518 56868
rect 9585 56865 9597 56868
rect 9631 56865 9643 56899
rect 9585 56859 9643 56865
rect 1397 56831 1455 56837
rect 1397 56797 1409 56831
rect 1443 56797 1455 56831
rect 1397 56791 1455 56797
rect 1817 56831 1875 56837
rect 1817 56797 1829 56831
rect 1863 56797 1875 56831
rect 2682 56828 2688 56840
rect 2643 56800 2688 56828
rect 1817 56791 1875 56797
rect 2682 56788 2688 56800
rect 2740 56788 2746 56840
rect 2777 56831 2835 56837
rect 2777 56797 2789 56831
rect 2823 56797 2835 56831
rect 3970 56828 3976 56840
rect 3931 56800 3976 56828
rect 2777 56791 2835 56797
rect 1581 56763 1639 56769
rect 1581 56729 1593 56763
rect 1627 56729 1639 56763
rect 1581 56723 1639 56729
rect 1673 56763 1731 56769
rect 1673 56729 1685 56763
rect 1719 56760 1731 56763
rect 2498 56760 2504 56772
rect 1719 56732 2504 56760
rect 1719 56729 1731 56732
rect 1673 56723 1731 56729
rect 1596 56692 1624 56723
rect 2498 56720 2504 56732
rect 2556 56720 2562 56772
rect 1762 56692 1768 56704
rect 1596 56664 1768 56692
rect 1762 56652 1768 56664
rect 1820 56652 1826 56704
rect 2314 56652 2320 56704
rect 2372 56692 2378 56704
rect 2792 56692 2820 56791
rect 3970 56788 3976 56800
rect 4028 56788 4034 56840
rect 9306 56828 9312 56840
rect 9267 56800 9312 56828
rect 9306 56788 9312 56800
rect 9364 56788 9370 56840
rect 2372 56664 2820 56692
rect 2372 56652 2378 56664
rect 1104 56602 10856 56624
rect 1104 56550 4214 56602
rect 4266 56550 4278 56602
rect 4330 56550 4342 56602
rect 4394 56550 4406 56602
rect 4458 56550 4470 56602
rect 4522 56550 7478 56602
rect 7530 56550 7542 56602
rect 7594 56550 7606 56602
rect 7658 56550 7670 56602
rect 7722 56550 7734 56602
rect 7786 56550 10856 56602
rect 1104 56528 10856 56550
rect 2133 56491 2191 56497
rect 2133 56457 2145 56491
rect 2179 56488 2191 56491
rect 3970 56488 3976 56500
rect 2179 56460 3976 56488
rect 2179 56457 2191 56460
rect 2133 56451 2191 56457
rect 3970 56448 3976 56460
rect 4028 56448 4034 56500
rect 2774 56380 2780 56432
rect 2832 56420 2838 56432
rect 2869 56423 2927 56429
rect 2869 56420 2881 56423
rect 2832 56392 2881 56420
rect 2832 56380 2838 56392
rect 2869 56389 2881 56392
rect 2915 56389 2927 56423
rect 2869 56383 2927 56389
rect 3326 56380 3332 56432
rect 3384 56420 3390 56432
rect 4154 56420 4160 56432
rect 3384 56392 4160 56420
rect 3384 56380 3390 56392
rect 842 56312 848 56364
rect 900 56352 906 56364
rect 1210 56352 1216 56364
rect 900 56324 1216 56352
rect 900 56312 906 56324
rect 1210 56312 1216 56324
rect 1268 56312 1274 56364
rect 1949 56355 2007 56361
rect 1949 56321 1961 56355
rect 1995 56352 2007 56355
rect 2593 56355 2651 56361
rect 2593 56352 2605 56355
rect 1995 56324 2605 56352
rect 1995 56321 2007 56324
rect 1949 56315 2007 56321
rect 2593 56321 2605 56324
rect 2639 56352 2651 56355
rect 2958 56352 2964 56364
rect 2639 56324 2964 56352
rect 2639 56321 2651 56324
rect 2593 56315 2651 56321
rect 2958 56312 2964 56324
rect 3016 56312 3022 56364
rect 3712 56361 3740 56392
rect 4154 56380 4160 56392
rect 4212 56380 4218 56432
rect 4706 56380 4712 56432
rect 4764 56420 4770 56432
rect 4982 56420 4988 56432
rect 4764 56392 4988 56420
rect 4764 56380 4770 56392
rect 4982 56380 4988 56392
rect 5040 56380 5046 56432
rect 3697 56355 3755 56361
rect 3697 56321 3709 56355
rect 3743 56321 3755 56355
rect 3697 56315 3755 56321
rect 3881 56355 3939 56361
rect 3881 56321 3893 56355
rect 3927 56352 3939 56355
rect 10137 56355 10195 56361
rect 10137 56352 10149 56355
rect 3927 56324 10149 56352
rect 3927 56321 3939 56324
rect 3881 56315 3939 56321
rect 10137 56321 10149 56324
rect 10183 56321 10195 56355
rect 10137 56315 10195 56321
rect 1765 56287 1823 56293
rect 1765 56253 1777 56287
rect 1811 56253 1823 56287
rect 1765 56247 1823 56253
rect 1780 56216 1808 56247
rect 2866 56244 2872 56296
rect 2924 56284 2930 56296
rect 3513 56287 3571 56293
rect 3513 56284 3525 56287
rect 2924 56256 3525 56284
rect 2924 56244 2930 56256
rect 3513 56253 3525 56256
rect 3559 56284 3571 56287
rect 8570 56284 8576 56296
rect 3559 56256 8576 56284
rect 3559 56253 3571 56256
rect 3513 56247 3571 56253
rect 8570 56244 8576 56256
rect 8628 56244 8634 56296
rect 3326 56216 3332 56228
rect 1780 56188 3332 56216
rect 3326 56176 3332 56188
rect 3384 56176 3390 56228
rect 9950 56148 9956 56160
rect 9911 56120 9956 56148
rect 9950 56108 9956 56120
rect 10008 56108 10014 56160
rect 842 56040 848 56092
rect 900 56080 906 56092
rect 900 56052 980 56080
rect 900 56040 906 56052
rect 566 55904 572 55956
rect 624 55944 630 55956
rect 842 55944 848 55956
rect 624 55916 848 55944
rect 624 55904 630 55916
rect 842 55904 848 55916
rect 900 55904 906 55956
rect 952 55876 980 56052
rect 1104 56058 10856 56080
rect 1104 56006 2582 56058
rect 2634 56006 2646 56058
rect 2698 56006 2710 56058
rect 2762 56006 2774 56058
rect 2826 56006 2838 56058
rect 2890 56006 5846 56058
rect 5898 56006 5910 56058
rect 5962 56006 5974 56058
rect 6026 56006 6038 56058
rect 6090 56006 6102 56058
rect 6154 56006 9110 56058
rect 9162 56006 9174 56058
rect 9226 56006 9238 56058
rect 9290 56006 9302 56058
rect 9354 56006 9366 56058
rect 9418 56006 10856 56058
rect 1104 55984 10856 56006
rect 1581 55947 1639 55953
rect 1581 55944 1593 55947
rect 1504 55916 1593 55944
rect 1504 55876 1532 55916
rect 1581 55913 1593 55916
rect 1627 55913 1639 55947
rect 1581 55907 1639 55913
rect 2777 55947 2835 55953
rect 2777 55913 2789 55947
rect 2823 55944 2835 55947
rect 3142 55944 3148 55956
rect 2823 55916 3148 55944
rect 2823 55913 2835 55916
rect 2777 55907 2835 55913
rect 3142 55904 3148 55916
rect 3200 55904 3206 55956
rect 952 55848 1532 55876
rect 3326 55836 3332 55888
rect 3384 55876 3390 55888
rect 3384 55848 3924 55876
rect 3384 55836 3390 55848
rect 2409 55811 2467 55817
rect 2409 55777 2421 55811
rect 2455 55808 2467 55811
rect 2455 55780 3004 55808
rect 2455 55777 2467 55780
rect 2409 55771 2467 55777
rect 658 55700 664 55752
rect 716 55740 722 55752
rect 1397 55743 1455 55749
rect 1397 55740 1409 55743
rect 716 55712 1409 55740
rect 716 55700 722 55712
rect 1397 55709 1409 55712
rect 1443 55709 1455 55743
rect 1397 55703 1455 55709
rect 2314 55700 2320 55752
rect 2372 55740 2378 55752
rect 2593 55743 2651 55749
rect 2593 55740 2605 55743
rect 2372 55712 2605 55740
rect 2372 55700 2378 55712
rect 2593 55709 2605 55712
rect 2639 55709 2651 55743
rect 2976 55740 3004 55780
rect 3326 55740 3332 55752
rect 2976 55712 3332 55740
rect 2593 55703 2651 55709
rect 3326 55700 3332 55712
rect 3384 55700 3390 55752
rect 3896 55749 3924 55848
rect 3970 55836 3976 55888
rect 4028 55876 4034 55888
rect 4801 55879 4859 55885
rect 4801 55876 4813 55879
rect 4028 55848 4813 55876
rect 4028 55836 4034 55848
rect 4801 55845 4813 55848
rect 4847 55845 4859 55879
rect 4801 55839 4859 55845
rect 5442 55768 5448 55820
rect 5500 55808 5506 55820
rect 9585 55811 9643 55817
rect 9585 55808 9597 55811
rect 5500 55780 9597 55808
rect 5500 55768 5506 55780
rect 9585 55777 9597 55780
rect 9631 55777 9643 55811
rect 9585 55771 9643 55777
rect 3881 55743 3939 55749
rect 3881 55709 3893 55743
rect 3927 55709 3939 55743
rect 3881 55703 3939 55709
rect 3973 55743 4031 55749
rect 3973 55709 3985 55743
rect 4019 55740 4031 55743
rect 4154 55740 4160 55752
rect 4019 55712 4160 55740
rect 4019 55709 4031 55712
rect 3973 55703 4031 55709
rect 3896 55672 3924 55703
rect 4154 55700 4160 55712
rect 4212 55700 4218 55752
rect 4614 55740 4620 55752
rect 4575 55712 4620 55740
rect 4614 55700 4620 55712
rect 4672 55700 4678 55752
rect 9306 55740 9312 55752
rect 9267 55712 9312 55740
rect 9306 55700 9312 55712
rect 9364 55700 9370 55752
rect 6362 55672 6368 55684
rect 3896 55644 6368 55672
rect 6362 55632 6368 55644
rect 6420 55632 6426 55684
rect 3142 55564 3148 55616
rect 3200 55604 3206 55616
rect 3418 55604 3424 55616
rect 3200 55576 3424 55604
rect 3200 55564 3206 55576
rect 3418 55564 3424 55576
rect 3476 55564 3482 55616
rect 4157 55607 4215 55613
rect 4157 55573 4169 55607
rect 4203 55604 4215 55607
rect 10134 55604 10140 55616
rect 4203 55576 10140 55604
rect 4203 55573 4215 55576
rect 4157 55567 4215 55573
rect 10134 55564 10140 55576
rect 10192 55564 10198 55616
rect 1104 55514 10856 55536
rect 1104 55462 4214 55514
rect 4266 55462 4278 55514
rect 4330 55462 4342 55514
rect 4394 55462 4406 55514
rect 4458 55462 4470 55514
rect 4522 55462 7478 55514
rect 7530 55462 7542 55514
rect 7594 55462 7606 55514
rect 7658 55462 7670 55514
rect 7722 55462 7734 55514
rect 7786 55462 10856 55514
rect 1104 55440 10856 55462
rect 1670 55400 1676 55412
rect 1596 55372 1676 55400
rect 1596 55341 1624 55372
rect 1670 55360 1676 55372
rect 1728 55360 1734 55412
rect 1762 55360 1768 55412
rect 1820 55400 1826 55412
rect 1946 55400 1952 55412
rect 1820 55372 1952 55400
rect 1820 55360 1826 55372
rect 1946 55360 1952 55372
rect 2004 55360 2010 55412
rect 3418 55400 3424 55412
rect 3379 55372 3424 55400
rect 3418 55360 3424 55372
rect 3476 55360 3482 55412
rect 5534 55360 5540 55412
rect 5592 55400 5598 55412
rect 9674 55400 9680 55412
rect 5592 55372 9680 55400
rect 5592 55360 5598 55372
rect 9674 55360 9680 55372
rect 9732 55360 9738 55412
rect 1581 55335 1639 55341
rect 1581 55301 1593 55335
rect 1627 55301 1639 55335
rect 1581 55295 1639 55301
rect 1780 55304 2360 55332
rect 1780 55273 1808 55304
rect 1397 55267 1455 55273
rect 1397 55264 1409 55267
rect 1044 55236 1409 55264
rect 1044 54856 1072 55236
rect 1397 55233 1409 55236
rect 1443 55233 1455 55267
rect 1670 55267 1728 55273
rect 1670 55264 1682 55267
rect 1397 55227 1455 55233
rect 1596 55236 1682 55264
rect 1596 55208 1624 55236
rect 1670 55233 1682 55236
rect 1716 55233 1728 55267
rect 1670 55227 1728 55233
rect 1770 55267 1828 55273
rect 1770 55233 1782 55267
rect 1816 55233 1828 55267
rect 1770 55227 1828 55233
rect 2332 55208 2360 55304
rect 2498 55264 2504 55276
rect 2459 55236 2504 55264
rect 2498 55224 2504 55236
rect 2556 55224 2562 55276
rect 3237 55267 3295 55273
rect 3237 55233 3249 55267
rect 3283 55264 3295 55267
rect 4154 55264 4160 55276
rect 3283 55236 4160 55264
rect 3283 55233 3295 55236
rect 3237 55227 3295 55233
rect 4154 55224 4160 55236
rect 4212 55224 4218 55276
rect 9309 55267 9367 55273
rect 9309 55233 9321 55267
rect 9355 55264 9367 55267
rect 9490 55264 9496 55276
rect 9355 55236 9496 55264
rect 9355 55233 9367 55236
rect 9309 55227 9367 55233
rect 9490 55224 9496 55236
rect 9548 55224 9554 55276
rect 1578 55156 1584 55208
rect 1636 55156 1642 55208
rect 2314 55156 2320 55208
rect 2372 55156 2378 55208
rect 2590 55156 2596 55208
rect 2648 55196 2654 55208
rect 2958 55196 2964 55208
rect 2648 55168 2964 55196
rect 2648 55156 2654 55168
rect 2958 55156 2964 55168
rect 3016 55156 3022 55208
rect 2866 55088 2872 55140
rect 2924 55128 2930 55140
rect 2924 55100 3464 55128
rect 2924 55088 2930 55100
rect 3436 55072 3464 55100
rect 1946 55060 1952 55072
rect 1907 55032 1952 55060
rect 1946 55020 1952 55032
rect 2004 55020 2010 55072
rect 2498 55020 2504 55072
rect 2556 55060 2562 55072
rect 2685 55063 2743 55069
rect 2685 55060 2697 55063
rect 2556 55032 2697 55060
rect 2556 55020 2562 55032
rect 2685 55029 2697 55032
rect 2731 55029 2743 55063
rect 2685 55023 2743 55029
rect 3418 55020 3424 55072
rect 3476 55020 3482 55072
rect 6546 55020 6552 55072
rect 6604 55060 6610 55072
rect 9539 55063 9597 55069
rect 9539 55060 9551 55063
rect 6604 55032 9551 55060
rect 6604 55020 6610 55032
rect 9539 55029 9551 55032
rect 9585 55029 9597 55063
rect 9539 55023 9597 55029
rect 1104 54970 10856 54992
rect 1104 54918 2582 54970
rect 2634 54918 2646 54970
rect 2698 54918 2710 54970
rect 2762 54918 2774 54970
rect 2826 54918 2838 54970
rect 2890 54918 5846 54970
rect 5898 54918 5910 54970
rect 5962 54918 5974 54970
rect 6026 54918 6038 54970
rect 6090 54918 6102 54970
rect 6154 54918 9110 54970
rect 9162 54918 9174 54970
rect 9226 54918 9238 54970
rect 9290 54918 9302 54970
rect 9354 54918 9366 54970
rect 9418 54918 10856 54970
rect 1104 54896 10856 54918
rect 5534 54856 5540 54868
rect 1044 54828 5540 54856
rect 5534 54816 5540 54828
rect 5592 54816 5598 54868
rect 8294 54720 8300 54732
rect 1412 54692 8300 54720
rect 1412 54661 1440 54692
rect 8294 54680 8300 54692
rect 8352 54680 8358 54732
rect 1397 54655 1455 54661
rect 1397 54621 1409 54655
rect 1443 54621 1455 54655
rect 1397 54615 1455 54621
rect 1486 54612 1492 54664
rect 1544 54652 1550 54664
rect 1673 54655 1731 54661
rect 1673 54652 1685 54655
rect 1544 54624 1685 54652
rect 1544 54612 1550 54624
rect 1673 54621 1685 54624
rect 1719 54621 1731 54655
rect 1673 54615 1731 54621
rect 1765 54655 1823 54661
rect 1765 54621 1777 54655
rect 1811 54652 1823 54655
rect 2314 54652 2320 54664
rect 1811 54624 2320 54652
rect 1811 54621 1823 54624
rect 1765 54615 1823 54621
rect 2314 54612 2320 54624
rect 2372 54612 2378 54664
rect 2409 54655 2467 54661
rect 2409 54621 2421 54655
rect 2455 54652 2467 54655
rect 6638 54652 6644 54664
rect 2455 54624 6644 54652
rect 2455 54621 2467 54624
rect 2409 54615 2467 54621
rect 6638 54612 6644 54624
rect 6696 54612 6702 54664
rect 10134 54652 10140 54664
rect 10095 54624 10140 54652
rect 10134 54612 10140 54624
rect 10192 54612 10198 54664
rect 1578 54584 1584 54596
rect 1539 54556 1584 54584
rect 1578 54544 1584 54556
rect 1636 54544 1642 54596
rect 1949 54519 2007 54525
rect 1949 54485 1961 54519
rect 1995 54516 2007 54519
rect 2314 54516 2320 54528
rect 1995 54488 2320 54516
rect 1995 54485 2007 54488
rect 1949 54479 2007 54485
rect 2314 54476 2320 54488
rect 2372 54476 2378 54528
rect 2593 54519 2651 54525
rect 2593 54485 2605 54519
rect 2639 54516 2651 54519
rect 2774 54516 2780 54528
rect 2639 54488 2780 54516
rect 2639 54485 2651 54488
rect 2593 54479 2651 54485
rect 2774 54476 2780 54488
rect 2832 54476 2838 54528
rect 9858 54476 9864 54528
rect 9916 54516 9922 54528
rect 9953 54519 10011 54525
rect 9953 54516 9965 54519
rect 9916 54488 9965 54516
rect 9916 54476 9922 54488
rect 9953 54485 9965 54488
rect 9999 54485 10011 54519
rect 9953 54479 10011 54485
rect 1104 54426 10856 54448
rect 1104 54374 4214 54426
rect 4266 54374 4278 54426
rect 4330 54374 4342 54426
rect 4394 54374 4406 54426
rect 4458 54374 4470 54426
rect 4522 54374 7478 54426
rect 7530 54374 7542 54426
rect 7594 54374 7606 54426
rect 7658 54374 7670 54426
rect 7722 54374 7734 54426
rect 7786 54374 10856 54426
rect 1104 54352 10856 54374
rect 2869 54315 2927 54321
rect 2869 54281 2881 54315
rect 2915 54312 2927 54315
rect 3050 54312 3056 54324
rect 2915 54284 3056 54312
rect 2915 54281 2927 54284
rect 2869 54275 2927 54281
rect 3050 54272 3056 54284
rect 3108 54272 3114 54324
rect 2314 54204 2320 54256
rect 2372 54244 2378 54256
rect 10226 54244 10232 54256
rect 2372 54216 10232 54244
rect 2372 54204 2378 54216
rect 10226 54204 10232 54216
rect 10284 54204 10290 54256
rect 1397 54179 1455 54185
rect 1397 54145 1409 54179
rect 1443 54145 1455 54179
rect 1397 54139 1455 54145
rect 2133 54179 2191 54185
rect 2133 54145 2145 54179
rect 2179 54145 2191 54179
rect 3050 54176 3056 54188
rect 3011 54148 3056 54176
rect 2133 54139 2191 54145
rect 1412 54040 1440 54139
rect 2148 54108 2176 54139
rect 3050 54136 3056 54148
rect 3108 54136 3114 54188
rect 9858 54176 9864 54188
rect 9819 54148 9864 54176
rect 9858 54136 9864 54148
rect 9916 54136 9922 54188
rect 4430 54108 4436 54120
rect 2148 54080 4436 54108
rect 4430 54068 4436 54080
rect 4488 54068 4494 54120
rect 4522 54040 4528 54052
rect 1412 54012 4528 54040
rect 4522 54000 4528 54012
rect 4580 54000 4586 54052
rect 10042 54040 10048 54052
rect 10003 54012 10048 54040
rect 10042 54000 10048 54012
rect 10100 54000 10106 54052
rect 1394 53932 1400 53984
rect 1452 53972 1458 53984
rect 1581 53975 1639 53981
rect 1581 53972 1593 53975
rect 1452 53944 1593 53972
rect 1452 53932 1458 53944
rect 1581 53941 1593 53944
rect 1627 53941 1639 53975
rect 2314 53972 2320 53984
rect 2275 53944 2320 53972
rect 1581 53935 1639 53941
rect 2314 53932 2320 53944
rect 2372 53932 2378 53984
rect 1104 53882 10856 53904
rect 1104 53830 2582 53882
rect 2634 53830 2646 53882
rect 2698 53830 2710 53882
rect 2762 53830 2774 53882
rect 2826 53830 2838 53882
rect 2890 53830 5846 53882
rect 5898 53830 5910 53882
rect 5962 53830 5974 53882
rect 6026 53830 6038 53882
rect 6090 53830 6102 53882
rect 6154 53830 9110 53882
rect 9162 53830 9174 53882
rect 9226 53830 9238 53882
rect 9290 53830 9302 53882
rect 9354 53830 9366 53882
rect 9418 53830 10856 53882
rect 1104 53808 10856 53830
rect 1397 53567 1455 53573
rect 1397 53533 1409 53567
rect 1443 53564 1455 53567
rect 1486 53564 1492 53576
rect 1443 53536 1492 53564
rect 1443 53533 1455 53536
rect 1397 53527 1455 53533
rect 1486 53524 1492 53536
rect 1544 53524 1550 53576
rect 9861 53567 9919 53573
rect 9861 53533 9873 53567
rect 9907 53564 9919 53567
rect 9950 53564 9956 53576
rect 9907 53536 9956 53564
rect 9907 53533 9919 53536
rect 9861 53527 9919 53533
rect 9950 53524 9956 53536
rect 10008 53524 10014 53576
rect 1578 53428 1584 53440
rect 1539 53400 1584 53428
rect 1578 53388 1584 53400
rect 1636 53388 1642 53440
rect 10042 53428 10048 53440
rect 10003 53400 10048 53428
rect 10042 53388 10048 53400
rect 10100 53388 10106 53440
rect 1104 53338 10856 53360
rect 1104 53286 4214 53338
rect 4266 53286 4278 53338
rect 4330 53286 4342 53338
rect 4394 53286 4406 53338
rect 4458 53286 4470 53338
rect 4522 53286 7478 53338
rect 7530 53286 7542 53338
rect 7594 53286 7606 53338
rect 7658 53286 7670 53338
rect 7722 53286 7734 53338
rect 7786 53286 10856 53338
rect 1104 53264 10856 53286
rect 2501 53227 2559 53233
rect 2501 53193 2513 53227
rect 2547 53224 2559 53227
rect 3050 53224 3056 53236
rect 2547 53196 3056 53224
rect 2547 53193 2559 53196
rect 2501 53187 2559 53193
rect 3050 53184 3056 53196
rect 3108 53184 3114 53236
rect 9217 53227 9275 53233
rect 9217 53193 9229 53227
rect 9263 53193 9275 53227
rect 9217 53187 9275 53193
rect 3510 53116 3516 53168
rect 3568 53156 3574 53168
rect 3970 53156 3976 53168
rect 3568 53128 3976 53156
rect 3568 53116 3574 53128
rect 3970 53116 3976 53128
rect 4028 53116 4034 53168
rect 5350 53116 5356 53168
rect 5408 53156 5414 53168
rect 6178 53156 6184 53168
rect 5408 53128 6184 53156
rect 5408 53116 5414 53128
rect 6178 53116 6184 53128
rect 6236 53116 6242 53168
rect 9232 53156 9260 53187
rect 9232 53128 9904 53156
rect 1397 53091 1455 53097
rect 1397 53057 1409 53091
rect 1443 53057 1455 53091
rect 2314 53088 2320 53100
rect 2275 53060 2320 53088
rect 1397 53051 1455 53057
rect 1412 52952 1440 53051
rect 2314 53048 2320 53060
rect 2372 53048 2378 53100
rect 2958 53048 2964 53100
rect 3016 53088 3022 53100
rect 9876 53097 9904 53128
rect 3237 53091 3295 53097
rect 3237 53088 3249 53091
rect 3016 53060 3249 53088
rect 3016 53048 3022 53060
rect 3237 53057 3249 53060
rect 3283 53057 3295 53091
rect 3237 53051 3295 53057
rect 3421 53091 3479 53097
rect 3421 53057 3433 53091
rect 3467 53088 3479 53091
rect 9401 53091 9459 53097
rect 9401 53088 9413 53091
rect 3467 53060 9413 53088
rect 3467 53057 3479 53060
rect 3421 53051 3479 53057
rect 9401 53057 9413 53060
rect 9447 53057 9459 53091
rect 9401 53051 9459 53057
rect 9861 53091 9919 53097
rect 9861 53057 9873 53091
rect 9907 53057 9919 53091
rect 9861 53051 9919 53057
rect 2133 53023 2191 53029
rect 2133 52989 2145 53023
rect 2179 53020 2191 53023
rect 2498 53020 2504 53032
rect 2179 52992 2504 53020
rect 2179 52989 2191 52992
rect 2133 52983 2191 52989
rect 2498 52980 2504 52992
rect 2556 52980 2562 53032
rect 3050 53020 3056 53032
rect 3011 52992 3056 53020
rect 3050 52980 3056 52992
rect 3108 53020 3114 53032
rect 3326 53020 3332 53032
rect 3108 52992 3332 53020
rect 3108 52980 3114 52992
rect 3326 52980 3332 52992
rect 3384 52980 3390 53032
rect 5074 52952 5080 52964
rect 1412 52924 5080 52952
rect 5074 52912 5080 52924
rect 5132 52912 5138 52964
rect 1394 52844 1400 52896
rect 1452 52884 1458 52896
rect 1581 52887 1639 52893
rect 1581 52884 1593 52887
rect 1452 52856 1593 52884
rect 1452 52844 1458 52856
rect 1581 52853 1593 52856
rect 1627 52853 1639 52887
rect 10042 52884 10048 52896
rect 10003 52856 10048 52884
rect 1581 52847 1639 52853
rect 10042 52844 10048 52856
rect 10100 52844 10106 52896
rect 1104 52794 10856 52816
rect 1104 52742 2582 52794
rect 2634 52742 2646 52794
rect 2698 52742 2710 52794
rect 2762 52742 2774 52794
rect 2826 52742 2838 52794
rect 2890 52742 5846 52794
rect 5898 52742 5910 52794
rect 5962 52742 5974 52794
rect 6026 52742 6038 52794
rect 6090 52742 6102 52794
rect 6154 52742 9110 52794
rect 9162 52742 9174 52794
rect 9226 52742 9238 52794
rect 9290 52742 9302 52794
rect 9354 52742 9366 52794
rect 9418 52742 10856 52794
rect 1104 52720 10856 52742
rect 2314 52612 2320 52624
rect 2275 52584 2320 52612
rect 2314 52572 2320 52584
rect 2372 52572 2378 52624
rect 1397 52479 1455 52485
rect 1397 52445 1409 52479
rect 1443 52445 1455 52479
rect 1397 52439 1455 52445
rect 2133 52479 2191 52485
rect 2133 52445 2145 52479
rect 2179 52476 2191 52479
rect 5626 52476 5632 52488
rect 2179 52448 5632 52476
rect 2179 52445 2191 52448
rect 2133 52439 2191 52445
rect 1412 52408 1440 52439
rect 5626 52436 5632 52448
rect 5684 52436 5690 52488
rect 10134 52476 10140 52488
rect 10095 52448 10140 52476
rect 10134 52436 10140 52448
rect 10192 52436 10198 52488
rect 2590 52408 2596 52420
rect 1412 52380 2596 52408
rect 2590 52368 2596 52380
rect 2648 52368 2654 52420
rect 1486 52300 1492 52352
rect 1544 52340 1550 52352
rect 1581 52343 1639 52349
rect 1581 52340 1593 52343
rect 1544 52312 1593 52340
rect 1544 52300 1550 52312
rect 1581 52309 1593 52312
rect 1627 52309 1639 52343
rect 1581 52303 1639 52309
rect 9858 52300 9864 52352
rect 9916 52340 9922 52352
rect 9953 52343 10011 52349
rect 9953 52340 9965 52343
rect 9916 52312 9965 52340
rect 9916 52300 9922 52312
rect 9953 52309 9965 52312
rect 9999 52309 10011 52343
rect 9953 52303 10011 52309
rect 1104 52250 10856 52272
rect 1104 52198 4214 52250
rect 4266 52198 4278 52250
rect 4330 52198 4342 52250
rect 4394 52198 4406 52250
rect 4458 52198 4470 52250
rect 4522 52198 7478 52250
rect 7530 52198 7542 52250
rect 7594 52198 7606 52250
rect 7658 52198 7670 52250
rect 7722 52198 7734 52250
rect 7786 52198 10856 52250
rect 1104 52176 10856 52198
rect 2222 52136 2228 52148
rect 2183 52108 2228 52136
rect 2222 52096 2228 52108
rect 2280 52096 2286 52148
rect 4065 52139 4123 52145
rect 4065 52105 4077 52139
rect 4111 52136 4123 52139
rect 10134 52136 10140 52148
rect 4111 52108 10140 52136
rect 4111 52105 4123 52108
rect 4065 52099 4123 52105
rect 10134 52096 10140 52108
rect 10192 52096 10198 52148
rect 1397 52003 1455 52009
rect 1397 51969 1409 52003
rect 1443 52000 1455 52003
rect 2222 52000 2228 52012
rect 1443 51972 2228 52000
rect 1443 51969 1455 51972
rect 1397 51963 1455 51969
rect 2222 51960 2228 51972
rect 2280 51960 2286 52012
rect 2406 52000 2412 52012
rect 2367 51972 2412 52000
rect 2406 51960 2412 51972
rect 2464 51960 2470 52012
rect 2958 51960 2964 52012
rect 3016 52000 3022 52012
rect 3053 52003 3111 52009
rect 3053 52000 3065 52003
rect 3016 51972 3065 52000
rect 3016 51960 3022 51972
rect 3053 51969 3065 51972
rect 3099 52000 3111 52003
rect 3326 52000 3332 52012
rect 3099 51972 3332 52000
rect 3099 51969 3111 51972
rect 3053 51963 3111 51969
rect 3326 51960 3332 51972
rect 3384 52000 3390 52012
rect 3881 52003 3939 52009
rect 3881 52000 3893 52003
rect 3384 51972 3893 52000
rect 3384 51960 3390 51972
rect 3881 51969 3893 51972
rect 3927 51969 3939 52003
rect 9858 52000 9864 52012
rect 9819 51972 9864 52000
rect 3881 51963 3939 51969
rect 9858 51960 9864 51972
rect 9916 51960 9922 52012
rect 2498 51892 2504 51944
rect 2556 51932 2562 51944
rect 2869 51935 2927 51941
rect 2869 51932 2881 51935
rect 2556 51904 2881 51932
rect 2556 51892 2562 51904
rect 2869 51901 2881 51904
rect 2915 51901 2927 51935
rect 3697 51935 3755 51941
rect 3697 51932 3709 51935
rect 2869 51895 2927 51901
rect 2976 51904 3709 51932
rect 2976 51876 3004 51904
rect 3697 51901 3709 51904
rect 3743 51901 3755 51935
rect 3697 51895 3755 51901
rect 2958 51824 2964 51876
rect 3016 51824 3022 51876
rect 3237 51867 3295 51873
rect 3237 51833 3249 51867
rect 3283 51864 3295 51867
rect 10134 51864 10140 51876
rect 3283 51836 10140 51864
rect 3283 51833 3295 51836
rect 3237 51827 3295 51833
rect 10134 51824 10140 51836
rect 10192 51824 10198 51876
rect 1578 51796 1584 51808
rect 1539 51768 1584 51796
rect 1578 51756 1584 51768
rect 1636 51756 1642 51808
rect 10042 51796 10048 51808
rect 10003 51768 10048 51796
rect 10042 51756 10048 51768
rect 10100 51756 10106 51808
rect 1104 51706 10856 51728
rect 1104 51654 2582 51706
rect 2634 51654 2646 51706
rect 2698 51654 2710 51706
rect 2762 51654 2774 51706
rect 2826 51654 2838 51706
rect 2890 51654 5846 51706
rect 5898 51654 5910 51706
rect 5962 51654 5974 51706
rect 6026 51654 6038 51706
rect 6090 51654 6102 51706
rect 6154 51654 9110 51706
rect 9162 51654 9174 51706
rect 9226 51654 9238 51706
rect 9290 51654 9302 51706
rect 9354 51654 9366 51706
rect 9418 51654 10856 51706
rect 1104 51632 10856 51654
rect 2406 51552 2412 51604
rect 2464 51592 2470 51604
rect 2777 51595 2835 51601
rect 2777 51592 2789 51595
rect 2464 51564 2789 51592
rect 2464 51552 2470 51564
rect 2777 51561 2789 51564
rect 2823 51561 2835 51595
rect 2777 51555 2835 51561
rect 1118 51524 1124 51536
rect 584 51496 1124 51524
rect 584 51468 612 51496
rect 1118 51484 1124 51496
rect 1176 51484 1182 51536
rect 566 51416 572 51468
rect 624 51416 630 51468
rect 1762 51416 1768 51468
rect 1820 51416 1826 51468
rect 2314 51416 2320 51468
rect 2372 51456 2378 51468
rect 2372 51428 2636 51456
rect 2372 51416 2378 51428
rect 1118 51348 1124 51400
rect 1176 51388 1182 51400
rect 1397 51391 1455 51397
rect 1397 51388 1409 51391
rect 1176 51360 1409 51388
rect 1176 51348 1182 51360
rect 1397 51357 1409 51360
rect 1443 51357 1455 51391
rect 1780 51388 1808 51416
rect 2406 51388 2412 51400
rect 1780 51360 2412 51388
rect 1397 51351 1455 51357
rect 2406 51348 2412 51360
rect 2464 51348 2470 51400
rect 2608 51397 2636 51428
rect 2501 51391 2559 51397
rect 2501 51357 2513 51391
rect 2547 51357 2559 51391
rect 2501 51351 2559 51357
rect 2593 51391 2651 51397
rect 2593 51357 2605 51391
rect 2639 51388 2651 51391
rect 3050 51388 3056 51400
rect 2639 51360 3056 51388
rect 2639 51357 2651 51360
rect 2593 51351 2651 51357
rect 2516 51320 2544 51351
rect 3050 51348 3056 51360
rect 3108 51348 3114 51400
rect 9858 51388 9864 51400
rect 9819 51360 9864 51388
rect 9858 51348 9864 51360
rect 9916 51348 9922 51400
rect 2958 51320 2964 51332
rect 2516 51292 2964 51320
rect 2958 51280 2964 51292
rect 3016 51280 3022 51332
rect 1578 51252 1584 51264
rect 1539 51224 1584 51252
rect 1578 51212 1584 51224
rect 1636 51212 1642 51264
rect 10042 51252 10048 51264
rect 10003 51224 10048 51252
rect 10042 51212 10048 51224
rect 10100 51212 10106 51264
rect 1104 51162 10856 51184
rect 1104 51110 4214 51162
rect 4266 51110 4278 51162
rect 4330 51110 4342 51162
rect 4394 51110 4406 51162
rect 4458 51110 4470 51162
rect 4522 51110 7478 51162
rect 7530 51110 7542 51162
rect 7594 51110 7606 51162
rect 7658 51110 7670 51162
rect 7722 51110 7734 51162
rect 7786 51110 10856 51162
rect 1104 51088 10856 51110
rect 1302 51048 1308 51060
rect 124 51020 1308 51048
rect 124 50300 152 51020
rect 1302 51008 1308 51020
rect 1360 51008 1366 51060
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 3970 51048 3976 51060
rect 3476 51020 3976 51048
rect 3476 51008 3482 51020
rect 3970 51008 3976 51020
rect 4028 51008 4034 51060
rect 5166 51008 5172 51060
rect 5224 51048 5230 51060
rect 6730 51048 6736 51060
rect 5224 51020 6736 51048
rect 5224 51008 5230 51020
rect 6730 51008 6736 51020
rect 6788 51008 6794 51060
rect 9858 51008 9864 51060
rect 9916 51048 9922 51060
rect 9953 51051 10011 51057
rect 9953 51048 9965 51051
rect 9916 51020 9965 51048
rect 9916 51008 9922 51020
rect 9953 51017 9965 51020
rect 9999 51017 10011 51051
rect 9953 51011 10011 51017
rect 1210 50980 1216 50992
rect 1044 50952 1216 50980
rect 1044 50504 1072 50952
rect 1210 50940 1216 50952
rect 1268 50940 1274 50992
rect 5258 50940 5264 50992
rect 5316 50940 5322 50992
rect 1397 50915 1455 50921
rect 1397 50912 1409 50915
rect 1228 50884 1409 50912
rect 1228 50856 1256 50884
rect 1397 50881 1409 50884
rect 1443 50881 1455 50915
rect 1397 50875 1455 50881
rect 2133 50915 2191 50921
rect 2133 50881 2145 50915
rect 2179 50881 2191 50915
rect 2133 50875 2191 50881
rect 1210 50804 1216 50856
rect 1268 50804 1274 50856
rect 1302 50804 1308 50856
rect 1360 50844 1366 50856
rect 2148 50844 2176 50875
rect 3786 50872 3792 50924
rect 3844 50912 3850 50924
rect 4062 50912 4068 50924
rect 3844 50884 4068 50912
rect 3844 50872 3850 50884
rect 4062 50872 4068 50884
rect 4120 50872 4126 50924
rect 1360 50816 2176 50844
rect 5276 50844 5304 50940
rect 10134 50912 10140 50924
rect 10095 50884 10140 50912
rect 10134 50872 10140 50884
rect 10192 50872 10198 50924
rect 5626 50844 5632 50856
rect 5276 50816 5632 50844
rect 1360 50804 1366 50816
rect 5626 50804 5632 50816
rect 5684 50804 5690 50856
rect 1581 50779 1639 50785
rect 1581 50776 1593 50779
rect 1320 50748 1593 50776
rect 1320 50720 1348 50748
rect 1581 50745 1593 50748
rect 1627 50745 1639 50779
rect 1581 50739 1639 50745
rect 1946 50736 1952 50788
rect 2004 50776 2010 50788
rect 2317 50779 2375 50785
rect 2317 50776 2329 50779
rect 2004 50748 2329 50776
rect 2004 50736 2010 50748
rect 2317 50745 2329 50748
rect 2363 50745 2375 50779
rect 2317 50739 2375 50745
rect 1302 50668 1308 50720
rect 1360 50668 1366 50720
rect 1104 50618 10856 50640
rect 1104 50566 2582 50618
rect 2634 50566 2646 50618
rect 2698 50566 2710 50618
rect 2762 50566 2774 50618
rect 2826 50566 2838 50618
rect 2890 50566 5846 50618
rect 5898 50566 5910 50618
rect 5962 50566 5974 50618
rect 6026 50566 6038 50618
rect 6090 50566 6102 50618
rect 6154 50566 9110 50618
rect 9162 50566 9174 50618
rect 9226 50566 9238 50618
rect 9290 50566 9302 50618
rect 9354 50566 9366 50618
rect 9418 50566 10856 50618
rect 1104 50544 10856 50566
rect 1302 50504 1308 50516
rect 1044 50476 1308 50504
rect 1302 50464 1308 50476
rect 1360 50464 1366 50516
rect 1412 50476 1808 50504
rect 198 50396 204 50448
rect 256 50436 262 50448
rect 256 50408 980 50436
rect 256 50396 262 50408
rect 750 50328 756 50380
rect 808 50328 814 50380
rect 198 50300 204 50312
rect 124 50272 204 50300
rect 198 50260 204 50272
rect 256 50260 262 50312
rect 768 50028 796 50328
rect 952 50232 980 50408
rect 1412 50309 1440 50476
rect 1780 50436 1808 50476
rect 4706 50464 4712 50516
rect 4764 50504 4770 50516
rect 6822 50504 6828 50516
rect 4764 50476 6828 50504
rect 4764 50464 4770 50476
rect 6822 50464 6828 50476
rect 6880 50464 6886 50516
rect 6546 50436 6552 50448
rect 1780 50408 6552 50436
rect 6546 50396 6552 50408
rect 6604 50396 6610 50448
rect 1946 50368 1952 50380
rect 1680 50340 1952 50368
rect 1397 50303 1455 50309
rect 1397 50269 1409 50303
rect 1443 50269 1455 50303
rect 1397 50263 1455 50269
rect 1486 50260 1492 50312
rect 1544 50300 1550 50312
rect 1581 50303 1639 50309
rect 1581 50300 1593 50303
rect 1544 50272 1593 50300
rect 1544 50260 1550 50272
rect 1581 50269 1593 50272
rect 1627 50300 1639 50303
rect 1680 50300 1708 50340
rect 1946 50328 1952 50340
rect 2004 50328 2010 50380
rect 4706 50328 4712 50380
rect 4764 50368 4770 50380
rect 4982 50368 4988 50380
rect 4764 50340 4988 50368
rect 4764 50328 4770 50340
rect 4982 50328 4988 50340
rect 5040 50328 5046 50380
rect 1627 50272 1708 50300
rect 1627 50269 1639 50272
rect 1581 50263 1639 50269
rect 1762 50260 1768 50312
rect 1820 50300 1826 50312
rect 2409 50303 2467 50309
rect 1820 50272 1865 50300
rect 1820 50260 1826 50272
rect 2409 50269 2421 50303
rect 2455 50300 2467 50303
rect 5534 50300 5540 50312
rect 2455 50272 5540 50300
rect 2455 50269 2467 50272
rect 2409 50263 2467 50269
rect 5534 50260 5540 50272
rect 5592 50260 5598 50312
rect 9858 50300 9864 50312
rect 9819 50272 9864 50300
rect 9858 50260 9864 50272
rect 9916 50260 9922 50312
rect 1673 50235 1731 50241
rect 1673 50232 1685 50235
rect 952 50204 1685 50232
rect 1673 50201 1685 50204
rect 1719 50201 1731 50235
rect 1673 50195 1731 50201
rect 1946 50164 1952 50176
rect 1907 50136 1952 50164
rect 1946 50124 1952 50136
rect 2004 50124 2010 50176
rect 2593 50167 2651 50173
rect 2593 50133 2605 50167
rect 2639 50164 2651 50167
rect 2774 50164 2780 50176
rect 2639 50136 2780 50164
rect 2639 50133 2651 50136
rect 2593 50127 2651 50133
rect 2774 50124 2780 50136
rect 2832 50124 2838 50176
rect 10042 50164 10048 50176
rect 10003 50136 10048 50164
rect 10042 50124 10048 50136
rect 10100 50124 10106 50176
rect 1104 50074 10856 50096
rect 934 50028 940 50040
rect 768 50000 940 50028
rect 934 49988 940 50000
rect 992 49988 998 50040
rect 1104 50022 4214 50074
rect 4266 50022 4278 50074
rect 4330 50022 4342 50074
rect 4394 50022 4406 50074
rect 4458 50022 4470 50074
rect 4522 50022 7478 50074
rect 7530 50022 7542 50074
rect 7594 50022 7606 50074
rect 7658 50022 7670 50074
rect 7722 50022 7734 50074
rect 7786 50022 10856 50074
rect 1104 50000 10856 50022
rect 3145 49963 3203 49969
rect 3145 49929 3157 49963
rect 3191 49960 3203 49963
rect 3234 49960 3240 49972
rect 3191 49932 3240 49960
rect 3191 49929 3203 49932
rect 3145 49923 3203 49929
rect 3234 49920 3240 49932
rect 3292 49920 3298 49972
rect 9582 49920 9588 49972
rect 9640 49960 9646 49972
rect 10045 49963 10103 49969
rect 10045 49960 10057 49963
rect 9640 49932 10057 49960
rect 9640 49920 9646 49932
rect 10045 49929 10057 49932
rect 10091 49929 10103 49963
rect 10045 49923 10103 49929
rect 1670 49892 1676 49904
rect 1631 49864 1676 49892
rect 1670 49852 1676 49864
rect 1728 49852 1734 49904
rect 4522 49892 4528 49904
rect 2746 49864 4528 49892
rect 1397 49827 1455 49833
rect 1397 49793 1409 49827
rect 1443 49793 1455 49827
rect 1397 49787 1455 49793
rect 1412 49756 1440 49787
rect 1486 49784 1492 49836
rect 1544 49824 1550 49836
rect 1581 49827 1639 49833
rect 1581 49824 1593 49827
rect 1544 49796 1593 49824
rect 1544 49784 1550 49796
rect 1581 49793 1593 49796
rect 1627 49793 1639 49827
rect 1762 49824 1768 49836
rect 1723 49796 1768 49824
rect 1581 49787 1639 49793
rect 1762 49784 1768 49796
rect 1820 49784 1826 49836
rect 2409 49827 2467 49833
rect 2409 49793 2421 49827
rect 2455 49824 2467 49827
rect 2746 49824 2774 49864
rect 4522 49852 4528 49864
rect 4580 49852 4586 49904
rect 2455 49796 2774 49824
rect 3329 49827 3387 49833
rect 2455 49793 2467 49796
rect 2409 49787 2467 49793
rect 3329 49793 3341 49827
rect 3375 49793 3387 49827
rect 3329 49787 3387 49793
rect 1412 49728 3280 49756
rect 1946 49620 1952 49632
rect 1907 49592 1952 49620
rect 1946 49580 1952 49592
rect 2004 49580 2010 49632
rect 2222 49580 2228 49632
rect 2280 49620 2286 49632
rect 2593 49623 2651 49629
rect 2593 49620 2605 49623
rect 2280 49592 2605 49620
rect 2280 49580 2286 49592
rect 2593 49589 2605 49592
rect 2639 49589 2651 49623
rect 3252 49620 3280 49728
rect 3344 49700 3372 49787
rect 9674 49784 9680 49836
rect 9732 49824 9738 49836
rect 9861 49827 9919 49833
rect 9861 49824 9873 49827
rect 9732 49796 9873 49824
rect 9732 49784 9738 49796
rect 9861 49793 9873 49796
rect 9907 49793 9919 49827
rect 9861 49787 9919 49793
rect 3326 49648 3332 49700
rect 3384 49648 3390 49700
rect 6270 49620 6276 49632
rect 3252 49592 6276 49620
rect 2593 49583 2651 49589
rect 6270 49580 6276 49592
rect 6328 49580 6334 49632
rect 1104 49530 10856 49552
rect 1104 49478 2582 49530
rect 2634 49478 2646 49530
rect 2698 49478 2710 49530
rect 2762 49478 2774 49530
rect 2826 49478 2838 49530
rect 2890 49478 5846 49530
rect 5898 49478 5910 49530
rect 5962 49478 5974 49530
rect 6026 49478 6038 49530
rect 6090 49478 6102 49530
rect 6154 49478 9110 49530
rect 9162 49478 9174 49530
rect 9226 49478 9238 49530
rect 9290 49478 9302 49530
rect 9354 49478 9366 49530
rect 9418 49478 10856 49530
rect 1104 49456 10856 49478
rect 2777 49419 2835 49425
rect 2777 49385 2789 49419
rect 2823 49416 2835 49419
rect 3326 49416 3332 49428
rect 2823 49388 3332 49416
rect 2823 49385 2835 49388
rect 2777 49379 2835 49385
rect 3326 49376 3332 49388
rect 3384 49376 3390 49428
rect 3510 49376 3516 49428
rect 3568 49416 3574 49428
rect 3568 49388 3924 49416
rect 3568 49376 3574 49388
rect 3896 49360 3924 49388
rect 2498 49308 2504 49360
rect 2556 49348 2562 49360
rect 3234 49348 3240 49360
rect 2556 49320 3240 49348
rect 2556 49308 2562 49320
rect 3234 49308 3240 49320
rect 3292 49308 3298 49360
rect 3878 49308 3884 49360
rect 3936 49308 3942 49360
rect 5258 49280 5264 49292
rect 1412 49252 5264 49280
rect 1412 49221 1440 49252
rect 5258 49240 5264 49252
rect 5316 49240 5322 49292
rect 1397 49215 1455 49221
rect 1397 49181 1409 49215
rect 1443 49181 1455 49215
rect 1397 49175 1455 49181
rect 1486 49172 1492 49224
rect 1544 49212 1550 49224
rect 1581 49215 1639 49221
rect 1581 49212 1593 49215
rect 1544 49184 1593 49212
rect 1544 49172 1550 49184
rect 1581 49181 1593 49184
rect 1627 49181 1639 49215
rect 1762 49212 1768 49224
rect 1723 49184 1768 49212
rect 1581 49175 1639 49181
rect 1762 49172 1768 49184
rect 1820 49172 1826 49224
rect 2409 49215 2467 49221
rect 2409 49181 2421 49215
rect 2455 49181 2467 49215
rect 2409 49175 2467 49181
rect 2593 49215 2651 49221
rect 2593 49181 2605 49215
rect 2639 49212 2651 49215
rect 2774 49212 2780 49224
rect 2639 49184 2780 49212
rect 2639 49181 2651 49184
rect 2593 49175 2651 49181
rect 1670 49104 1676 49156
rect 1728 49144 1734 49156
rect 2424 49144 2452 49175
rect 2774 49172 2780 49184
rect 2832 49212 2838 49224
rect 3050 49212 3056 49224
rect 2832 49184 3056 49212
rect 2832 49172 2838 49184
rect 3050 49172 3056 49184
rect 3108 49172 3114 49224
rect 3789 49215 3847 49221
rect 3789 49181 3801 49215
rect 3835 49212 3847 49215
rect 3970 49212 3976 49224
rect 3835 49184 3976 49212
rect 3835 49181 3847 49184
rect 3789 49175 3847 49181
rect 3970 49172 3976 49184
rect 4028 49172 4034 49224
rect 9861 49215 9919 49221
rect 9861 49181 9873 49215
rect 9907 49212 9919 49215
rect 9950 49212 9956 49224
rect 9907 49184 9956 49212
rect 9907 49181 9919 49184
rect 9861 49175 9919 49181
rect 9950 49172 9956 49184
rect 10008 49172 10014 49224
rect 2682 49144 2688 49156
rect 1728 49116 1773 49144
rect 2424 49116 2688 49144
rect 1728 49104 1734 49116
rect 2682 49104 2688 49116
rect 2740 49104 2746 49156
rect 2866 49104 2872 49156
rect 2924 49144 2930 49156
rect 6454 49144 6460 49156
rect 2924 49116 6460 49144
rect 2924 49104 2930 49116
rect 6454 49104 6460 49116
rect 6512 49104 6518 49156
rect 1394 49036 1400 49088
rect 1452 49076 1458 49088
rect 1949 49079 2007 49085
rect 1949 49076 1961 49079
rect 1452 49048 1961 49076
rect 1452 49036 1458 49048
rect 1949 49045 1961 49048
rect 1995 49045 2007 49079
rect 3970 49076 3976 49088
rect 3931 49048 3976 49076
rect 1949 49039 2007 49045
rect 3970 49036 3976 49048
rect 4028 49036 4034 49088
rect 10042 49076 10048 49088
rect 10003 49048 10048 49076
rect 10042 49036 10048 49048
rect 10100 49036 10106 49088
rect 1104 48986 10856 49008
rect 1104 48934 4214 48986
rect 4266 48934 4278 48986
rect 4330 48934 4342 48986
rect 4394 48934 4406 48986
rect 4458 48934 4470 48986
rect 4522 48934 7478 48986
rect 7530 48934 7542 48986
rect 7594 48934 7606 48986
rect 7658 48934 7670 48986
rect 7722 48934 7734 48986
rect 7786 48934 10856 48986
rect 1104 48912 10856 48934
rect 1949 48875 2007 48881
rect 1949 48841 1961 48875
rect 1995 48872 2007 48875
rect 3050 48872 3056 48884
rect 1995 48844 3056 48872
rect 1995 48841 2007 48844
rect 1949 48835 2007 48841
rect 3050 48832 3056 48844
rect 3108 48832 3114 48884
rect 3145 48875 3203 48881
rect 3145 48841 3157 48875
rect 3191 48872 3203 48875
rect 3191 48844 3556 48872
rect 3191 48841 3203 48844
rect 3145 48835 3203 48841
rect 2866 48804 2872 48816
rect 1412 48776 2872 48804
rect 1412 48745 1440 48776
rect 2866 48764 2872 48776
rect 2924 48764 2930 48816
rect 3326 48764 3332 48816
rect 3384 48764 3390 48816
rect 3528 48804 3556 48844
rect 3602 48832 3608 48884
rect 3660 48872 3666 48884
rect 3660 48844 4108 48872
rect 3660 48832 3666 48844
rect 3528 48776 4016 48804
rect 1397 48739 1455 48745
rect 1397 48705 1409 48739
rect 1443 48705 1455 48739
rect 1397 48699 1455 48705
rect 1486 48696 1492 48748
rect 1544 48736 1550 48748
rect 1581 48739 1639 48745
rect 1581 48736 1593 48739
rect 1544 48708 1593 48736
rect 1544 48696 1550 48708
rect 1581 48705 1593 48708
rect 1627 48705 1639 48739
rect 1581 48699 1639 48705
rect 1673 48739 1731 48745
rect 1673 48705 1685 48739
rect 1719 48705 1731 48739
rect 1673 48699 1731 48705
rect 1302 48628 1308 48680
rect 1360 48668 1366 48680
rect 1688 48668 1716 48699
rect 1762 48696 1768 48748
rect 1820 48736 1826 48748
rect 2777 48739 2835 48745
rect 2777 48736 2789 48739
rect 1820 48708 1865 48736
rect 2148 48708 2789 48736
rect 1820 48696 1826 48708
rect 1360 48640 1716 48668
rect 1360 48628 1366 48640
rect 1670 48600 1676 48612
rect 1320 48572 1676 48600
rect 1320 48544 1348 48572
rect 1670 48560 1676 48572
rect 1728 48600 1734 48612
rect 2148 48600 2176 48708
rect 2777 48705 2789 48708
rect 2823 48705 2835 48739
rect 2777 48699 2835 48705
rect 2961 48739 3019 48745
rect 2961 48705 2973 48739
rect 3007 48736 3019 48739
rect 3142 48736 3148 48748
rect 3007 48708 3148 48736
rect 3007 48705 3019 48708
rect 2961 48699 3019 48705
rect 3142 48696 3148 48708
rect 3200 48696 3206 48748
rect 3344 48680 3372 48764
rect 3418 48696 3424 48748
rect 3476 48696 3482 48748
rect 3605 48739 3663 48745
rect 3605 48705 3617 48739
rect 3651 48736 3663 48739
rect 3651 48708 3924 48736
rect 3651 48705 3663 48708
rect 3605 48699 3663 48705
rect 3326 48628 3332 48680
rect 3384 48628 3390 48680
rect 1728 48572 2176 48600
rect 1728 48560 1734 48572
rect 2314 48560 2320 48612
rect 2372 48560 2378 48612
rect 3050 48560 3056 48612
rect 3108 48600 3114 48612
rect 3108 48572 3372 48600
rect 3108 48560 3114 48572
rect 1302 48492 1308 48544
rect 1360 48492 1366 48544
rect 1486 48492 1492 48544
rect 1544 48532 1550 48544
rect 2332 48532 2360 48560
rect 3344 48544 3372 48572
rect 3436 48544 3464 48696
rect 1544 48504 2360 48532
rect 1544 48492 1550 48504
rect 3326 48492 3332 48544
rect 3384 48492 3390 48544
rect 3418 48492 3424 48544
rect 3476 48492 3482 48544
rect 3786 48532 3792 48544
rect 3747 48504 3792 48532
rect 3786 48492 3792 48504
rect 3844 48492 3850 48544
rect 3896 48532 3924 48708
rect 3988 48668 4016 48776
rect 4080 48748 4108 48844
rect 9858 48832 9864 48884
rect 9916 48872 9922 48884
rect 9953 48875 10011 48881
rect 9953 48872 9965 48875
rect 9916 48844 9965 48872
rect 9916 48832 9922 48844
rect 9953 48841 9965 48844
rect 9999 48841 10011 48875
rect 9953 48835 10011 48841
rect 9646 48776 10180 48804
rect 4062 48696 4068 48748
rect 4120 48696 4126 48748
rect 9646 48668 9674 48776
rect 10152 48745 10180 48776
rect 10137 48739 10195 48745
rect 10137 48705 10149 48739
rect 10183 48705 10195 48739
rect 10137 48699 10195 48705
rect 3988 48640 9674 48668
rect 4522 48560 4528 48612
rect 4580 48600 4586 48612
rect 5534 48600 5540 48612
rect 4580 48572 5540 48600
rect 4580 48560 4586 48572
rect 5534 48560 5540 48572
rect 5592 48560 5598 48612
rect 8478 48532 8484 48544
rect 3896 48504 8484 48532
rect 8478 48492 8484 48504
rect 8536 48492 8542 48544
rect 1104 48442 10856 48464
rect 1104 48390 2582 48442
rect 2634 48390 2646 48442
rect 2698 48390 2710 48442
rect 2762 48390 2774 48442
rect 2826 48390 2838 48442
rect 2890 48390 5846 48442
rect 5898 48390 5910 48442
rect 5962 48390 5974 48442
rect 6026 48390 6038 48442
rect 6090 48390 6102 48442
rect 6154 48390 9110 48442
rect 9162 48390 9174 48442
rect 9226 48390 9238 48442
rect 9290 48390 9302 48442
rect 9354 48390 9366 48442
rect 9418 48390 10856 48442
rect 1104 48368 10856 48390
rect 2222 48288 2228 48340
rect 2280 48328 2286 48340
rect 2280 48300 2544 48328
rect 2280 48288 2286 48300
rect 2516 48272 2544 48300
rect 842 48260 848 48272
rect 676 48232 848 48260
rect 676 47988 704 48232
rect 842 48220 848 48232
rect 900 48220 906 48272
rect 2498 48220 2504 48272
rect 2556 48220 2562 48272
rect 3694 48220 3700 48272
rect 3752 48260 3758 48272
rect 4338 48260 4344 48272
rect 3752 48232 4344 48260
rect 3752 48220 3758 48232
rect 4338 48220 4344 48232
rect 4396 48220 4402 48272
rect 9217 48263 9275 48269
rect 9217 48229 9229 48263
rect 9263 48260 9275 48263
rect 9674 48260 9680 48272
rect 9263 48232 9680 48260
rect 9263 48229 9275 48232
rect 9217 48223 9275 48229
rect 9674 48220 9680 48232
rect 9732 48220 9738 48272
rect 750 48152 756 48204
rect 808 48192 814 48204
rect 2685 48195 2743 48201
rect 2685 48192 2697 48195
rect 808 48164 2697 48192
rect 808 48152 814 48164
rect 2685 48161 2697 48164
rect 2731 48161 2743 48195
rect 2685 48155 2743 48161
rect 4522 48152 4528 48204
rect 4580 48192 4586 48204
rect 7098 48192 7104 48204
rect 4580 48164 7104 48192
rect 4580 48152 4586 48164
rect 7098 48152 7104 48164
rect 7156 48152 7162 48204
rect 934 48084 940 48136
rect 992 48084 998 48136
rect 1397 48127 1455 48133
rect 1397 48093 1409 48127
rect 1443 48093 1455 48127
rect 2406 48124 2412 48136
rect 2367 48096 2412 48124
rect 1397 48087 1455 48093
rect 750 48016 756 48068
rect 808 48056 814 48068
rect 952 48056 980 48084
rect 808 48028 980 48056
rect 1412 48056 1440 48087
rect 2406 48084 2412 48096
rect 2464 48084 2470 48136
rect 5258 48084 5264 48136
rect 5316 48124 5322 48136
rect 9401 48127 9459 48133
rect 9401 48124 9413 48127
rect 5316 48096 9413 48124
rect 5316 48084 5322 48096
rect 9401 48093 9413 48096
rect 9447 48093 9459 48127
rect 9401 48087 9459 48093
rect 9490 48084 9496 48136
rect 9548 48124 9554 48136
rect 9861 48127 9919 48133
rect 9861 48124 9873 48127
rect 9548 48096 9873 48124
rect 9548 48084 9554 48096
rect 9861 48093 9873 48096
rect 9907 48093 9919 48127
rect 9861 48087 9919 48093
rect 7006 48056 7012 48068
rect 1412 48028 7012 48056
rect 808 48016 814 48028
rect 7006 48016 7012 48028
rect 7064 48016 7070 48068
rect 842 47988 848 48000
rect 676 47960 848 47988
rect 842 47948 848 47960
rect 900 47948 906 48000
rect 1578 47988 1584 48000
rect 1539 47960 1584 47988
rect 1578 47948 1584 47960
rect 1636 47948 1642 48000
rect 10042 47988 10048 48000
rect 10003 47960 10048 47988
rect 10042 47948 10048 47960
rect 10100 47948 10106 48000
rect 1104 47898 10856 47920
rect 1104 47846 4214 47898
rect 4266 47846 4278 47898
rect 4330 47846 4342 47898
rect 4394 47846 4406 47898
rect 4458 47846 4470 47898
rect 4522 47846 7478 47898
rect 7530 47846 7542 47898
rect 7594 47846 7606 47898
rect 7658 47846 7670 47898
rect 7722 47846 7734 47898
rect 7786 47846 10856 47898
rect 1104 47824 10856 47846
rect 1946 47676 1952 47728
rect 2004 47716 2010 47728
rect 2314 47716 2320 47728
rect 2004 47688 2320 47716
rect 2004 47676 2010 47688
rect 2314 47676 2320 47688
rect 2372 47676 2378 47728
rect 1394 47648 1400 47660
rect 1355 47620 1400 47648
rect 1394 47608 1400 47620
rect 1452 47608 1458 47660
rect 2869 47651 2927 47657
rect 2869 47617 2881 47651
rect 2915 47648 2927 47651
rect 3786 47648 3792 47660
rect 2915 47620 3792 47648
rect 2915 47617 2927 47620
rect 2869 47611 2927 47617
rect 3786 47608 3792 47620
rect 3844 47608 3850 47660
rect 8294 47608 8300 47660
rect 8352 47648 8358 47660
rect 9861 47651 9919 47657
rect 9861 47648 9873 47651
rect 8352 47620 9873 47648
rect 8352 47608 8358 47620
rect 9861 47617 9873 47620
rect 9907 47617 9919 47651
rect 9861 47611 9919 47617
rect 1946 47540 1952 47592
rect 2004 47580 2010 47592
rect 2593 47583 2651 47589
rect 2593 47580 2605 47583
rect 2004 47552 2605 47580
rect 2004 47540 2010 47552
rect 2593 47549 2605 47552
rect 2639 47549 2651 47583
rect 2593 47543 2651 47549
rect 1578 47444 1584 47456
rect 1539 47416 1584 47444
rect 1578 47404 1584 47416
rect 1636 47404 1642 47456
rect 3786 47404 3792 47456
rect 3844 47444 3850 47456
rect 3970 47444 3976 47456
rect 3844 47416 3976 47444
rect 3844 47404 3850 47416
rect 3970 47404 3976 47416
rect 4028 47404 4034 47456
rect 10042 47444 10048 47456
rect 10003 47416 10048 47444
rect 10042 47404 10048 47416
rect 10100 47404 10106 47456
rect 1104 47354 10856 47376
rect 1104 47302 2582 47354
rect 2634 47302 2646 47354
rect 2698 47302 2710 47354
rect 2762 47302 2774 47354
rect 2826 47302 2838 47354
rect 2890 47302 5846 47354
rect 5898 47302 5910 47354
rect 5962 47302 5974 47354
rect 6026 47302 6038 47354
rect 6090 47302 6102 47354
rect 6154 47302 9110 47354
rect 9162 47302 9174 47354
rect 9226 47302 9238 47354
rect 9290 47302 9302 47354
rect 9354 47302 9366 47354
rect 9418 47302 10856 47354
rect 1104 47280 10856 47302
rect 1578 47200 1584 47252
rect 1636 47240 1642 47252
rect 1762 47240 1768 47252
rect 1636 47212 1768 47240
rect 1636 47200 1642 47212
rect 1762 47200 1768 47212
rect 1820 47200 1826 47252
rect 1946 47240 1952 47252
rect 1907 47212 1952 47240
rect 1946 47200 1952 47212
rect 2004 47200 2010 47252
rect 2406 47200 2412 47252
rect 2464 47240 2470 47252
rect 2777 47243 2835 47249
rect 2777 47240 2789 47243
rect 2464 47212 2789 47240
rect 2464 47200 2470 47212
rect 2777 47209 2789 47212
rect 2823 47209 2835 47243
rect 2777 47203 2835 47209
rect 7745 47243 7803 47249
rect 7745 47209 7757 47243
rect 7791 47240 7803 47243
rect 9490 47240 9496 47252
rect 7791 47212 9496 47240
rect 7791 47209 7803 47212
rect 7745 47203 7803 47209
rect 9490 47200 9496 47212
rect 9548 47200 9554 47252
rect 9950 47240 9956 47252
rect 9911 47212 9956 47240
rect 9950 47200 9956 47212
rect 10008 47200 10014 47252
rect 3970 47172 3976 47184
rect 3931 47144 3976 47172
rect 3970 47132 3976 47144
rect 4028 47132 4034 47184
rect 4430 47132 4436 47184
rect 4488 47172 4494 47184
rect 6454 47172 6460 47184
rect 4488 47144 6460 47172
rect 4488 47132 4494 47144
rect 6454 47132 6460 47144
rect 6512 47132 6518 47184
rect 1780 47076 2636 47104
rect 1780 47045 1808 47076
rect 1673 47039 1731 47045
rect 1673 47005 1685 47039
rect 1719 47005 1731 47039
rect 1673 46999 1731 47005
rect 1765 47039 1823 47045
rect 1765 47005 1777 47039
rect 1811 47005 1823 47039
rect 2498 47036 2504 47048
rect 2459 47008 2504 47036
rect 1765 46999 1823 47005
rect 1688 46968 1716 46999
rect 2498 46996 2504 47008
rect 2556 46996 2562 47048
rect 2608 47045 2636 47076
rect 2682 47064 2688 47116
rect 2740 47104 2746 47116
rect 5537 47107 5595 47113
rect 5537 47104 5549 47107
rect 2740 47076 5549 47104
rect 2740 47064 2746 47076
rect 5537 47073 5549 47076
rect 5583 47073 5595 47107
rect 6546 47104 6552 47116
rect 5537 47067 5595 47073
rect 5736 47076 6552 47104
rect 2593 47039 2651 47045
rect 2593 47005 2605 47039
rect 2639 47036 2651 47039
rect 2958 47036 2964 47048
rect 2639 47008 2964 47036
rect 2639 47005 2651 47008
rect 2593 46999 2651 47005
rect 2958 46996 2964 47008
rect 3016 46996 3022 47048
rect 3789 47039 3847 47045
rect 3789 47005 3801 47039
rect 3835 47036 3847 47039
rect 4430 47036 4436 47048
rect 3835 47008 4436 47036
rect 3835 47005 3847 47008
rect 3789 46999 3847 47005
rect 4430 46996 4436 47008
rect 4488 46996 4494 47048
rect 5736 47045 5764 47076
rect 6546 47064 6552 47076
rect 6604 47064 6610 47116
rect 4525 47039 4583 47045
rect 4525 47005 4537 47039
rect 4571 47005 4583 47039
rect 4525 46999 4583 47005
rect 4709 47039 4767 47045
rect 4709 47005 4721 47039
rect 4755 47036 4767 47039
rect 5721 47039 5779 47045
rect 5721 47036 5733 47039
rect 4755 47008 5733 47036
rect 4755 47005 4767 47008
rect 4709 46999 4767 47005
rect 5721 47005 5733 47008
rect 5767 47005 5779 47039
rect 5721 46999 5779 47005
rect 5905 47039 5963 47045
rect 5905 47005 5917 47039
rect 5951 47036 5963 47039
rect 7929 47039 7987 47045
rect 7929 47036 7941 47039
rect 5951 47008 7941 47036
rect 5951 47005 5963 47008
rect 5905 46999 5963 47005
rect 7929 47005 7941 47008
rect 7975 47005 7987 47039
rect 7929 46999 7987 47005
rect 10137 47039 10195 47045
rect 10137 47005 10149 47039
rect 10183 47005 10195 47039
rect 10137 46999 10195 47005
rect 4246 46968 4252 46980
rect 1688 46940 4252 46968
rect 4246 46928 4252 46940
rect 4304 46968 4310 46980
rect 4540 46968 4568 46999
rect 4304 46940 4568 46968
rect 4893 46971 4951 46977
rect 4304 46928 4310 46940
rect 4893 46937 4905 46971
rect 4939 46968 4951 46971
rect 10152 46968 10180 46999
rect 4939 46940 10180 46968
rect 4939 46937 4951 46940
rect 4893 46931 4951 46937
rect 1104 46810 10856 46832
rect 14 46724 20 46776
rect 72 46764 78 46776
rect 72 46736 888 46764
rect 1104 46758 4214 46810
rect 4266 46758 4278 46810
rect 4330 46758 4342 46810
rect 4394 46758 4406 46810
rect 4458 46758 4470 46810
rect 4522 46758 7478 46810
rect 7530 46758 7542 46810
rect 7594 46758 7606 46810
rect 7658 46758 7670 46810
rect 7722 46758 7734 46810
rect 7786 46758 10856 46810
rect 1104 46736 10856 46758
rect 72 46724 78 46736
rect 750 46696 756 46708
rect 676 46668 756 46696
rect 676 46504 704 46668
rect 750 46656 756 46668
rect 808 46656 814 46708
rect 860 46628 888 46736
rect 3050 46656 3056 46708
rect 3108 46696 3114 46708
rect 3418 46696 3424 46708
rect 3108 46668 3424 46696
rect 3108 46656 3114 46668
rect 3418 46656 3424 46668
rect 3476 46656 3482 46708
rect 7837 46699 7895 46705
rect 7837 46665 7849 46699
rect 7883 46696 7895 46699
rect 8294 46696 8300 46708
rect 7883 46668 8300 46696
rect 7883 46665 7895 46668
rect 7837 46659 7895 46665
rect 8294 46656 8300 46668
rect 8352 46656 8358 46708
rect 860 46600 2268 46628
rect 2240 46569 2268 46600
rect 2225 46563 2283 46569
rect 2225 46529 2237 46563
rect 2271 46529 2283 46563
rect 2225 46523 2283 46529
rect 3237 46563 3295 46569
rect 3237 46529 3249 46563
rect 3283 46560 3295 46563
rect 3418 46560 3424 46572
rect 3283 46532 3424 46560
rect 3283 46529 3295 46532
rect 3237 46523 3295 46529
rect 3418 46520 3424 46532
rect 3476 46520 3482 46572
rect 6546 46560 6552 46572
rect 6507 46532 6552 46560
rect 6546 46520 6552 46532
rect 6604 46520 6610 46572
rect 6733 46563 6791 46569
rect 6733 46529 6745 46563
rect 6779 46560 6791 46563
rect 8021 46563 8079 46569
rect 8021 46560 8033 46563
rect 6779 46532 8033 46560
rect 6779 46529 6791 46532
rect 6733 46523 6791 46529
rect 8021 46529 8033 46532
rect 8067 46529 8079 46563
rect 8021 46523 8079 46529
rect 8110 46520 8116 46572
rect 8168 46560 8174 46572
rect 9861 46563 9919 46569
rect 9861 46560 9873 46563
rect 8168 46532 9873 46560
rect 8168 46520 8174 46532
rect 9861 46529 9873 46532
rect 9907 46529 9919 46563
rect 9861 46523 9919 46529
rect 658 46452 664 46504
rect 716 46452 722 46504
rect 1946 46492 1952 46504
rect 1907 46464 1952 46492
rect 1946 46452 1952 46464
rect 2004 46452 2010 46504
rect 4062 46452 4068 46504
rect 4120 46492 4126 46504
rect 6365 46495 6423 46501
rect 6365 46492 6377 46495
rect 4120 46464 6377 46492
rect 4120 46452 4126 46464
rect 6365 46461 6377 46464
rect 6411 46461 6423 46495
rect 6365 46455 6423 46461
rect 10042 46424 10048 46436
rect 10003 46396 10048 46424
rect 10042 46384 10048 46396
rect 10100 46384 10106 46436
rect 14 46316 20 46368
rect 72 46356 78 46368
rect 1026 46356 1032 46368
rect 72 46328 1032 46356
rect 72 46316 78 46328
rect 1026 46316 1032 46328
rect 1084 46316 1090 46368
rect 2498 46316 2504 46368
rect 2556 46356 2562 46368
rect 3421 46359 3479 46365
rect 3421 46356 3433 46359
rect 2556 46328 3433 46356
rect 2556 46316 2562 46328
rect 3421 46325 3433 46328
rect 3467 46325 3479 46359
rect 3421 46319 3479 46325
rect 4522 46316 4528 46368
rect 4580 46356 4586 46368
rect 4706 46356 4712 46368
rect 4580 46328 4712 46356
rect 4580 46316 4586 46328
rect 4706 46316 4712 46328
rect 4764 46316 4770 46368
rect 1104 46266 10856 46288
rect 1104 46214 2582 46266
rect 2634 46214 2646 46266
rect 2698 46214 2710 46266
rect 2762 46214 2774 46266
rect 2826 46214 2838 46266
rect 2890 46214 5846 46266
rect 5898 46214 5910 46266
rect 5962 46214 5974 46266
rect 6026 46214 6038 46266
rect 6090 46214 6102 46266
rect 6154 46214 9110 46266
rect 9162 46214 9174 46266
rect 9226 46214 9238 46266
rect 9290 46214 9302 46266
rect 9354 46214 9366 46266
rect 9418 46214 10856 46266
rect 1104 46192 10856 46214
rect 106 46112 112 46164
rect 164 46152 170 46164
rect 1026 46152 1032 46164
rect 164 46124 1032 46152
rect 164 46112 170 46124
rect 1026 46112 1032 46124
rect 1084 46112 1090 46164
rect 1946 46112 1952 46164
rect 2004 46152 2010 46164
rect 2409 46155 2467 46161
rect 2409 46152 2421 46155
rect 2004 46124 2421 46152
rect 2004 46112 2010 46124
rect 2409 46121 2421 46124
rect 2455 46121 2467 46155
rect 2409 46115 2467 46121
rect 4706 46112 4712 46164
rect 4764 46152 4770 46164
rect 4890 46152 4896 46164
rect 4764 46124 4896 46152
rect 4764 46112 4770 46124
rect 4890 46112 4896 46124
rect 4948 46112 4954 46164
rect 3326 46044 3332 46096
rect 3384 46084 3390 46096
rect 3510 46084 3516 46096
rect 3384 46056 3516 46084
rect 3384 46044 3390 46056
rect 3510 46044 3516 46056
rect 3568 46044 3574 46096
rect 1486 45976 1492 46028
rect 1544 46016 1550 46028
rect 1946 46016 1952 46028
rect 1544 45988 1952 46016
rect 1544 45976 1550 45988
rect 1946 45976 1952 45988
rect 2004 45976 2010 46028
rect 2958 46016 2964 46028
rect 2240 45988 2964 46016
rect 2240 45957 2268 45988
rect 2958 45976 2964 45988
rect 3016 45976 3022 46028
rect 2041 45951 2099 45957
rect 2041 45948 2053 45951
rect 1596 45920 2053 45948
rect 1596 45824 1624 45920
rect 2041 45917 2053 45920
rect 2087 45917 2099 45951
rect 2041 45911 2099 45917
rect 2225 45951 2283 45957
rect 2225 45917 2237 45951
rect 2271 45917 2283 45951
rect 2866 45948 2872 45960
rect 2827 45920 2872 45948
rect 2225 45911 2283 45917
rect 2056 45880 2084 45911
rect 2866 45908 2872 45920
rect 2924 45908 2930 45960
rect 3050 45908 3056 45960
rect 3108 45948 3114 45960
rect 3326 45948 3332 45960
rect 3108 45920 3332 45948
rect 3108 45908 3114 45920
rect 3326 45908 3332 45920
rect 3384 45908 3390 45960
rect 6914 45908 6920 45960
rect 6972 45948 6978 45960
rect 9861 45951 9919 45957
rect 9861 45948 9873 45951
rect 6972 45920 9873 45948
rect 6972 45908 6978 45920
rect 9861 45917 9873 45920
rect 9907 45917 9919 45951
rect 9861 45911 9919 45917
rect 4062 45880 4068 45892
rect 2056 45852 4068 45880
rect 4062 45840 4068 45852
rect 4120 45840 4126 45892
rect 4522 45840 4528 45892
rect 4580 45880 4586 45892
rect 4982 45880 4988 45892
rect 4580 45852 4988 45880
rect 4580 45840 4586 45852
rect 4982 45840 4988 45852
rect 5040 45840 5046 45892
rect 1578 45772 1584 45824
rect 1636 45772 1642 45824
rect 3050 45812 3056 45824
rect 3011 45784 3056 45812
rect 3050 45772 3056 45784
rect 3108 45772 3114 45824
rect 10042 45812 10048 45824
rect 10003 45784 10048 45812
rect 10042 45772 10048 45784
rect 10100 45772 10106 45824
rect 1104 45722 10856 45744
rect 1104 45670 4214 45722
rect 4266 45670 4278 45722
rect 4330 45670 4342 45722
rect 4394 45670 4406 45722
rect 4458 45670 4470 45722
rect 4522 45670 7478 45722
rect 7530 45670 7542 45722
rect 7594 45670 7606 45722
rect 7658 45670 7670 45722
rect 7722 45670 7734 45722
rect 7786 45670 10856 45722
rect 1104 45648 10856 45670
rect 2314 45608 2320 45620
rect 2275 45580 2320 45608
rect 2314 45568 2320 45580
rect 2372 45568 2378 45620
rect 3786 45500 3792 45552
rect 3844 45540 3850 45552
rect 5534 45540 5540 45552
rect 3844 45512 5540 45540
rect 3844 45500 3850 45512
rect 5534 45500 5540 45512
rect 5592 45500 5598 45552
rect 1302 45432 1308 45484
rect 1360 45472 1366 45484
rect 1397 45475 1455 45481
rect 1397 45472 1409 45475
rect 1360 45444 1409 45472
rect 1360 45432 1366 45444
rect 1397 45441 1409 45444
rect 1443 45441 1455 45475
rect 1397 45435 1455 45441
rect 2133 45475 2191 45481
rect 2133 45441 2145 45475
rect 2179 45472 2191 45475
rect 2866 45472 2872 45484
rect 2179 45444 2774 45472
rect 2827 45444 2872 45472
rect 2179 45441 2191 45444
rect 2133 45435 2191 45441
rect 2746 45404 2774 45444
rect 2866 45432 2872 45444
rect 2924 45432 2930 45484
rect 5350 45432 5356 45484
rect 5408 45472 5414 45484
rect 6549 45475 6607 45481
rect 6549 45472 6561 45475
rect 5408 45444 6561 45472
rect 5408 45432 5414 45444
rect 6549 45441 6561 45444
rect 6595 45441 6607 45475
rect 6549 45435 6607 45441
rect 4154 45404 4160 45416
rect 2746 45376 4160 45404
rect 4154 45364 4160 45376
rect 4212 45364 4218 45416
rect 2590 45296 2596 45348
rect 2648 45336 2654 45348
rect 3053 45339 3111 45345
rect 3053 45336 3065 45339
rect 2648 45308 3065 45336
rect 2648 45296 2654 45308
rect 3053 45305 3065 45308
rect 3099 45305 3111 45339
rect 3053 45299 3111 45305
rect 6365 45339 6423 45345
rect 6365 45305 6377 45339
rect 6411 45336 6423 45339
rect 6914 45336 6920 45348
rect 6411 45308 6920 45336
rect 6411 45305 6423 45308
rect 6365 45299 6423 45305
rect 6914 45296 6920 45308
rect 6972 45296 6978 45348
rect 1578 45268 1584 45280
rect 1539 45240 1584 45268
rect 1578 45228 1584 45240
rect 1636 45228 1642 45280
rect 1104 45178 10856 45200
rect 1104 45126 2582 45178
rect 2634 45126 2646 45178
rect 2698 45126 2710 45178
rect 2762 45126 2774 45178
rect 2826 45126 2838 45178
rect 2890 45126 5846 45178
rect 5898 45126 5910 45178
rect 5962 45126 5974 45178
rect 6026 45126 6038 45178
rect 6090 45126 6102 45178
rect 6154 45126 9110 45178
rect 9162 45126 9174 45178
rect 9226 45126 9238 45178
rect 9290 45126 9302 45178
rect 9354 45126 9366 45178
rect 9418 45126 10856 45178
rect 1104 45104 10856 45126
rect 5350 45064 5356 45076
rect 5311 45036 5356 45064
rect 5350 45024 5356 45036
rect 5408 45024 5414 45076
rect 6641 45067 6699 45073
rect 6641 45033 6653 45067
rect 6687 45064 6699 45067
rect 8110 45064 8116 45076
rect 6687 45036 8116 45064
rect 6687 45033 6699 45036
rect 6641 45027 6699 45033
rect 8110 45024 8116 45036
rect 8168 45024 8174 45076
rect 1486 44956 1492 45008
rect 1544 44996 1550 45008
rect 1544 44968 1624 44996
rect 1544 44956 1550 44968
rect 1486 44860 1492 44872
rect 1447 44832 1492 44860
rect 1486 44820 1492 44832
rect 1544 44820 1550 44872
rect 1596 44736 1624 44968
rect 1765 44931 1823 44937
rect 1765 44897 1777 44931
rect 1811 44928 1823 44931
rect 2314 44928 2320 44940
rect 1811 44900 2320 44928
rect 1811 44897 1823 44900
rect 1765 44891 1823 44897
rect 2314 44888 2320 44900
rect 2372 44888 2378 44940
rect 8570 44928 8576 44940
rect 3712 44900 8576 44928
rect 2777 44863 2835 44869
rect 2777 44829 2789 44863
rect 2823 44860 2835 44863
rect 3712 44860 3740 44900
rect 8570 44888 8576 44900
rect 8628 44888 8634 44940
rect 2823 44832 3740 44860
rect 5077 44863 5135 44869
rect 2823 44829 2835 44832
rect 2777 44823 2835 44829
rect 5077 44829 5089 44863
rect 5123 44829 5135 44863
rect 5077 44823 5135 44829
rect 5169 44863 5227 44869
rect 5169 44829 5181 44863
rect 5215 44829 5227 44863
rect 5169 44823 5227 44829
rect 1578 44684 1584 44736
rect 1636 44684 1642 44736
rect 2958 44724 2964 44736
rect 2919 44696 2964 44724
rect 2958 44684 2964 44696
rect 3016 44684 3022 44736
rect 5092 44724 5120 44823
rect 5184 44792 5212 44823
rect 5534 44820 5540 44872
rect 5592 44860 5598 44872
rect 5813 44863 5871 44869
rect 5813 44860 5825 44863
rect 5592 44832 5825 44860
rect 5592 44820 5598 44832
rect 5813 44829 5825 44832
rect 5859 44829 5871 44863
rect 5813 44823 5871 44829
rect 5997 44863 6055 44869
rect 5997 44829 6009 44863
rect 6043 44829 6055 44863
rect 5997 44823 6055 44829
rect 6181 44863 6239 44869
rect 6181 44829 6193 44863
rect 6227 44860 6239 44863
rect 6825 44863 6883 44869
rect 6825 44860 6837 44863
rect 6227 44832 6837 44860
rect 6227 44829 6239 44832
rect 6181 44823 6239 44829
rect 6825 44829 6837 44832
rect 6871 44829 6883 44863
rect 9858 44860 9864 44872
rect 9819 44832 9864 44860
rect 6825 44823 6883 44829
rect 6012 44792 6040 44823
rect 9858 44820 9864 44832
rect 9916 44820 9922 44872
rect 6546 44792 6552 44804
rect 5184 44764 6552 44792
rect 6546 44752 6552 44764
rect 6604 44752 6610 44804
rect 5626 44724 5632 44736
rect 5092 44696 5632 44724
rect 5626 44684 5632 44696
rect 5684 44684 5690 44736
rect 6178 44684 6184 44736
rect 6236 44724 6242 44736
rect 6638 44724 6644 44736
rect 6236 44696 6644 44724
rect 6236 44684 6242 44696
rect 6638 44684 6644 44696
rect 6696 44684 6702 44736
rect 10042 44724 10048 44736
rect 10003 44696 10048 44724
rect 10042 44684 10048 44696
rect 10100 44684 10106 44736
rect 1104 44634 10856 44656
rect 1104 44582 4214 44634
rect 4266 44582 4278 44634
rect 4330 44582 4342 44634
rect 4394 44582 4406 44634
rect 4458 44582 4470 44634
rect 4522 44582 7478 44634
rect 7530 44582 7542 44634
rect 7594 44582 7606 44634
rect 7658 44582 7670 44634
rect 7722 44582 7734 44634
rect 7786 44582 10856 44634
rect 1104 44560 10856 44582
rect 2958 44480 2964 44532
rect 3016 44520 3022 44532
rect 3326 44520 3332 44532
rect 3016 44492 3332 44520
rect 3016 44480 3022 44492
rect 3326 44480 3332 44492
rect 3384 44480 3390 44532
rect 6365 44523 6423 44529
rect 6365 44489 6377 44523
rect 6411 44520 6423 44523
rect 9858 44520 9864 44532
rect 6411 44492 9864 44520
rect 6411 44489 6423 44492
rect 6365 44483 6423 44489
rect 9858 44480 9864 44492
rect 9916 44480 9922 44532
rect 842 44344 848 44396
rect 900 44384 906 44396
rect 1673 44387 1731 44393
rect 900 44356 1164 44384
rect 900 44344 906 44356
rect 1136 44316 1164 44356
rect 1673 44353 1685 44387
rect 1719 44384 1731 44387
rect 2961 44387 3019 44393
rect 1719 44356 2912 44384
rect 1719 44353 1731 44356
rect 1673 44347 1731 44353
rect 1949 44319 2007 44325
rect 1949 44316 1961 44319
rect 1136 44288 1961 44316
rect 1949 44285 1961 44288
rect 1995 44285 2007 44319
rect 2884 44316 2912 44356
rect 2961 44353 2973 44387
rect 3007 44384 3019 44387
rect 3786 44384 3792 44396
rect 3007 44356 3792 44384
rect 3007 44353 3019 44356
rect 2961 44347 3019 44353
rect 3786 44344 3792 44356
rect 3844 44344 3850 44396
rect 6546 44384 6552 44396
rect 6507 44356 6552 44384
rect 6546 44344 6552 44356
rect 6604 44344 6610 44396
rect 9858 44384 9864 44396
rect 9819 44356 9864 44384
rect 9858 44344 9864 44356
rect 9916 44344 9922 44396
rect 3326 44316 3332 44328
rect 2884 44288 3332 44316
rect 1949 44279 2007 44285
rect 3326 44276 3332 44288
rect 3384 44276 3390 44328
rect 3142 44180 3148 44192
rect 3103 44152 3148 44180
rect 3142 44140 3148 44152
rect 3200 44140 3206 44192
rect 10042 44180 10048 44192
rect 10003 44152 10048 44180
rect 10042 44140 10048 44152
rect 10100 44140 10106 44192
rect 1104 44090 10856 44112
rect 1104 44038 2582 44090
rect 2634 44038 2646 44090
rect 2698 44038 2710 44090
rect 2762 44038 2774 44090
rect 2826 44038 2838 44090
rect 2890 44038 5846 44090
rect 5898 44038 5910 44090
rect 5962 44038 5974 44090
rect 6026 44038 6038 44090
rect 6090 44038 6102 44090
rect 6154 44038 9110 44090
rect 9162 44038 9174 44090
rect 9226 44038 9238 44090
rect 9290 44038 9302 44090
rect 9354 44038 9366 44090
rect 9418 44038 10856 44090
rect 1104 44016 10856 44038
rect 1486 43936 1492 43988
rect 1544 43976 1550 43988
rect 1857 43979 1915 43985
rect 1857 43976 1869 43979
rect 1544 43948 1869 43976
rect 1544 43936 1550 43948
rect 1857 43945 1869 43948
rect 1903 43945 1915 43979
rect 1857 43939 1915 43945
rect 2685 43979 2743 43985
rect 2685 43945 2697 43979
rect 2731 43976 2743 43979
rect 3326 43976 3332 43988
rect 2731 43948 3332 43976
rect 2731 43945 2743 43948
rect 2685 43939 2743 43945
rect 3326 43936 3332 43948
rect 3384 43936 3390 43988
rect 3786 43936 3792 43988
rect 3844 43976 3850 43988
rect 3970 43976 3976 43988
rect 3844 43948 3976 43976
rect 3844 43936 3850 43948
rect 3970 43936 3976 43948
rect 4028 43936 4034 43988
rect 4893 43979 4951 43985
rect 4893 43945 4905 43979
rect 4939 43976 4951 43979
rect 6546 43976 6552 43988
rect 4939 43948 6552 43976
rect 4939 43945 4951 43948
rect 4893 43939 4951 43945
rect 6546 43936 6552 43948
rect 6604 43936 6610 43988
rect 5626 43908 5632 43920
rect 1504 43880 5632 43908
rect 1504 43849 1532 43880
rect 5626 43868 5632 43880
rect 5684 43868 5690 43920
rect 1489 43843 1547 43849
rect 1489 43809 1501 43843
rect 1535 43809 1547 43843
rect 4525 43843 4583 43849
rect 4525 43840 4537 43843
rect 1489 43803 1547 43809
rect 1688 43812 2544 43840
rect 1688 43781 1716 43812
rect 2516 43781 2544 43812
rect 3160 43812 4537 43840
rect 3160 43784 3188 43812
rect 4525 43809 4537 43812
rect 4571 43809 4583 43843
rect 4525 43803 4583 43809
rect 1673 43775 1731 43781
rect 1673 43741 1685 43775
rect 1719 43741 1731 43775
rect 1673 43735 1731 43741
rect 2317 43775 2375 43781
rect 2317 43741 2329 43775
rect 2363 43741 2375 43775
rect 2317 43735 2375 43741
rect 2501 43775 2559 43781
rect 2501 43741 2513 43775
rect 2547 43772 2559 43775
rect 2590 43772 2596 43784
rect 2547 43744 2596 43772
rect 2547 43741 2559 43744
rect 2501 43735 2559 43741
rect 842 43664 848 43716
rect 900 43704 906 43716
rect 2332 43704 2360 43735
rect 2590 43732 2596 43744
rect 2648 43772 2654 43784
rect 3050 43772 3056 43784
rect 2648 43744 3056 43772
rect 2648 43732 2654 43744
rect 3050 43732 3056 43744
rect 3108 43732 3114 43784
rect 3142 43732 3148 43784
rect 3200 43732 3206 43784
rect 3326 43732 3332 43784
rect 3384 43772 3390 43784
rect 3789 43775 3847 43781
rect 3789 43772 3801 43775
rect 3384 43744 3801 43772
rect 3384 43732 3390 43744
rect 3789 43741 3801 43744
rect 3835 43741 3847 43775
rect 3789 43735 3847 43741
rect 4709 43775 4767 43781
rect 4709 43741 4721 43775
rect 4755 43772 4767 43775
rect 6638 43772 6644 43784
rect 4755 43744 6644 43772
rect 4755 43741 4767 43744
rect 4709 43735 4767 43741
rect 6638 43732 6644 43744
rect 6696 43732 6702 43784
rect 9861 43775 9919 43781
rect 9861 43741 9873 43775
rect 9907 43772 9919 43775
rect 9950 43772 9956 43784
rect 9907 43744 9956 43772
rect 9907 43741 9919 43744
rect 9861 43735 9919 43741
rect 9950 43732 9956 43744
rect 10008 43732 10014 43784
rect 5534 43704 5540 43716
rect 900 43676 5540 43704
rect 900 43664 906 43676
rect 5534 43664 5540 43676
rect 5592 43664 5598 43716
rect 3970 43636 3976 43648
rect 3931 43608 3976 43636
rect 3970 43596 3976 43608
rect 4028 43596 4034 43648
rect 10042 43636 10048 43648
rect 10003 43608 10048 43636
rect 10042 43596 10048 43608
rect 10100 43596 10106 43648
rect 1104 43546 10856 43568
rect 1104 43494 4214 43546
rect 4266 43494 4278 43546
rect 4330 43494 4342 43546
rect 4394 43494 4406 43546
rect 4458 43494 4470 43546
rect 4522 43494 7478 43546
rect 7530 43494 7542 43546
rect 7594 43494 7606 43546
rect 7658 43494 7670 43546
rect 7722 43494 7734 43546
rect 7786 43494 10856 43546
rect 1104 43472 10856 43494
rect 934 43392 940 43444
rect 992 43432 998 43444
rect 992 43404 1716 43432
rect 992 43392 998 43404
rect 1688 43296 1716 43404
rect 3142 43392 3148 43444
rect 3200 43392 3206 43444
rect 3326 43432 3332 43444
rect 3287 43404 3332 43432
rect 3326 43392 3332 43404
rect 3384 43392 3390 43444
rect 6362 43392 6368 43444
rect 6420 43432 6426 43444
rect 6914 43432 6920 43444
rect 6420 43404 6920 43432
rect 6420 43392 6426 43404
rect 6914 43392 6920 43404
rect 6972 43392 6978 43444
rect 9950 43432 9956 43444
rect 9911 43404 9956 43432
rect 9950 43392 9956 43404
rect 10008 43392 10014 43444
rect 1762 43324 1768 43376
rect 1820 43364 1826 43376
rect 3053 43367 3111 43373
rect 3053 43364 3065 43367
rect 1820 43336 3065 43364
rect 1820 43324 1826 43336
rect 3053 43333 3065 43336
rect 3099 43333 3111 43367
rect 3160 43364 3188 43392
rect 3160 43336 3372 43364
rect 3053 43327 3111 43333
rect 3344 43308 3372 43336
rect 2777 43299 2835 43305
rect 1688 43268 1808 43296
rect 1486 43228 1492 43240
rect 1447 43200 1492 43228
rect 1486 43188 1492 43200
rect 1544 43188 1550 43240
rect 1780 43237 1808 43268
rect 2777 43265 2789 43299
rect 2823 43265 2835 43299
rect 2958 43296 2964 43308
rect 2919 43268 2964 43296
rect 2777 43259 2835 43265
rect 1765 43231 1823 43237
rect 1765 43197 1777 43231
rect 1811 43197 1823 43231
rect 2792 43228 2820 43259
rect 2958 43256 2964 43268
rect 3016 43256 3022 43308
rect 3142 43296 3148 43308
rect 3103 43268 3148 43296
rect 3142 43256 3148 43268
rect 3200 43256 3206 43308
rect 3326 43256 3332 43308
rect 3384 43256 3390 43308
rect 3694 43256 3700 43308
rect 3752 43296 3758 43308
rect 3789 43299 3847 43305
rect 3789 43296 3801 43299
rect 3752 43268 3801 43296
rect 3752 43256 3758 43268
rect 3789 43265 3801 43268
rect 3835 43265 3847 43299
rect 3789 43259 3847 43265
rect 9674 43256 9680 43308
rect 9732 43296 9738 43308
rect 10137 43299 10195 43305
rect 10137 43296 10149 43299
rect 9732 43268 10149 43296
rect 9732 43256 9738 43268
rect 10137 43265 10149 43268
rect 10183 43265 10195 43299
rect 10137 43259 10195 43265
rect 9766 43228 9772 43240
rect 2792 43200 9772 43228
rect 1765 43191 1823 43197
rect 9766 43188 9772 43200
rect 9824 43188 9830 43240
rect 842 43120 848 43172
rect 900 43160 906 43172
rect 2590 43160 2596 43172
rect 900 43132 2596 43160
rect 900 43120 906 43132
rect 2590 43120 2596 43132
rect 2648 43120 2654 43172
rect 3602 43120 3608 43172
rect 3660 43160 3666 43172
rect 3970 43160 3976 43172
rect 3660 43132 3832 43160
rect 3931 43132 3976 43160
rect 3660 43120 3666 43132
rect 3804 43104 3832 43132
rect 3970 43120 3976 43132
rect 4028 43120 4034 43172
rect 3786 43052 3792 43104
rect 3844 43052 3850 43104
rect 1104 43002 10856 43024
rect 1104 42950 2582 43002
rect 2634 42950 2646 43002
rect 2698 42950 2710 43002
rect 2762 42950 2774 43002
rect 2826 42950 2838 43002
rect 2890 42950 5846 43002
rect 5898 42950 5910 43002
rect 5962 42950 5974 43002
rect 6026 42950 6038 43002
rect 6090 42950 6102 43002
rect 6154 42950 9110 43002
rect 9162 42950 9174 43002
rect 9226 42950 9238 43002
rect 9290 42950 9302 43002
rect 9354 42950 9366 43002
rect 9418 42950 10856 43002
rect 1104 42928 10856 42950
rect 1486 42848 1492 42900
rect 1544 42888 1550 42900
rect 2133 42891 2191 42897
rect 2133 42888 2145 42891
rect 1544 42860 2145 42888
rect 1544 42848 1550 42860
rect 2133 42857 2145 42860
rect 2179 42857 2191 42891
rect 3326 42888 3332 42900
rect 2133 42851 2191 42857
rect 2608 42860 3332 42888
rect 1765 42755 1823 42761
rect 1765 42721 1777 42755
rect 1811 42752 1823 42755
rect 2608 42752 2636 42860
rect 3326 42848 3332 42860
rect 3384 42848 3390 42900
rect 1811 42724 2636 42752
rect 1811 42721 1823 42724
rect 1765 42715 1823 42721
rect 6270 42712 6276 42764
rect 6328 42752 6334 42764
rect 8386 42752 8392 42764
rect 6328 42724 8392 42752
rect 6328 42712 6334 42724
rect 8386 42712 8392 42724
rect 8444 42712 8450 42764
rect 842 42644 848 42696
rect 900 42684 906 42696
rect 1949 42687 2007 42693
rect 1949 42684 1961 42687
rect 900 42656 1961 42684
rect 900 42644 906 42656
rect 1949 42653 1961 42656
rect 1995 42653 2007 42687
rect 2593 42687 2651 42693
rect 2593 42684 2605 42687
rect 1949 42647 2007 42653
rect 2056 42656 2605 42684
rect 1670 42576 1676 42628
rect 1728 42616 1734 42628
rect 2056 42616 2084 42656
rect 2593 42653 2605 42656
rect 2639 42653 2651 42687
rect 2593 42647 2651 42653
rect 3142 42644 3148 42696
rect 3200 42684 3206 42696
rect 3510 42684 3516 42696
rect 3200 42656 3516 42684
rect 3200 42644 3206 42656
rect 3510 42644 3516 42656
rect 3568 42644 3574 42696
rect 3789 42687 3847 42693
rect 3789 42653 3801 42687
rect 3835 42684 3847 42687
rect 4154 42684 4160 42696
rect 3835 42656 4160 42684
rect 3835 42653 3847 42656
rect 3789 42647 3847 42653
rect 4154 42644 4160 42656
rect 4212 42644 4218 42696
rect 6454 42684 6460 42696
rect 6415 42656 6460 42684
rect 6454 42644 6460 42656
rect 6512 42644 6518 42696
rect 9861 42687 9919 42693
rect 9861 42653 9873 42687
rect 9907 42684 9919 42687
rect 9950 42684 9956 42696
rect 9907 42656 9956 42684
rect 9907 42653 9919 42656
rect 9861 42647 9919 42653
rect 9950 42644 9956 42656
rect 10008 42644 10014 42696
rect 1728 42588 2084 42616
rect 1728 42576 1734 42588
rect 2774 42508 2780 42560
rect 2832 42548 2838 42560
rect 3970 42548 3976 42560
rect 2832 42520 2877 42548
rect 3931 42520 3976 42548
rect 2832 42508 2838 42520
rect 3970 42508 3976 42520
rect 4028 42508 4034 42560
rect 6273 42551 6331 42557
rect 6273 42517 6285 42551
rect 6319 42548 6331 42551
rect 9858 42548 9864 42560
rect 6319 42520 9864 42548
rect 6319 42517 6331 42520
rect 6273 42511 6331 42517
rect 9858 42508 9864 42520
rect 9916 42508 9922 42560
rect 10042 42548 10048 42560
rect 10003 42520 10048 42548
rect 10042 42508 10048 42520
rect 10100 42508 10106 42560
rect 1104 42458 10856 42480
rect 1104 42406 4214 42458
rect 4266 42406 4278 42458
rect 4330 42406 4342 42458
rect 4394 42406 4406 42458
rect 4458 42406 4470 42458
rect 4522 42406 7478 42458
rect 7530 42406 7542 42458
rect 7594 42406 7606 42458
rect 7658 42406 7670 42458
rect 7722 42406 7734 42458
rect 7786 42406 10856 42458
rect 1104 42384 10856 42406
rect 3326 42304 3332 42356
rect 3384 42344 3390 42356
rect 3970 42344 3976 42356
rect 3384 42316 3976 42344
rect 3384 42304 3390 42316
rect 3970 42304 3976 42316
rect 4028 42304 4034 42356
rect 4430 42236 4436 42288
rect 4488 42276 4494 42288
rect 4798 42276 4804 42288
rect 4488 42248 4804 42276
rect 4488 42236 4494 42248
rect 4798 42236 4804 42248
rect 4856 42236 4862 42288
rect 1397 42211 1455 42217
rect 1397 42177 1409 42211
rect 1443 42208 1455 42211
rect 1762 42208 1768 42220
rect 1443 42180 1768 42208
rect 1443 42177 1455 42180
rect 1397 42171 1455 42177
rect 1762 42168 1768 42180
rect 1820 42168 1826 42220
rect 2130 42208 2136 42220
rect 2091 42180 2136 42208
rect 2130 42168 2136 42180
rect 2188 42168 2194 42220
rect 2866 42208 2872 42220
rect 2827 42180 2872 42208
rect 2866 42168 2872 42180
rect 2924 42168 2930 42220
rect 9490 42168 9496 42220
rect 9548 42208 9554 42220
rect 9861 42211 9919 42217
rect 9861 42208 9873 42211
rect 9548 42180 9873 42208
rect 9548 42168 9554 42180
rect 9861 42177 9873 42180
rect 9907 42177 9919 42211
rect 9861 42171 9919 42177
rect 2314 42140 2320 42152
rect 2148 42112 2320 42140
rect 2148 42084 2176 42112
rect 2314 42100 2320 42112
rect 2372 42100 2378 42152
rect 2130 42032 2136 42084
rect 2188 42032 2194 42084
rect 1578 42004 1584 42016
rect 1539 41976 1584 42004
rect 1578 41964 1584 41976
rect 1636 41964 1642 42016
rect 2314 42004 2320 42016
rect 2275 41976 2320 42004
rect 2314 41964 2320 41976
rect 2372 41964 2378 42016
rect 3050 42004 3056 42016
rect 3011 41976 3056 42004
rect 3050 41964 3056 41976
rect 3108 41964 3114 42016
rect 10042 42004 10048 42016
rect 10003 41976 10048 42004
rect 10042 41964 10048 41976
rect 10100 41964 10106 42016
rect 1104 41914 10856 41936
rect 1104 41862 2582 41914
rect 2634 41862 2646 41914
rect 2698 41862 2710 41914
rect 2762 41862 2774 41914
rect 2826 41862 2838 41914
rect 2890 41862 5846 41914
rect 5898 41862 5910 41914
rect 5962 41862 5974 41914
rect 6026 41862 6038 41914
rect 6090 41862 6102 41914
rect 6154 41862 9110 41914
rect 9162 41862 9174 41914
rect 9226 41862 9238 41914
rect 9290 41862 9302 41914
rect 9354 41862 9366 41914
rect 9418 41862 10856 41914
rect 1104 41840 10856 41862
rect 658 41760 664 41812
rect 716 41800 722 41812
rect 2639 41803 2697 41809
rect 2639 41800 2651 41803
rect 716 41772 2651 41800
rect 716 41760 722 41772
rect 2639 41769 2651 41772
rect 2685 41769 2697 41803
rect 2639 41763 2697 41769
rect 5077 41803 5135 41809
rect 5077 41769 5089 41803
rect 5123 41800 5135 41803
rect 9674 41800 9680 41812
rect 5123 41772 9680 41800
rect 5123 41769 5135 41772
rect 5077 41763 5135 41769
rect 9674 41760 9680 41772
rect 9732 41760 9738 41812
rect 9950 41800 9956 41812
rect 9911 41772 9956 41800
rect 9950 41760 9956 41772
rect 10008 41760 10014 41812
rect 1949 41735 2007 41741
rect 1949 41701 1961 41735
rect 1995 41732 2007 41735
rect 6362 41732 6368 41744
rect 1995 41704 6368 41732
rect 1995 41701 2007 41704
rect 1949 41695 2007 41701
rect 6362 41692 6368 41704
rect 6420 41692 6426 41744
rect 658 41624 664 41676
rect 716 41664 722 41676
rect 1394 41664 1400 41676
rect 716 41636 1400 41664
rect 716 41624 722 41636
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 2314 41624 2320 41676
rect 2372 41624 2378 41676
rect 2409 41667 2467 41673
rect 2409 41633 2421 41667
rect 2455 41664 2467 41667
rect 2866 41664 2872 41676
rect 2455 41636 2872 41664
rect 2455 41633 2467 41636
rect 2409 41627 2467 41633
rect 2866 41624 2872 41636
rect 2924 41624 2930 41676
rect 3694 41664 3700 41676
rect 2976 41636 3700 41664
rect 842 41488 848 41540
rect 900 41528 906 41540
rect 1394 41528 1400 41540
rect 900 41500 1400 41528
rect 900 41488 906 41500
rect 1394 41488 1400 41500
rect 1452 41488 1458 41540
rect 1762 41528 1768 41540
rect 1723 41500 1768 41528
rect 1762 41488 1768 41500
rect 1820 41488 1826 41540
rect 2332 41472 2360 41624
rect 2682 41556 2688 41608
rect 2740 41596 2746 41608
rect 2976 41596 3004 41636
rect 3694 41624 3700 41636
rect 3752 41624 3758 41676
rect 5258 41624 5264 41676
rect 5316 41664 5322 41676
rect 5316 41636 6408 41664
rect 5316 41624 5322 41636
rect 6380 41608 6408 41636
rect 2740 41568 3004 41596
rect 2740 41556 2746 41568
rect 3050 41556 3056 41608
rect 3108 41596 3114 41608
rect 4709 41599 4767 41605
rect 4709 41596 4721 41599
rect 3108 41568 4721 41596
rect 3108 41556 3114 41568
rect 4709 41565 4721 41568
rect 4755 41565 4767 41599
rect 4709 41559 4767 41565
rect 4893 41599 4951 41605
rect 4893 41565 4905 41599
rect 4939 41565 4951 41599
rect 4893 41559 4951 41565
rect 4908 41528 4936 41559
rect 5442 41556 5448 41608
rect 5500 41596 5506 41608
rect 5902 41596 5908 41608
rect 5500 41568 5908 41596
rect 5500 41556 5506 41568
rect 5902 41556 5908 41568
rect 5960 41556 5966 41608
rect 6362 41556 6368 41608
rect 6420 41556 6426 41608
rect 9766 41556 9772 41608
rect 9824 41596 9830 41608
rect 10137 41599 10195 41605
rect 10137 41596 10149 41599
rect 9824 41568 10149 41596
rect 9824 41556 9830 41568
rect 10137 41565 10149 41568
rect 10183 41565 10195 41599
rect 10137 41559 10195 41565
rect 5810 41528 5816 41540
rect 4908 41500 5816 41528
rect 5810 41488 5816 41500
rect 5868 41528 5874 41540
rect 6638 41528 6644 41540
rect 5868 41500 6644 41528
rect 5868 41488 5874 41500
rect 6638 41488 6644 41500
rect 6696 41488 6702 41540
rect 2314 41420 2320 41472
rect 2372 41420 2378 41472
rect 5074 41420 5080 41472
rect 5132 41460 5138 41472
rect 7006 41460 7012 41472
rect 5132 41432 7012 41460
rect 5132 41420 5138 41432
rect 7006 41420 7012 41432
rect 7064 41420 7070 41472
rect 1104 41370 10856 41392
rect 1104 41318 4214 41370
rect 4266 41318 4278 41370
rect 4330 41318 4342 41370
rect 4394 41318 4406 41370
rect 4458 41318 4470 41370
rect 4522 41318 7478 41370
rect 7530 41318 7542 41370
rect 7594 41318 7606 41370
rect 7658 41318 7670 41370
rect 7722 41318 7734 41370
rect 7786 41318 10856 41370
rect 1104 41296 10856 41318
rect 750 41216 756 41268
rect 808 41256 814 41268
rect 1486 41256 1492 41268
rect 808 41228 1492 41256
rect 808 41216 814 41228
rect 1486 41216 1492 41228
rect 1544 41216 1550 41268
rect 1762 41216 1768 41268
rect 1820 41256 1826 41268
rect 1949 41259 2007 41265
rect 1949 41256 1961 41259
rect 1820 41228 1961 41256
rect 1820 41216 1826 41228
rect 1949 41225 1961 41228
rect 1995 41225 2007 41259
rect 1949 41219 2007 41225
rect 2682 41216 2688 41268
rect 2740 41216 2746 41268
rect 2866 41256 2872 41268
rect 2827 41228 2872 41256
rect 2866 41216 2872 41228
rect 2924 41216 2930 41268
rect 5353 41259 5411 41265
rect 5353 41225 5365 41259
rect 5399 41256 5411 41259
rect 6454 41256 6460 41268
rect 5399 41228 6460 41256
rect 5399 41225 5411 41228
rect 5353 41219 5411 41225
rect 6454 41216 6460 41228
rect 6512 41216 6518 41268
rect 2700 41188 2728 41216
rect 3510 41188 3516 41200
rect 2700 41160 3516 41188
rect 3510 41148 3516 41160
rect 3568 41148 3574 41200
rect 5534 41148 5540 41200
rect 5592 41188 5598 41200
rect 6914 41188 6920 41200
rect 5592 41160 6920 41188
rect 5592 41148 5598 41160
rect 6914 41148 6920 41160
rect 6972 41148 6978 41200
rect 1394 41080 1400 41132
rect 1452 41120 1458 41132
rect 1765 41123 1823 41129
rect 1765 41120 1777 41123
rect 1452 41092 1777 41120
rect 1452 41080 1458 41092
rect 1765 41089 1777 41092
rect 1811 41120 1823 41123
rect 2685 41123 2743 41129
rect 2685 41120 2697 41123
rect 1811 41092 2697 41120
rect 1811 41089 1823 41092
rect 1765 41083 1823 41089
rect 2685 41089 2697 41092
rect 2731 41089 2743 41123
rect 2685 41083 2743 41089
rect 2774 41080 2780 41132
rect 2832 41120 2838 41132
rect 3329 41123 3387 41129
rect 3329 41120 3341 41123
rect 2832 41092 3341 41120
rect 2832 41080 2838 41092
rect 3329 41089 3341 41092
rect 3375 41089 3387 41123
rect 3329 41083 3387 41089
rect 5169 41123 5227 41129
rect 5169 41089 5181 41123
rect 5215 41089 5227 41123
rect 5169 41083 5227 41089
rect 1581 41055 1639 41061
rect 1581 41021 1593 41055
rect 1627 41021 1639 41055
rect 1581 41015 1639 41021
rect 2501 41055 2559 41061
rect 2501 41021 2513 41055
rect 2547 41052 2559 41055
rect 3050 41052 3056 41064
rect 2547 41024 3056 41052
rect 2547 41021 2559 41024
rect 2501 41015 2559 41021
rect 1596 40916 1624 41015
rect 3050 41012 3056 41024
rect 3108 41012 3114 41064
rect 4430 41012 4436 41064
rect 4488 41052 4494 41064
rect 4985 41055 5043 41061
rect 4985 41052 4997 41055
rect 4488 41024 4997 41052
rect 4488 41012 4494 41024
rect 4985 41021 4997 41024
rect 5031 41021 5043 41055
rect 5184 41052 5212 41083
rect 5626 41080 5632 41132
rect 5684 41120 5690 41132
rect 5902 41120 5908 41132
rect 5684 41092 5908 41120
rect 5684 41080 5690 41092
rect 5902 41080 5908 41092
rect 5960 41080 5966 41132
rect 7006 41080 7012 41132
rect 7064 41120 7070 41132
rect 9861 41123 9919 41129
rect 9861 41120 9873 41123
rect 7064 41092 9873 41120
rect 7064 41080 7070 41092
rect 9861 41089 9873 41092
rect 9907 41089 9919 41123
rect 9861 41083 9919 41089
rect 5810 41052 5816 41064
rect 5184 41024 5816 41052
rect 4985 41015 5043 41021
rect 5810 41012 5816 41024
rect 5868 41052 5874 41064
rect 6454 41052 6460 41064
rect 5868 41024 6460 41052
rect 5868 41012 5874 41024
rect 6454 41012 6460 41024
rect 6512 41012 6518 41064
rect 2774 40944 2780 40996
rect 2832 40984 2838 40996
rect 3513 40987 3571 40993
rect 3513 40984 3525 40987
rect 2832 40956 3525 40984
rect 2832 40944 2838 40956
rect 3513 40953 3525 40956
rect 3559 40953 3571 40987
rect 10042 40984 10048 40996
rect 10003 40956 10048 40984
rect 3513 40947 3571 40953
rect 10042 40944 10048 40956
rect 10100 40944 10106 40996
rect 3050 40916 3056 40928
rect 1596 40888 3056 40916
rect 3050 40876 3056 40888
rect 3108 40876 3114 40928
rect 4982 40876 4988 40928
rect 5040 40916 5046 40928
rect 5442 40916 5448 40928
rect 5040 40888 5448 40916
rect 5040 40876 5046 40888
rect 5442 40876 5448 40888
rect 5500 40876 5506 40928
rect 1104 40826 10856 40848
rect 1104 40774 2582 40826
rect 2634 40774 2646 40826
rect 2698 40774 2710 40826
rect 2762 40774 2774 40826
rect 2826 40774 2838 40826
rect 2890 40774 5846 40826
rect 5898 40774 5910 40826
rect 5962 40774 5974 40826
rect 6026 40774 6038 40826
rect 6090 40774 6102 40826
rect 6154 40774 9110 40826
rect 9162 40774 9174 40826
rect 9226 40774 9238 40826
rect 9290 40774 9302 40826
rect 9354 40774 9366 40826
rect 9418 40774 10856 40826
rect 1104 40752 10856 40774
rect 1026 40672 1032 40724
rect 1084 40712 1090 40724
rect 9217 40715 9275 40721
rect 1084 40684 2452 40712
rect 1084 40672 1090 40684
rect 2130 40644 2136 40656
rect 1412 40616 2136 40644
rect 1412 40517 1440 40616
rect 2130 40604 2136 40616
rect 2188 40604 2194 40656
rect 2424 40585 2452 40684
rect 9217 40681 9229 40715
rect 9263 40712 9275 40715
rect 9490 40712 9496 40724
rect 9263 40684 9496 40712
rect 9263 40681 9275 40684
rect 9217 40675 9275 40681
rect 9490 40672 9496 40684
rect 9548 40672 9554 40724
rect 2866 40604 2872 40656
rect 2924 40644 2930 40656
rect 4430 40644 4436 40656
rect 2924 40616 4436 40644
rect 2924 40604 2930 40616
rect 4430 40604 4436 40616
rect 4488 40604 4494 40656
rect 4982 40604 4988 40656
rect 5040 40644 5046 40656
rect 5350 40644 5356 40656
rect 5040 40616 5356 40644
rect 5040 40604 5046 40616
rect 5350 40604 5356 40616
rect 5408 40604 5414 40656
rect 2409 40579 2467 40585
rect 2409 40545 2421 40579
rect 2455 40545 2467 40579
rect 2409 40539 2467 40545
rect 3878 40536 3884 40588
rect 3936 40536 3942 40588
rect 1397 40511 1455 40517
rect 1397 40477 1409 40511
rect 1443 40477 1455 40511
rect 2130 40508 2136 40520
rect 2091 40480 2136 40508
rect 1397 40471 1455 40477
rect 2130 40468 2136 40480
rect 2188 40468 2194 40520
rect 3789 40511 3847 40517
rect 3789 40477 3801 40511
rect 3835 40508 3847 40511
rect 3896 40508 3924 40536
rect 3835 40480 3924 40508
rect 3835 40477 3847 40480
rect 3789 40471 3847 40477
rect 5350 40468 5356 40520
rect 5408 40508 5414 40520
rect 9401 40511 9459 40517
rect 9401 40508 9413 40511
rect 5408 40480 9413 40508
rect 5408 40468 5414 40480
rect 9401 40477 9413 40480
rect 9447 40477 9459 40511
rect 9858 40508 9864 40520
rect 9819 40480 9864 40508
rect 9401 40471 9459 40477
rect 9858 40468 9864 40480
rect 9916 40468 9922 40520
rect 106 40400 112 40452
rect 164 40440 170 40452
rect 1762 40440 1768 40452
rect 164 40412 1768 40440
rect 164 40400 170 40412
rect 1762 40400 1768 40412
rect 1820 40400 1826 40452
rect 1578 40372 1584 40384
rect 1539 40344 1584 40372
rect 1578 40332 1584 40344
rect 1636 40332 1642 40384
rect 3970 40372 3976 40384
rect 3931 40344 3976 40372
rect 3970 40332 3976 40344
rect 4028 40332 4034 40384
rect 10042 40372 10048 40384
rect 10003 40344 10048 40372
rect 10042 40332 10048 40344
rect 10100 40332 10106 40384
rect 1104 40282 10856 40304
rect 1104 40230 4214 40282
rect 4266 40230 4278 40282
rect 4330 40230 4342 40282
rect 4394 40230 4406 40282
rect 4458 40230 4470 40282
rect 4522 40230 7478 40282
rect 7530 40230 7542 40282
rect 7594 40230 7606 40282
rect 7658 40230 7670 40282
rect 7722 40230 7734 40282
rect 7786 40230 10856 40282
rect 1104 40208 10856 40230
rect 2130 40128 2136 40180
rect 2188 40168 2194 40180
rect 2409 40171 2467 40177
rect 2409 40168 2421 40171
rect 2188 40140 2421 40168
rect 2188 40128 2194 40140
rect 2409 40137 2421 40140
rect 2455 40137 2467 40171
rect 2409 40131 2467 40137
rect 9217 40171 9275 40177
rect 9217 40137 9229 40171
rect 9263 40168 9275 40171
rect 9858 40168 9864 40180
rect 9263 40140 9864 40168
rect 9263 40137 9275 40140
rect 9217 40131 9275 40137
rect 9858 40128 9864 40140
rect 9916 40128 9922 40180
rect 658 40060 664 40112
rect 716 40100 722 40112
rect 716 40072 2452 40100
rect 716 40060 722 40072
rect 2424 40044 2452 40072
rect 2958 40060 2964 40112
rect 3016 40100 3022 40112
rect 3145 40103 3203 40109
rect 3145 40100 3157 40103
rect 3016 40072 3157 40100
rect 3016 40060 3022 40072
rect 3145 40069 3157 40072
rect 3191 40069 3203 40103
rect 3145 40063 3203 40069
rect 5442 40060 5448 40112
rect 5500 40060 5506 40112
rect 6914 40060 6920 40112
rect 6972 40100 6978 40112
rect 6972 40072 9444 40100
rect 6972 40060 6978 40072
rect 1026 39992 1032 40044
rect 1084 40032 1090 40044
rect 1394 40032 1400 40044
rect 1084 40004 1400 40032
rect 1084 39992 1090 40004
rect 1394 39992 1400 40004
rect 1452 40032 1458 40044
rect 2225 40035 2283 40041
rect 2225 40032 2237 40035
rect 1452 40004 2237 40032
rect 1452 39992 1458 40004
rect 2225 40001 2237 40004
rect 2271 40001 2283 40035
rect 2225 39995 2283 40001
rect 2406 39992 2412 40044
rect 2464 39992 2470 40044
rect 2498 39992 2504 40044
rect 2556 40032 2562 40044
rect 2774 40032 2780 40044
rect 2556 40004 2780 40032
rect 2556 39992 2562 40004
rect 2774 39992 2780 40004
rect 2832 40032 2838 40044
rect 2869 40035 2927 40041
rect 2869 40032 2881 40035
rect 2832 40004 2881 40032
rect 2832 39992 2838 40004
rect 2869 40001 2881 40004
rect 2915 40001 2927 40035
rect 2869 39995 2927 40001
rect 3789 40035 3847 40041
rect 3789 40001 3801 40035
rect 3835 40032 3847 40035
rect 5460 40032 5488 40060
rect 9416 40041 9444 40072
rect 3835 40004 5488 40032
rect 9401 40035 9459 40041
rect 3835 40001 3847 40004
rect 3789 39995 3847 40001
rect 9401 40001 9413 40035
rect 9447 40001 9459 40035
rect 9858 40032 9864 40044
rect 9819 40004 9864 40032
rect 9401 39995 9459 40001
rect 9858 39992 9864 40004
rect 9916 39992 9922 40044
rect 2041 39967 2099 39973
rect 2041 39933 2053 39967
rect 2087 39964 2099 39967
rect 2087 39936 2774 39964
rect 2087 39933 2099 39936
rect 2041 39927 2099 39933
rect 2746 39896 2774 39936
rect 5442 39924 5448 39976
rect 5500 39964 5506 39976
rect 5626 39964 5632 39976
rect 5500 39936 5632 39964
rect 5500 39924 5506 39936
rect 5626 39924 5632 39936
rect 5684 39924 5690 39976
rect 2866 39896 2872 39908
rect 2746 39868 2872 39896
rect 2866 39856 2872 39868
rect 2924 39856 2930 39908
rect 3970 39828 3976 39840
rect 3931 39800 3976 39828
rect 3970 39788 3976 39800
rect 4028 39788 4034 39840
rect 10042 39828 10048 39840
rect 10003 39800 10048 39828
rect 10042 39788 10048 39800
rect 10100 39788 10106 39840
rect 1104 39738 10856 39760
rect 1104 39686 2582 39738
rect 2634 39686 2646 39738
rect 2698 39686 2710 39738
rect 2762 39686 2774 39738
rect 2826 39686 2838 39738
rect 2890 39686 5846 39738
rect 5898 39686 5910 39738
rect 5962 39686 5974 39738
rect 6026 39686 6038 39738
rect 6090 39686 6102 39738
rect 6154 39686 9110 39738
rect 9162 39686 9174 39738
rect 9226 39686 9238 39738
rect 9290 39686 9302 39738
rect 9354 39686 9366 39738
rect 9418 39686 10856 39738
rect 1104 39664 10856 39686
rect 5629 39627 5687 39633
rect 5629 39593 5641 39627
rect 5675 39624 5687 39627
rect 6914 39624 6920 39636
rect 5675 39596 6920 39624
rect 5675 39593 5687 39596
rect 5629 39587 5687 39593
rect 6914 39584 6920 39596
rect 6972 39584 6978 39636
rect 9858 39624 9864 39636
rect 9819 39596 9864 39624
rect 9858 39584 9864 39596
rect 9916 39584 9922 39636
rect 3145 39559 3203 39565
rect 3145 39525 3157 39559
rect 3191 39556 3203 39559
rect 6362 39556 6368 39568
rect 3191 39528 6368 39556
rect 3191 39525 3203 39528
rect 3145 39519 3203 39525
rect 6362 39516 6368 39528
rect 6420 39516 6426 39568
rect 6641 39559 6699 39565
rect 6641 39525 6653 39559
rect 6687 39556 6699 39559
rect 7006 39556 7012 39568
rect 6687 39528 7012 39556
rect 6687 39525 6699 39528
rect 6641 39519 6699 39525
rect 7006 39516 7012 39528
rect 7064 39516 7070 39568
rect 3050 39488 3056 39500
rect 2884 39460 3056 39488
rect 2884 39432 2912 39460
rect 3050 39448 3056 39460
rect 3108 39448 3114 39500
rect 106 39380 112 39432
rect 164 39420 170 39432
rect 1397 39423 1455 39429
rect 1397 39420 1409 39423
rect 164 39392 1409 39420
rect 164 39380 170 39392
rect 1397 39389 1409 39392
rect 1443 39389 1455 39423
rect 1397 39383 1455 39389
rect 2498 39380 2504 39432
rect 2556 39380 2562 39432
rect 2866 39420 2872 39432
rect 2827 39392 2872 39420
rect 2866 39380 2872 39392
rect 2924 39380 2930 39432
rect 2961 39423 3019 39429
rect 2961 39389 2973 39423
rect 3007 39389 3019 39423
rect 2961 39383 3019 39389
rect 3789 39423 3847 39429
rect 3789 39389 3801 39423
rect 3835 39420 3847 39423
rect 4062 39420 4068 39432
rect 3835 39392 4068 39420
rect 3835 39389 3847 39392
rect 3789 39383 3847 39389
rect 2516 39352 2544 39380
rect 2774 39352 2780 39364
rect 2516 39324 2780 39352
rect 2774 39312 2780 39324
rect 2832 39352 2838 39364
rect 2976 39352 3004 39383
rect 4062 39380 4068 39392
rect 4120 39380 4126 39432
rect 5261 39423 5319 39429
rect 5261 39389 5273 39423
rect 5307 39389 5319 39423
rect 5261 39383 5319 39389
rect 5445 39423 5503 39429
rect 5445 39389 5457 39423
rect 5491 39420 5503 39423
rect 5626 39420 5632 39432
rect 5491 39392 5632 39420
rect 5491 39389 5503 39392
rect 5445 39383 5503 39389
rect 2832 39324 3004 39352
rect 2832 39312 2838 39324
rect 3050 39312 3056 39364
rect 3108 39352 3114 39364
rect 5276 39352 5304 39383
rect 5626 39380 5632 39392
rect 5684 39380 5690 39432
rect 6730 39380 6736 39432
rect 6788 39420 6794 39432
rect 6825 39423 6883 39429
rect 6825 39420 6837 39423
rect 6788 39392 6837 39420
rect 6788 39380 6794 39392
rect 6825 39389 6837 39392
rect 6871 39389 6883 39423
rect 6825 39383 6883 39389
rect 8754 39380 8760 39432
rect 8812 39420 8818 39432
rect 10045 39423 10103 39429
rect 10045 39420 10057 39423
rect 8812 39392 10057 39420
rect 8812 39380 8818 39392
rect 10045 39389 10057 39392
rect 10091 39389 10103 39423
rect 10045 39383 10103 39389
rect 3108 39324 5304 39352
rect 3108 39312 3114 39324
rect 1394 39244 1400 39296
rect 1452 39284 1458 39296
rect 1581 39287 1639 39293
rect 1581 39284 1593 39287
rect 1452 39256 1593 39284
rect 1452 39244 1458 39256
rect 1581 39253 1593 39256
rect 1627 39253 1639 39287
rect 3970 39284 3976 39296
rect 3931 39256 3976 39284
rect 1581 39247 1639 39253
rect 3970 39244 3976 39256
rect 4028 39244 4034 39296
rect 1104 39194 10856 39216
rect 1104 39142 4214 39194
rect 4266 39142 4278 39194
rect 4330 39142 4342 39194
rect 4394 39142 4406 39194
rect 4458 39142 4470 39194
rect 4522 39142 7478 39194
rect 7530 39142 7542 39194
rect 7594 39142 7606 39194
rect 7658 39142 7670 39194
rect 7722 39142 7734 39194
rect 7786 39142 10856 39194
rect 1104 39120 10856 39142
rect 1026 39040 1032 39092
rect 1084 39080 1090 39092
rect 2406 39080 2412 39092
rect 1084 39052 2412 39080
rect 1084 39040 1090 39052
rect 2406 39040 2412 39052
rect 2464 39040 2470 39092
rect 6730 39080 6736 39092
rect 6691 39052 6736 39080
rect 6730 39040 6736 39052
rect 6788 39040 6794 39092
rect 3694 39012 3700 39024
rect 2792 38984 3700 39012
rect 474 38904 480 38956
rect 532 38944 538 38956
rect 2792 38953 2820 38984
rect 3694 38972 3700 38984
rect 3752 38972 3758 39024
rect 4430 38972 4436 39024
rect 4488 39012 4494 39024
rect 5626 39012 5632 39024
rect 4488 38984 5632 39012
rect 4488 38972 4494 38984
rect 5626 38972 5632 38984
rect 5684 38972 5690 39024
rect 1765 38947 1823 38953
rect 1765 38944 1777 38947
rect 532 38916 1777 38944
rect 532 38904 538 38916
rect 1765 38913 1777 38916
rect 1811 38913 1823 38947
rect 1765 38907 1823 38913
rect 2777 38947 2835 38953
rect 2777 38913 2789 38947
rect 2823 38913 2835 38947
rect 2777 38907 2835 38913
rect 3513 38947 3571 38953
rect 3513 38913 3525 38947
rect 3559 38944 3571 38947
rect 4706 38944 4712 38956
rect 3559 38916 4712 38944
rect 3559 38913 3571 38916
rect 3513 38907 3571 38913
rect 4706 38904 4712 38916
rect 4764 38904 4770 38956
rect 5644 38944 5672 38972
rect 6454 38944 6460 38956
rect 5644 38916 6460 38944
rect 6454 38904 6460 38916
rect 6512 38944 6518 38956
rect 6549 38947 6607 38953
rect 6549 38944 6561 38947
rect 6512 38916 6561 38944
rect 6512 38904 6518 38916
rect 6549 38913 6561 38916
rect 6595 38913 6607 38947
rect 6549 38907 6607 38913
rect 8202 38904 8208 38956
rect 8260 38944 8266 38956
rect 9861 38947 9919 38953
rect 9861 38944 9873 38947
rect 8260 38916 9873 38944
rect 8260 38904 8266 38916
rect 9861 38913 9873 38916
rect 9907 38913 9919 38947
rect 9861 38907 9919 38913
rect 1489 38879 1547 38885
rect 1489 38845 1501 38879
rect 1535 38845 1547 38879
rect 1489 38839 1547 38845
rect 1504 38740 1532 38839
rect 4338 38836 4344 38888
rect 4396 38876 4402 38888
rect 6365 38879 6423 38885
rect 6365 38876 6377 38879
rect 4396 38848 6377 38876
rect 4396 38836 4402 38848
rect 6365 38845 6377 38848
rect 6411 38845 6423 38879
rect 6365 38839 6423 38845
rect 2774 38768 2780 38820
rect 2832 38808 2838 38820
rect 4246 38808 4252 38820
rect 2832 38780 4252 38808
rect 2832 38768 2838 38780
rect 4246 38768 4252 38780
rect 4304 38768 4310 38820
rect 4522 38768 4528 38820
rect 4580 38808 4586 38820
rect 4706 38808 4712 38820
rect 4580 38780 4712 38808
rect 4580 38768 4586 38780
rect 4706 38768 4712 38780
rect 4764 38768 4770 38820
rect 2958 38740 2964 38752
rect 1044 38712 1532 38740
rect 2919 38712 2964 38740
rect 1044 38536 1072 38712
rect 2958 38700 2964 38712
rect 3016 38700 3022 38752
rect 3694 38740 3700 38752
rect 3655 38712 3700 38740
rect 3694 38700 3700 38712
rect 3752 38700 3758 38752
rect 4614 38700 4620 38752
rect 4672 38740 4678 38752
rect 7098 38740 7104 38752
rect 4672 38712 7104 38740
rect 4672 38700 4678 38712
rect 7098 38700 7104 38712
rect 7156 38700 7162 38752
rect 10042 38740 10048 38752
rect 10003 38712 10048 38740
rect 10042 38700 10048 38712
rect 10100 38700 10106 38752
rect 1104 38650 10856 38672
rect 1104 38598 2582 38650
rect 2634 38598 2646 38650
rect 2698 38598 2710 38650
rect 2762 38598 2774 38650
rect 2826 38598 2838 38650
rect 2890 38598 5846 38650
rect 5898 38598 5910 38650
rect 5962 38598 5974 38650
rect 6026 38598 6038 38650
rect 6090 38598 6102 38650
rect 6154 38598 9110 38650
rect 9162 38598 9174 38650
rect 9226 38598 9238 38650
rect 9290 38598 9302 38650
rect 9354 38598 9366 38650
rect 9418 38598 10856 38650
rect 1104 38576 10856 38598
rect 1486 38536 1492 38548
rect 1044 38508 1492 38536
rect 1486 38496 1492 38508
rect 1544 38496 1550 38548
rect 2406 38496 2412 38548
rect 2464 38536 2470 38548
rect 2961 38539 3019 38545
rect 2961 38536 2973 38539
rect 2464 38508 2973 38536
rect 2464 38496 2470 38508
rect 2961 38505 2973 38508
rect 3007 38505 3019 38539
rect 2961 38499 3019 38505
rect 5261 38539 5319 38545
rect 5261 38505 5273 38539
rect 5307 38536 5319 38539
rect 5350 38536 5356 38548
rect 5307 38508 5356 38536
rect 5307 38505 5319 38508
rect 5261 38499 5319 38505
rect 5350 38496 5356 38508
rect 5408 38496 5414 38548
rect 382 38360 388 38412
rect 440 38400 446 38412
rect 1765 38403 1823 38409
rect 1765 38400 1777 38403
rect 440 38372 1777 38400
rect 440 38360 446 38372
rect 1765 38369 1777 38372
rect 1811 38369 1823 38403
rect 1765 38363 1823 38369
rect 4430 38360 4436 38412
rect 4488 38400 4494 38412
rect 4488 38372 5120 38400
rect 4488 38360 4494 38372
rect 1489 38335 1547 38341
rect 1489 38301 1501 38335
rect 1535 38301 1547 38335
rect 1489 38295 1547 38301
rect 1504 38264 1532 38295
rect 3694 38292 3700 38344
rect 3752 38332 3758 38344
rect 4246 38332 4252 38344
rect 3752 38304 4252 38332
rect 3752 38292 3758 38304
rect 4246 38292 4252 38304
rect 4304 38292 4310 38344
rect 5092 38341 5120 38372
rect 4985 38335 5043 38341
rect 4985 38301 4997 38335
rect 5031 38301 5043 38335
rect 4985 38295 5043 38301
rect 5077 38335 5135 38341
rect 5077 38301 5089 38335
rect 5123 38332 5135 38335
rect 5350 38332 5356 38344
rect 5123 38304 5356 38332
rect 5123 38301 5135 38304
rect 5077 38295 5135 38301
rect 2682 38264 2688 38276
rect 1504 38236 2688 38264
rect 2682 38224 2688 38236
rect 2740 38224 2746 38276
rect 2869 38267 2927 38273
rect 2869 38233 2881 38267
rect 2915 38264 2927 38267
rect 3510 38264 3516 38276
rect 2915 38236 3516 38264
rect 2915 38233 2927 38236
rect 2869 38227 2927 38233
rect 3510 38224 3516 38236
rect 3568 38224 3574 38276
rect 5000 38264 5028 38295
rect 5350 38292 5356 38304
rect 5408 38292 5414 38344
rect 8478 38292 8484 38344
rect 8536 38332 8542 38344
rect 9861 38335 9919 38341
rect 9861 38332 9873 38335
rect 8536 38304 9873 38332
rect 8536 38292 8542 38304
rect 9861 38301 9873 38304
rect 9907 38301 9919 38335
rect 9861 38295 9919 38301
rect 5718 38264 5724 38276
rect 5000 38236 5724 38264
rect 5718 38224 5724 38236
rect 5776 38224 5782 38276
rect 10042 38196 10048 38208
rect 10003 38168 10048 38196
rect 10042 38156 10048 38168
rect 10100 38156 10106 38208
rect 1104 38106 10856 38128
rect 1104 38054 4214 38106
rect 4266 38054 4278 38106
rect 4330 38054 4342 38106
rect 4394 38054 4406 38106
rect 4458 38054 4470 38106
rect 4522 38054 7478 38106
rect 7530 38054 7542 38106
rect 7594 38054 7606 38106
rect 7658 38054 7670 38106
rect 7722 38054 7734 38106
rect 7786 38054 10856 38106
rect 1104 38032 10856 38054
rect 1486 37952 1492 38004
rect 1544 37992 1550 38004
rect 1857 37995 1915 38001
rect 1857 37992 1869 37995
rect 1544 37964 1869 37992
rect 1544 37952 1550 37964
rect 1857 37961 1869 37964
rect 1903 37961 1915 37995
rect 2682 37992 2688 38004
rect 2643 37964 2688 37992
rect 1857 37955 1915 37961
rect 2682 37952 2688 37964
rect 2740 37952 2746 38004
rect 5077 37995 5135 38001
rect 5077 37961 5089 37995
rect 5123 37992 5135 37995
rect 9766 37992 9772 38004
rect 5123 37964 9772 37992
rect 5123 37961 5135 37964
rect 5077 37955 5135 37961
rect 9766 37952 9772 37964
rect 9824 37952 9830 38004
rect 1026 37884 1032 37936
rect 1084 37924 1090 37936
rect 2774 37924 2780 37936
rect 1084 37896 1532 37924
rect 1084 37884 1090 37896
rect 1504 37865 1532 37896
rect 2332 37896 2780 37924
rect 2332 37865 2360 37896
rect 2774 37884 2780 37896
rect 2832 37884 2838 37936
rect 3418 37924 3424 37936
rect 3379 37896 3424 37924
rect 3418 37884 3424 37896
rect 3476 37884 3482 37936
rect 1489 37859 1547 37865
rect 1489 37825 1501 37859
rect 1535 37825 1547 37859
rect 1489 37819 1547 37825
rect 1673 37859 1731 37865
rect 1673 37825 1685 37859
rect 1719 37825 1731 37859
rect 1673 37819 1731 37825
rect 2317 37859 2375 37865
rect 2317 37825 2329 37859
rect 2363 37825 2375 37859
rect 2317 37819 2375 37825
rect 2501 37859 2559 37865
rect 2501 37825 2513 37859
rect 2547 37856 2559 37859
rect 2590 37856 2596 37868
rect 2547 37828 2596 37856
rect 2547 37825 2559 37828
rect 2501 37819 2559 37825
rect 1026 37748 1032 37800
rect 1084 37788 1090 37800
rect 1688 37788 1716 37819
rect 2516 37788 2544 37819
rect 2590 37816 2596 37828
rect 2648 37816 2654 37868
rect 2958 37816 2964 37868
rect 3016 37856 3022 37868
rect 3237 37859 3295 37865
rect 3237 37856 3249 37859
rect 3016 37828 3249 37856
rect 3016 37816 3022 37828
rect 3237 37825 3249 37828
rect 3283 37825 3295 37859
rect 3237 37819 3295 37825
rect 4893 37859 4951 37865
rect 4893 37825 4905 37859
rect 4939 37856 4951 37859
rect 5350 37856 5356 37868
rect 4939 37828 5356 37856
rect 4939 37825 4951 37828
rect 4893 37819 4951 37825
rect 5350 37816 5356 37828
rect 5408 37816 5414 37868
rect 1084 37760 2544 37788
rect 4709 37791 4767 37797
rect 1084 37748 1090 37760
rect 4709 37757 4721 37791
rect 4755 37757 4767 37791
rect 4709 37751 4767 37757
rect 4724 37720 4752 37751
rect 2746 37692 4752 37720
rect 1578 37612 1584 37664
rect 1636 37652 1642 37664
rect 2746 37652 2774 37692
rect 1636 37624 2774 37652
rect 1636 37612 1642 37624
rect 1104 37562 10856 37584
rect 1104 37510 2582 37562
rect 2634 37510 2646 37562
rect 2698 37510 2710 37562
rect 2762 37510 2774 37562
rect 2826 37510 2838 37562
rect 2890 37510 5846 37562
rect 5898 37510 5910 37562
rect 5962 37510 5974 37562
rect 6026 37510 6038 37562
rect 6090 37510 6102 37562
rect 6154 37510 9110 37562
rect 9162 37510 9174 37562
rect 9226 37510 9238 37562
rect 9290 37510 9302 37562
rect 9354 37510 9366 37562
rect 9418 37510 10856 37562
rect 1104 37488 10856 37510
rect 2406 37380 2412 37392
rect 2240 37352 2412 37380
rect 2240 37244 2268 37352
rect 2406 37340 2412 37352
rect 2464 37340 2470 37392
rect 2317 37315 2375 37321
rect 2317 37281 2329 37315
rect 2363 37312 2375 37315
rect 5718 37312 5724 37324
rect 2363 37284 5724 37312
rect 2363 37281 2375 37284
rect 2317 37275 2375 37281
rect 5718 37272 5724 37284
rect 5776 37272 5782 37324
rect 2501 37247 2559 37253
rect 2501 37244 2513 37247
rect 2240 37216 2513 37244
rect 2501 37213 2513 37216
rect 2547 37244 2559 37247
rect 2590 37244 2596 37256
rect 2547 37216 2596 37244
rect 2547 37213 2559 37216
rect 2501 37207 2559 37213
rect 2590 37204 2596 37216
rect 2648 37204 2654 37256
rect 2685 37247 2743 37253
rect 2685 37213 2697 37247
rect 2731 37244 2743 37247
rect 2958 37244 2964 37256
rect 2731 37216 2964 37244
rect 2731 37213 2743 37216
rect 2685 37207 2743 37213
rect 2958 37204 2964 37216
rect 3016 37204 3022 37256
rect 3786 37244 3792 37256
rect 3747 37216 3792 37244
rect 3786 37204 3792 37216
rect 3844 37204 3850 37256
rect 8389 37247 8447 37253
rect 8389 37213 8401 37247
rect 8435 37244 8447 37247
rect 8570 37244 8576 37256
rect 8435 37216 8576 37244
rect 8435 37213 8447 37216
rect 8389 37207 8447 37213
rect 8570 37204 8576 37216
rect 8628 37204 8634 37256
rect 9861 37247 9919 37253
rect 9861 37213 9873 37247
rect 9907 37213 9919 37247
rect 9861 37207 9919 37213
rect 1673 37179 1731 37185
rect 1673 37145 1685 37179
rect 1719 37176 1731 37179
rect 2406 37176 2412 37188
rect 1719 37148 2412 37176
rect 1719 37145 1731 37148
rect 1673 37139 1731 37145
rect 2406 37136 2412 37148
rect 2464 37136 2470 37188
rect 6362 37136 6368 37188
rect 6420 37176 6426 37188
rect 9876 37176 9904 37207
rect 6420 37148 9904 37176
rect 6420 37136 6426 37148
rect 1765 37111 1823 37117
rect 1765 37077 1777 37111
rect 1811 37108 1823 37111
rect 2682 37108 2688 37120
rect 1811 37080 2688 37108
rect 1811 37077 1823 37080
rect 1765 37071 1823 37077
rect 2682 37068 2688 37080
rect 2740 37068 2746 37120
rect 3970 37108 3976 37120
rect 3931 37080 3976 37108
rect 3970 37068 3976 37080
rect 4028 37068 4034 37120
rect 8202 37108 8208 37120
rect 8163 37080 8208 37108
rect 8202 37068 8208 37080
rect 8260 37068 8266 37120
rect 10042 37108 10048 37120
rect 10003 37080 10048 37108
rect 10042 37068 10048 37080
rect 10100 37068 10106 37120
rect 1104 37018 10856 37040
rect 1104 36966 4214 37018
rect 4266 36966 4278 37018
rect 4330 36966 4342 37018
rect 4394 36966 4406 37018
rect 4458 36966 4470 37018
rect 4522 36966 7478 37018
rect 7530 36966 7542 37018
rect 7594 36966 7606 37018
rect 7658 36966 7670 37018
rect 7722 36966 7734 37018
rect 7786 36966 10856 37018
rect 1104 36944 10856 36966
rect 2406 36904 2412 36916
rect 2367 36876 2412 36904
rect 2406 36864 2412 36876
rect 2464 36864 2470 36916
rect 3053 36907 3111 36913
rect 3053 36873 3065 36907
rect 3099 36904 3111 36907
rect 3786 36904 3792 36916
rect 3099 36876 3792 36904
rect 3099 36873 3111 36876
rect 3053 36867 3111 36873
rect 3786 36864 3792 36876
rect 3844 36864 3850 36916
rect 6362 36904 6368 36916
rect 6323 36876 6368 36904
rect 6362 36864 6368 36876
rect 6420 36864 6426 36916
rect 7009 36907 7067 36913
rect 7009 36873 7021 36907
rect 7055 36904 7067 36907
rect 8478 36904 8484 36916
rect 7055 36876 8484 36904
rect 7055 36873 7067 36876
rect 7009 36867 7067 36873
rect 8478 36864 8484 36876
rect 8536 36864 8542 36916
rect 6822 36836 6828 36848
rect 2884 36808 6828 36836
rect 2225 36771 2283 36777
rect 2225 36737 2237 36771
rect 2271 36768 2283 36771
rect 2590 36768 2596 36780
rect 2271 36740 2596 36768
rect 2271 36737 2283 36740
rect 2225 36731 2283 36737
rect 2590 36728 2596 36740
rect 2648 36728 2654 36780
rect 2884 36777 2912 36808
rect 6822 36796 6828 36808
rect 6880 36796 6886 36848
rect 2869 36771 2927 36777
rect 2869 36737 2881 36771
rect 2915 36737 2927 36771
rect 2869 36731 2927 36737
rect 3142 36728 3148 36780
rect 3200 36768 3206 36780
rect 3510 36768 3516 36780
rect 3200 36740 3516 36768
rect 3200 36728 3206 36740
rect 3510 36728 3516 36740
rect 3568 36728 3574 36780
rect 6546 36768 6552 36780
rect 6507 36740 6552 36768
rect 6546 36728 6552 36740
rect 6604 36728 6610 36780
rect 7190 36768 7196 36780
rect 7151 36740 7196 36768
rect 7190 36728 7196 36740
rect 7248 36728 7254 36780
rect 9858 36768 9864 36780
rect 9819 36740 9864 36768
rect 9858 36728 9864 36740
rect 9916 36728 9922 36780
rect 1578 36660 1584 36712
rect 1636 36700 1642 36712
rect 2041 36703 2099 36709
rect 2041 36700 2053 36703
rect 1636 36672 2053 36700
rect 1636 36660 1642 36672
rect 2041 36669 2053 36672
rect 2087 36700 2099 36703
rect 2406 36700 2412 36712
rect 2087 36672 2412 36700
rect 2087 36669 2099 36672
rect 2041 36663 2099 36669
rect 2406 36660 2412 36672
rect 2464 36660 2470 36712
rect 934 36592 940 36644
rect 992 36632 998 36644
rect 4062 36632 4068 36644
rect 992 36604 4068 36632
rect 992 36592 998 36604
rect 4062 36592 4068 36604
rect 4120 36592 4126 36644
rect 4614 36592 4620 36644
rect 4672 36632 4678 36644
rect 5442 36632 5448 36644
rect 4672 36604 5448 36632
rect 4672 36592 4678 36604
rect 5442 36592 5448 36604
rect 5500 36592 5506 36644
rect 5074 36524 5080 36576
rect 5132 36564 5138 36576
rect 5350 36564 5356 36576
rect 5132 36536 5356 36564
rect 5132 36524 5138 36536
rect 5350 36524 5356 36536
rect 5408 36524 5414 36576
rect 5534 36524 5540 36576
rect 5592 36564 5598 36576
rect 6454 36564 6460 36576
rect 5592 36536 6460 36564
rect 5592 36524 5598 36536
rect 6454 36524 6460 36536
rect 6512 36524 6518 36576
rect 10042 36564 10048 36576
rect 10003 36536 10048 36564
rect 10042 36524 10048 36536
rect 10100 36524 10106 36576
rect 1104 36474 10856 36496
rect 1104 36422 2582 36474
rect 2634 36422 2646 36474
rect 2698 36422 2710 36474
rect 2762 36422 2774 36474
rect 2826 36422 2838 36474
rect 2890 36422 5846 36474
rect 5898 36422 5910 36474
rect 5962 36422 5974 36474
rect 6026 36422 6038 36474
rect 6090 36422 6102 36474
rect 6154 36422 9110 36474
rect 9162 36422 9174 36474
rect 9226 36422 9238 36474
rect 9290 36422 9302 36474
rect 9354 36422 9366 36474
rect 9418 36422 10856 36474
rect 1104 36400 10856 36422
rect 1946 36360 1952 36372
rect 1907 36332 1952 36360
rect 1946 36320 1952 36332
rect 2004 36320 2010 36372
rect 3970 36360 3976 36372
rect 3931 36332 3976 36360
rect 3970 36320 3976 36332
rect 4028 36320 4034 36372
rect 4525 36363 4583 36369
rect 4525 36329 4537 36363
rect 4571 36360 4583 36363
rect 9858 36360 9864 36372
rect 4571 36332 9864 36360
rect 4571 36329 4583 36332
rect 4525 36323 4583 36329
rect 9858 36320 9864 36332
rect 9916 36320 9922 36372
rect 6638 36292 6644 36304
rect 2516 36264 6644 36292
rect 2516 36165 2544 36264
rect 6638 36252 6644 36264
rect 6696 36252 6702 36304
rect 6270 36224 6276 36236
rect 3804 36196 6276 36224
rect 3804 36165 3832 36196
rect 6270 36184 6276 36196
rect 6328 36184 6334 36236
rect 2501 36159 2559 36165
rect 2501 36125 2513 36159
rect 2547 36125 2559 36159
rect 2501 36119 2559 36125
rect 3789 36159 3847 36165
rect 3789 36125 3801 36159
rect 3835 36125 3847 36159
rect 4706 36156 4712 36168
rect 4667 36128 4712 36156
rect 3789 36119 3847 36125
rect 4706 36116 4712 36128
rect 4764 36116 4770 36168
rect 9858 36156 9864 36168
rect 9819 36128 9864 36156
rect 9858 36116 9864 36128
rect 9916 36116 9922 36168
rect 1857 36091 1915 36097
rect 1857 36057 1869 36091
rect 1903 36088 1915 36091
rect 1946 36088 1952 36100
rect 1903 36060 1952 36088
rect 1903 36057 1915 36060
rect 1857 36051 1915 36057
rect 1946 36048 1952 36060
rect 2004 36048 2010 36100
rect 2685 36023 2743 36029
rect 2685 35989 2697 36023
rect 2731 36020 2743 36023
rect 2774 36020 2780 36032
rect 2731 35992 2780 36020
rect 2731 35989 2743 35992
rect 2685 35983 2743 35989
rect 2774 35980 2780 35992
rect 2832 35980 2838 36032
rect 10042 36020 10048 36032
rect 10003 35992 10048 36020
rect 10042 35980 10048 35992
rect 10100 35980 10106 36032
rect 1104 35930 10856 35952
rect 1104 35878 4214 35930
rect 4266 35878 4278 35930
rect 4330 35878 4342 35930
rect 4394 35878 4406 35930
rect 4458 35878 4470 35930
rect 4522 35878 7478 35930
rect 7530 35878 7542 35930
rect 7594 35878 7606 35930
rect 7658 35878 7670 35930
rect 7722 35878 7734 35930
rect 7786 35878 10856 35930
rect 1104 35856 10856 35878
rect 2961 35819 3019 35825
rect 2961 35785 2973 35819
rect 3007 35816 3019 35819
rect 4706 35816 4712 35828
rect 3007 35788 4712 35816
rect 3007 35785 3019 35788
rect 2961 35779 3019 35785
rect 4706 35776 4712 35788
rect 4764 35776 4770 35828
rect 5445 35819 5503 35825
rect 5445 35785 5457 35819
rect 5491 35816 5503 35819
rect 6546 35816 6552 35828
rect 5491 35788 6552 35816
rect 5491 35785 5503 35788
rect 5445 35779 5503 35785
rect 6546 35776 6552 35788
rect 6604 35776 6610 35828
rect 6733 35819 6791 35825
rect 6733 35785 6745 35819
rect 6779 35816 6791 35819
rect 7190 35816 7196 35828
rect 6779 35788 7196 35816
rect 6779 35785 6791 35788
rect 6733 35779 6791 35785
rect 7190 35776 7196 35788
rect 7248 35776 7254 35828
rect 1397 35683 1455 35689
rect 1397 35649 1409 35683
rect 1443 35680 1455 35683
rect 2130 35680 2136 35692
rect 1443 35652 2136 35680
rect 1443 35649 1455 35652
rect 1397 35643 1455 35649
rect 2130 35640 2136 35652
rect 2188 35640 2194 35692
rect 2777 35683 2835 35689
rect 2777 35649 2789 35683
rect 2823 35680 2835 35683
rect 2958 35680 2964 35692
rect 2823 35652 2964 35680
rect 2823 35649 2835 35652
rect 2777 35643 2835 35649
rect 2958 35640 2964 35652
rect 3016 35640 3022 35692
rect 3970 35680 3976 35692
rect 3931 35652 3976 35680
rect 3970 35640 3976 35652
rect 4028 35640 4034 35692
rect 4341 35683 4399 35689
rect 4341 35649 4353 35683
rect 4387 35680 4399 35683
rect 5261 35683 5319 35689
rect 5261 35680 5273 35683
rect 4387 35652 5273 35680
rect 4387 35649 4399 35652
rect 4341 35643 4399 35649
rect 5261 35649 5273 35652
rect 5307 35680 5319 35683
rect 5534 35680 5540 35692
rect 5307 35652 5540 35680
rect 5307 35649 5319 35652
rect 5261 35643 5319 35649
rect 5534 35640 5540 35652
rect 5592 35680 5598 35692
rect 6270 35680 6276 35692
rect 5592 35652 6276 35680
rect 5592 35640 5598 35652
rect 6270 35640 6276 35652
rect 6328 35680 6334 35692
rect 6549 35683 6607 35689
rect 6549 35680 6561 35683
rect 6328 35652 6561 35680
rect 6328 35640 6334 35652
rect 6549 35649 6561 35652
rect 6595 35649 6607 35683
rect 6549 35643 6607 35649
rect 2593 35615 2651 35621
rect 2593 35612 2605 35615
rect 1412 35584 2605 35612
rect 1412 35556 1440 35584
rect 2593 35581 2605 35584
rect 2639 35581 2651 35615
rect 2593 35575 2651 35581
rect 4614 35572 4620 35624
rect 4672 35612 4678 35624
rect 5077 35615 5135 35621
rect 5077 35612 5089 35615
rect 4672 35584 5089 35612
rect 4672 35572 4678 35584
rect 5077 35581 5089 35584
rect 5123 35581 5135 35615
rect 6362 35612 6368 35624
rect 6323 35584 6368 35612
rect 5077 35575 5135 35581
rect 6362 35572 6368 35584
rect 6420 35572 6426 35624
rect 1394 35504 1400 35556
rect 1452 35504 1458 35556
rect 2130 35504 2136 35556
rect 2188 35544 2194 35556
rect 2406 35544 2412 35556
rect 2188 35516 2412 35544
rect 2188 35504 2194 35516
rect 2406 35504 2412 35516
rect 2464 35504 2470 35556
rect 1578 35476 1584 35488
rect 1539 35448 1584 35476
rect 1578 35436 1584 35448
rect 1636 35436 1642 35488
rect 1104 35386 10856 35408
rect 1104 35334 2582 35386
rect 2634 35334 2646 35386
rect 2698 35334 2710 35386
rect 2762 35334 2774 35386
rect 2826 35334 2838 35386
rect 2890 35334 5846 35386
rect 5898 35334 5910 35386
rect 5962 35334 5974 35386
rect 6026 35334 6038 35386
rect 6090 35334 6102 35386
rect 6154 35334 9110 35386
rect 9162 35334 9174 35386
rect 9226 35334 9238 35386
rect 9290 35334 9302 35386
rect 9354 35334 9366 35386
rect 9418 35334 10856 35386
rect 1104 35312 10856 35334
rect 3789 35275 3847 35281
rect 3789 35241 3801 35275
rect 3835 35272 3847 35275
rect 9858 35272 9864 35284
rect 3835 35244 9864 35272
rect 3835 35241 3847 35244
rect 3789 35235 3847 35241
rect 9858 35232 9864 35244
rect 9916 35232 9922 35284
rect 1486 35164 1492 35216
rect 1544 35204 1550 35216
rect 2590 35204 2596 35216
rect 1544 35176 2596 35204
rect 1544 35164 1550 35176
rect 2590 35164 2596 35176
rect 2648 35164 2654 35216
rect 1397 35071 1455 35077
rect 1397 35037 1409 35071
rect 1443 35068 1455 35071
rect 1670 35068 1676 35080
rect 1443 35040 1676 35068
rect 1443 35037 1455 35040
rect 1397 35031 1455 35037
rect 1670 35028 1676 35040
rect 1728 35028 1734 35080
rect 2038 35028 2044 35080
rect 2096 35068 2102 35080
rect 2133 35071 2191 35077
rect 2133 35068 2145 35071
rect 2096 35040 2145 35068
rect 2096 35028 2102 35040
rect 2133 35037 2145 35040
rect 2179 35037 2191 35071
rect 2133 35031 2191 35037
rect 3142 35028 3148 35080
rect 3200 35068 3206 35080
rect 3973 35071 4031 35077
rect 3973 35068 3985 35071
rect 3200 35040 3985 35068
rect 3200 35028 3206 35040
rect 3973 35037 3985 35040
rect 4019 35037 4031 35071
rect 3973 35031 4031 35037
rect 4062 35028 4068 35080
rect 4120 35068 4126 35080
rect 9861 35071 9919 35077
rect 9861 35068 9873 35071
rect 4120 35040 9873 35068
rect 4120 35028 4126 35040
rect 9861 35037 9873 35040
rect 9907 35037 9919 35071
rect 9861 35031 9919 35037
rect 1578 34932 1584 34944
rect 1539 34904 1584 34932
rect 1578 34892 1584 34904
rect 1636 34892 1642 34944
rect 2314 34932 2320 34944
rect 2275 34904 2320 34932
rect 2314 34892 2320 34904
rect 2372 34892 2378 34944
rect 10042 34932 10048 34944
rect 10003 34904 10048 34932
rect 10042 34892 10048 34904
rect 10100 34892 10106 34944
rect 1104 34842 10856 34864
rect 1104 34790 4214 34842
rect 4266 34790 4278 34842
rect 4330 34790 4342 34842
rect 4394 34790 4406 34842
rect 4458 34790 4470 34842
rect 4522 34790 7478 34842
rect 7530 34790 7542 34842
rect 7594 34790 7606 34842
rect 7658 34790 7670 34842
rect 7722 34790 7734 34842
rect 7786 34790 10856 34842
rect 1104 34768 10856 34790
rect 1486 34688 1492 34740
rect 1544 34728 1550 34740
rect 1581 34731 1639 34737
rect 1581 34728 1593 34731
rect 1544 34700 1593 34728
rect 1544 34688 1550 34700
rect 1581 34697 1593 34700
rect 1627 34697 1639 34731
rect 1581 34691 1639 34697
rect 3789 34731 3847 34737
rect 3789 34697 3801 34731
rect 3835 34728 3847 34731
rect 4062 34728 4068 34740
rect 3835 34700 4068 34728
rect 3835 34697 3847 34700
rect 3789 34691 3847 34697
rect 4062 34688 4068 34700
rect 4120 34688 4126 34740
rect 9582 34688 9588 34740
rect 9640 34728 9646 34740
rect 10045 34731 10103 34737
rect 10045 34728 10057 34731
rect 9640 34700 10057 34728
rect 9640 34688 9646 34700
rect 10045 34697 10057 34700
rect 10091 34697 10103 34731
rect 10045 34691 10103 34697
rect 566 34552 572 34604
rect 624 34592 630 34604
rect 1397 34595 1455 34601
rect 1397 34592 1409 34595
rect 624 34564 1409 34592
rect 624 34552 630 34564
rect 1397 34561 1409 34564
rect 1443 34561 1455 34595
rect 1397 34555 1455 34561
rect 1854 34552 1860 34604
rect 1912 34592 1918 34604
rect 2133 34595 2191 34601
rect 2133 34592 2145 34595
rect 1912 34564 2145 34592
rect 1912 34552 1918 34564
rect 2133 34561 2145 34564
rect 2179 34561 2191 34595
rect 2133 34555 2191 34561
rect 2590 34552 2596 34604
rect 2648 34592 2654 34604
rect 2869 34595 2927 34601
rect 2869 34592 2881 34595
rect 2648 34564 2881 34592
rect 2648 34552 2654 34564
rect 2869 34561 2881 34564
rect 2915 34561 2927 34595
rect 2869 34555 2927 34561
rect 3973 34595 4031 34601
rect 3973 34561 3985 34595
rect 4019 34561 4031 34595
rect 3973 34555 4031 34561
rect 2222 34524 2228 34536
rect 584 34496 2228 34524
rect 584 34468 612 34496
rect 2222 34484 2228 34496
rect 2280 34484 2286 34536
rect 3988 34468 4016 34555
rect 5534 34552 5540 34604
rect 5592 34592 5598 34604
rect 9861 34595 9919 34601
rect 9861 34592 9873 34595
rect 5592 34564 9873 34592
rect 5592 34552 5598 34564
rect 9861 34561 9873 34564
rect 9907 34561 9919 34595
rect 9861 34555 9919 34561
rect 566 34416 572 34468
rect 624 34416 630 34468
rect 1854 34416 1860 34468
rect 1912 34456 1918 34468
rect 2130 34456 2136 34468
rect 1912 34428 2136 34456
rect 1912 34416 1918 34428
rect 2130 34416 2136 34428
rect 2188 34416 2194 34468
rect 3970 34416 3976 34468
rect 4028 34416 4034 34468
rect 2222 34348 2228 34400
rect 2280 34388 2286 34400
rect 2317 34391 2375 34397
rect 2317 34388 2329 34391
rect 2280 34360 2329 34388
rect 2280 34348 2286 34360
rect 2317 34357 2329 34360
rect 2363 34357 2375 34391
rect 3050 34388 3056 34400
rect 3011 34360 3056 34388
rect 2317 34351 2375 34357
rect 3050 34348 3056 34360
rect 3108 34348 3114 34400
rect 1104 34298 10856 34320
rect 1104 34246 2582 34298
rect 2634 34246 2646 34298
rect 2698 34246 2710 34298
rect 2762 34246 2774 34298
rect 2826 34246 2838 34298
rect 2890 34246 5846 34298
rect 5898 34246 5910 34298
rect 5962 34246 5974 34298
rect 6026 34246 6038 34298
rect 6090 34246 6102 34298
rect 6154 34246 9110 34298
rect 9162 34246 9174 34298
rect 9226 34246 9238 34298
rect 9290 34246 9302 34298
rect 9354 34246 9366 34298
rect 9418 34246 10856 34298
rect 1104 34224 10856 34246
rect 842 34144 848 34196
rect 900 34184 906 34196
rect 1949 34187 2007 34193
rect 1949 34184 1961 34187
rect 900 34156 1961 34184
rect 900 34144 906 34156
rect 1949 34153 1961 34156
rect 1995 34153 2007 34187
rect 1949 34147 2007 34153
rect 5353 34187 5411 34193
rect 5353 34153 5365 34187
rect 5399 34184 5411 34187
rect 8570 34184 8576 34196
rect 5399 34156 8576 34184
rect 5399 34153 5411 34156
rect 5353 34147 5411 34153
rect 8570 34144 8576 34156
rect 8628 34144 8634 34196
rect 198 34076 204 34128
rect 256 34116 262 34128
rect 2777 34119 2835 34125
rect 2777 34116 2789 34119
rect 256 34088 2789 34116
rect 256 34076 262 34088
rect 2777 34085 2789 34088
rect 2823 34085 2835 34119
rect 2777 34079 2835 34085
rect 5626 34076 5632 34128
rect 5684 34116 5690 34128
rect 5810 34116 5816 34128
rect 5684 34088 5816 34116
rect 5684 34076 5690 34088
rect 5810 34076 5816 34088
rect 5868 34076 5874 34128
rect 842 33940 848 33992
rect 900 33980 906 33992
rect 4985 33983 5043 33989
rect 4985 33980 4997 33983
rect 900 33952 4997 33980
rect 900 33940 906 33952
rect 4985 33949 4997 33952
rect 5031 33949 5043 33983
rect 4985 33943 5043 33949
rect 5169 33983 5227 33989
rect 5169 33949 5181 33983
rect 5215 33980 5227 33983
rect 5626 33980 5632 33992
rect 5215 33952 5632 33980
rect 5215 33949 5227 33952
rect 5169 33943 5227 33949
rect 5626 33940 5632 33952
rect 5684 33980 5690 33992
rect 6270 33980 6276 33992
rect 5684 33952 6276 33980
rect 5684 33940 5690 33952
rect 6270 33940 6276 33952
rect 6328 33940 6334 33992
rect 1857 33915 1915 33921
rect 1857 33881 1869 33915
rect 1903 33912 1915 33915
rect 2130 33912 2136 33924
rect 1903 33884 2136 33912
rect 1903 33881 1915 33884
rect 1857 33875 1915 33881
rect 2130 33872 2136 33884
rect 2188 33872 2194 33924
rect 2593 33915 2651 33921
rect 2593 33881 2605 33915
rect 2639 33912 2651 33915
rect 2958 33912 2964 33924
rect 2639 33884 2964 33912
rect 2639 33881 2651 33884
rect 2593 33875 2651 33881
rect 2958 33872 2964 33884
rect 3016 33872 3022 33924
rect 2406 33804 2412 33856
rect 2464 33844 2470 33856
rect 6362 33844 6368 33856
rect 2464 33816 6368 33844
rect 2464 33804 2470 33816
rect 6362 33804 6368 33816
rect 6420 33804 6426 33856
rect 1104 33754 10856 33776
rect 1104 33702 4214 33754
rect 4266 33702 4278 33754
rect 4330 33702 4342 33754
rect 4394 33702 4406 33754
rect 4458 33702 4470 33754
rect 4522 33702 7478 33754
rect 7530 33702 7542 33754
rect 7594 33702 7606 33754
rect 7658 33702 7670 33754
rect 7722 33702 7734 33754
rect 7786 33702 10856 33754
rect 1104 33680 10856 33702
rect 1854 33640 1860 33652
rect 1412 33612 1860 33640
rect 1412 33584 1440 33612
rect 1854 33600 1860 33612
rect 1912 33600 1918 33652
rect 2130 33640 2136 33652
rect 2091 33612 2136 33640
rect 2130 33600 2136 33612
rect 2188 33600 2194 33652
rect 2958 33640 2964 33652
rect 2919 33612 2964 33640
rect 2958 33600 2964 33612
rect 3016 33600 3022 33652
rect 3789 33643 3847 33649
rect 3789 33609 3801 33643
rect 3835 33640 3847 33643
rect 3970 33640 3976 33652
rect 3835 33612 3976 33640
rect 3835 33609 3847 33612
rect 3789 33603 3847 33609
rect 3970 33600 3976 33612
rect 4028 33600 4034 33652
rect 4249 33643 4307 33649
rect 4249 33609 4261 33643
rect 4295 33640 4307 33643
rect 5534 33640 5540 33652
rect 4295 33612 5540 33640
rect 4295 33609 4307 33612
rect 4249 33603 4307 33609
rect 5534 33600 5540 33612
rect 5592 33600 5598 33652
rect 5721 33643 5779 33649
rect 5721 33609 5733 33643
rect 5767 33640 5779 33643
rect 8754 33640 8760 33652
rect 5767 33612 8760 33640
rect 5767 33609 5779 33612
rect 5721 33603 5779 33609
rect 8754 33600 8760 33612
rect 8812 33600 8818 33652
rect 1394 33532 1400 33584
rect 1452 33532 1458 33584
rect 2406 33572 2412 33584
rect 1872 33544 2412 33572
rect 1872 33513 1900 33544
rect 2406 33532 2412 33544
rect 2464 33532 2470 33584
rect 2976 33544 5488 33572
rect 1857 33507 1915 33513
rect 1857 33473 1869 33507
rect 1903 33473 1915 33507
rect 1857 33467 1915 33473
rect 1946 33464 1952 33516
rect 2004 33504 2010 33516
rect 2777 33507 2835 33513
rect 2777 33504 2789 33507
rect 2004 33476 2789 33504
rect 2004 33464 2010 33476
rect 2777 33473 2789 33476
rect 2823 33473 2835 33507
rect 2777 33467 2835 33473
rect 2593 33439 2651 33445
rect 2593 33436 2605 33439
rect 1964 33408 2605 33436
rect 1964 33380 1992 33408
rect 2593 33405 2605 33408
rect 2639 33436 2651 33439
rect 2976 33436 3004 33544
rect 5460 33513 5488 33544
rect 3605 33507 3663 33513
rect 3605 33473 3617 33507
rect 3651 33473 3663 33507
rect 3605 33467 3663 33473
rect 4433 33507 4491 33513
rect 4433 33473 4445 33507
rect 4479 33504 4491 33507
rect 5445 33507 5503 33513
rect 4479 33476 4660 33504
rect 4479 33473 4491 33476
rect 4433 33467 4491 33473
rect 2639 33408 3004 33436
rect 3421 33439 3479 33445
rect 2639 33405 2651 33408
rect 2593 33399 2651 33405
rect 3421 33405 3433 33439
rect 3467 33405 3479 33439
rect 3421 33399 3479 33405
rect 1026 33328 1032 33380
rect 1084 33368 1090 33380
rect 1854 33368 1860 33380
rect 1084 33340 1860 33368
rect 1084 33328 1090 33340
rect 1854 33328 1860 33340
rect 1912 33328 1918 33380
rect 1946 33328 1952 33380
rect 2004 33328 2010 33380
rect 2406 33328 2412 33380
rect 2464 33368 2470 33380
rect 3436 33368 3464 33399
rect 2464 33340 3464 33368
rect 2464 33328 2470 33340
rect 2958 33260 2964 33312
rect 3016 33300 3022 33312
rect 3620 33300 3648 33467
rect 4632 33448 4660 33476
rect 5445 33473 5457 33507
rect 5491 33473 5503 33507
rect 5445 33467 5503 33473
rect 5537 33507 5595 33513
rect 5537 33473 5549 33507
rect 5583 33504 5595 33507
rect 5626 33504 5632 33516
rect 5583 33476 5632 33504
rect 5583 33473 5595 33476
rect 5537 33467 5595 33473
rect 5626 33464 5632 33476
rect 5684 33464 5690 33516
rect 9858 33504 9864 33516
rect 9819 33476 9864 33504
rect 9858 33464 9864 33476
rect 9916 33464 9922 33516
rect 4614 33396 4620 33448
rect 4672 33396 4678 33448
rect 5626 33328 5632 33380
rect 5684 33368 5690 33380
rect 5810 33368 5816 33380
rect 5684 33340 5816 33368
rect 5684 33328 5690 33340
rect 5810 33328 5816 33340
rect 5868 33328 5874 33380
rect 10042 33368 10048 33380
rect 10003 33340 10048 33368
rect 10042 33328 10048 33340
rect 10100 33328 10106 33380
rect 3016 33272 3648 33300
rect 3016 33260 3022 33272
rect 1104 33210 10856 33232
rect 1104 33158 2582 33210
rect 2634 33158 2646 33210
rect 2698 33158 2710 33210
rect 2762 33158 2774 33210
rect 2826 33158 2838 33210
rect 2890 33158 5846 33210
rect 5898 33158 5910 33210
rect 5962 33158 5974 33210
rect 6026 33158 6038 33210
rect 6090 33158 6102 33210
rect 6154 33158 9110 33210
rect 9162 33158 9174 33210
rect 9226 33158 9238 33210
rect 9290 33158 9302 33210
rect 9354 33158 9366 33210
rect 9418 33158 10856 33210
rect 1104 33136 10856 33158
rect 290 33056 296 33108
rect 348 33096 354 33108
rect 2225 33099 2283 33105
rect 2225 33096 2237 33099
rect 348 33068 2237 33096
rect 348 33056 354 33068
rect 2225 33065 2237 33068
rect 2271 33065 2283 33099
rect 3142 33096 3148 33108
rect 3103 33068 3148 33096
rect 2225 33059 2283 33065
rect 3142 33056 3148 33068
rect 3200 33056 3206 33108
rect 3694 32988 3700 33040
rect 3752 33028 3758 33040
rect 4709 33031 4767 33037
rect 4709 33028 4721 33031
rect 3752 33000 4721 33028
rect 3752 32988 3758 33000
rect 4709 32997 4721 33000
rect 4755 32997 4767 33031
rect 4709 32991 4767 32997
rect 1670 32920 1676 32972
rect 1728 32960 1734 32972
rect 9674 32960 9680 32972
rect 1728 32932 2912 32960
rect 1728 32920 1734 32932
rect 2314 32852 2320 32904
rect 2372 32892 2378 32904
rect 2777 32895 2835 32901
rect 2777 32892 2789 32895
rect 2372 32864 2789 32892
rect 2372 32852 2378 32864
rect 2777 32861 2789 32864
rect 2823 32861 2835 32895
rect 2777 32855 2835 32861
rect 2133 32827 2191 32833
rect 2133 32793 2145 32827
rect 2179 32824 2191 32827
rect 2590 32824 2596 32836
rect 2179 32796 2596 32824
rect 2179 32793 2191 32796
rect 2133 32787 2191 32793
rect 2590 32784 2596 32796
rect 2648 32784 2654 32836
rect 2884 32824 2912 32932
rect 4540 32932 9680 32960
rect 2958 32852 2964 32904
rect 3016 32892 3022 32904
rect 4540 32901 4568 32932
rect 9674 32920 9680 32932
rect 9732 32920 9738 32972
rect 3789 32895 3847 32901
rect 3016 32864 3061 32892
rect 3016 32852 3022 32864
rect 3789 32861 3801 32895
rect 3835 32892 3847 32895
rect 4341 32895 4399 32901
rect 4341 32892 4353 32895
rect 3835 32864 4353 32892
rect 3835 32861 3847 32864
rect 3789 32855 3847 32861
rect 4341 32861 4353 32864
rect 4387 32861 4399 32895
rect 4341 32855 4399 32861
rect 4525 32895 4583 32901
rect 4525 32861 4537 32895
rect 4571 32861 4583 32895
rect 4525 32855 4583 32861
rect 3804 32824 3832 32855
rect 7834 32852 7840 32904
rect 7892 32892 7898 32904
rect 9861 32895 9919 32901
rect 9861 32892 9873 32895
rect 7892 32864 9873 32892
rect 7892 32852 7898 32864
rect 9861 32861 9873 32864
rect 9907 32861 9919 32895
rect 9861 32855 9919 32861
rect 2884 32796 3832 32824
rect 3970 32756 3976 32768
rect 3931 32728 3976 32756
rect 3970 32716 3976 32728
rect 4028 32716 4034 32768
rect 10042 32756 10048 32768
rect 10003 32728 10048 32756
rect 10042 32716 10048 32728
rect 10100 32716 10106 32768
rect 1104 32666 10856 32688
rect 1104 32614 4214 32666
rect 4266 32614 4278 32666
rect 4330 32614 4342 32666
rect 4394 32614 4406 32666
rect 4458 32614 4470 32666
rect 4522 32614 7478 32666
rect 7530 32614 7542 32666
rect 7594 32614 7606 32666
rect 7658 32614 7670 32666
rect 7722 32614 7734 32666
rect 7786 32614 10856 32666
rect 1104 32592 10856 32614
rect 750 32512 756 32564
rect 808 32552 814 32564
rect 2590 32552 2596 32564
rect 808 32524 2360 32552
rect 2551 32524 2596 32552
rect 808 32512 814 32524
rect 2332 32484 2360 32524
rect 2590 32512 2596 32524
rect 2648 32512 2654 32564
rect 3234 32552 3240 32564
rect 3195 32524 3240 32552
rect 3234 32512 3240 32524
rect 3292 32512 3298 32564
rect 2332 32456 3832 32484
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32416 1639 32419
rect 1762 32416 1768 32428
rect 1627 32388 1768 32416
rect 1627 32385 1639 32388
rect 1581 32379 1639 32385
rect 1762 32376 1768 32388
rect 1820 32376 1826 32428
rect 1854 32376 1860 32428
rect 1912 32416 1918 32428
rect 2409 32419 2467 32425
rect 2409 32416 2421 32419
rect 1912 32388 2421 32416
rect 1912 32376 1918 32388
rect 2409 32385 2421 32388
rect 2455 32385 2467 32419
rect 2409 32379 2467 32385
rect 3145 32419 3203 32425
rect 3145 32385 3157 32419
rect 3191 32416 3203 32419
rect 3694 32416 3700 32428
rect 3191 32388 3700 32416
rect 3191 32385 3203 32388
rect 3145 32379 3203 32385
rect 3694 32376 3700 32388
rect 3752 32376 3758 32428
rect 3804 32425 3832 32456
rect 4430 32444 4436 32496
rect 4488 32484 4494 32496
rect 4798 32484 4804 32496
rect 4488 32456 4804 32484
rect 4488 32444 4494 32456
rect 4798 32444 4804 32456
rect 4856 32444 4862 32496
rect 3789 32419 3847 32425
rect 3789 32385 3801 32419
rect 3835 32385 3847 32419
rect 3789 32379 3847 32385
rect 842 32308 848 32360
rect 900 32348 906 32360
rect 2225 32351 2283 32357
rect 2225 32348 2237 32351
rect 900 32320 2237 32348
rect 900 32308 906 32320
rect 2225 32317 2237 32320
rect 2271 32317 2283 32351
rect 2225 32311 2283 32317
rect 3234 32308 3240 32360
rect 3292 32348 3298 32360
rect 3418 32348 3424 32360
rect 3292 32320 3424 32348
rect 3292 32308 3298 32320
rect 3418 32308 3424 32320
rect 3476 32308 3482 32360
rect 1765 32283 1823 32289
rect 1765 32249 1777 32283
rect 1811 32280 1823 32283
rect 5626 32280 5632 32292
rect 1811 32252 5632 32280
rect 1811 32249 1823 32252
rect 1765 32243 1823 32249
rect 5626 32240 5632 32252
rect 5684 32240 5690 32292
rect 3970 32212 3976 32224
rect 3931 32184 3976 32212
rect 3970 32172 3976 32184
rect 4028 32172 4034 32224
rect 1104 32122 10856 32144
rect 1104 32070 2582 32122
rect 2634 32070 2646 32122
rect 2698 32070 2710 32122
rect 2762 32070 2774 32122
rect 2826 32070 2838 32122
rect 2890 32070 5846 32122
rect 5898 32070 5910 32122
rect 5962 32070 5974 32122
rect 6026 32070 6038 32122
rect 6090 32070 6102 32122
rect 6154 32070 9110 32122
rect 9162 32070 9174 32122
rect 9226 32070 9238 32122
rect 9290 32070 9302 32122
rect 9354 32070 9366 32122
rect 9418 32070 10856 32122
rect 1104 32048 10856 32070
rect 1762 32008 1768 32020
rect 1723 31980 1768 32008
rect 1762 31968 1768 31980
rect 1820 31968 1826 32020
rect 2406 32008 2412 32020
rect 1964 31980 2412 32008
rect 934 31900 940 31952
rect 992 31940 998 31952
rect 1670 31940 1676 31952
rect 992 31912 1676 31940
rect 992 31900 998 31912
rect 1670 31900 1676 31912
rect 1728 31900 1734 31952
rect 1397 31875 1455 31881
rect 1397 31841 1409 31875
rect 1443 31872 1455 31875
rect 1964 31872 1992 31980
rect 2406 31968 2412 31980
rect 2464 32008 2470 32020
rect 2961 32011 3019 32017
rect 2464 31980 2728 32008
rect 2464 31968 2470 31980
rect 2700 31952 2728 31980
rect 2961 31977 2973 32011
rect 3007 32008 3019 32011
rect 4614 32008 4620 32020
rect 3007 31980 4620 32008
rect 3007 31977 3019 31980
rect 2961 31971 3019 31977
rect 4614 31968 4620 31980
rect 4672 31968 4678 32020
rect 4890 31968 4896 32020
rect 4948 31968 4954 32020
rect 2038 31900 2044 31952
rect 2096 31940 2102 31952
rect 2096 31912 2360 31940
rect 2096 31900 2102 31912
rect 1443 31844 1992 31872
rect 1443 31841 1455 31844
rect 1397 31835 1455 31841
rect 1486 31764 1492 31816
rect 1544 31804 1550 31816
rect 1581 31807 1639 31813
rect 1581 31804 1593 31807
rect 1544 31776 1593 31804
rect 1544 31764 1550 31776
rect 1581 31773 1593 31776
rect 1627 31804 1639 31807
rect 1854 31804 1860 31816
rect 1627 31776 1860 31804
rect 1627 31773 1639 31776
rect 1581 31767 1639 31773
rect 1854 31764 1860 31776
rect 1912 31764 1918 31816
rect 2332 31804 2360 31912
rect 2682 31900 2688 31952
rect 2740 31900 2746 31952
rect 3418 31900 3424 31952
rect 3476 31940 3482 31952
rect 3878 31940 3884 31952
rect 3476 31912 3884 31940
rect 3476 31900 3482 31912
rect 3878 31900 3884 31912
rect 3936 31900 3942 31952
rect 4430 31832 4436 31884
rect 4488 31872 4494 31884
rect 4488 31844 4844 31872
rect 4488 31832 4494 31844
rect 4816 31816 4844 31844
rect 2406 31804 2412 31816
rect 2332 31776 2412 31804
rect 2406 31764 2412 31776
rect 2464 31764 2470 31816
rect 2593 31807 2651 31813
rect 2593 31773 2605 31807
rect 2639 31773 2651 31807
rect 2774 31804 2780 31816
rect 2735 31776 2780 31804
rect 2593 31767 2651 31773
rect 1670 31696 1676 31748
rect 1728 31736 1734 31748
rect 2130 31736 2136 31748
rect 1728 31708 2136 31736
rect 1728 31696 1734 31708
rect 2130 31696 2136 31708
rect 2188 31696 2194 31748
rect 934 31628 940 31680
rect 992 31668 998 31680
rect 1762 31668 1768 31680
rect 992 31640 1768 31668
rect 992 31628 998 31640
rect 1762 31628 1768 31640
rect 1820 31628 1826 31680
rect 1854 31628 1860 31680
rect 1912 31668 1918 31680
rect 2608 31668 2636 31767
rect 2774 31764 2780 31776
rect 2832 31764 2838 31816
rect 3326 31764 3332 31816
rect 3384 31804 3390 31816
rect 3789 31807 3847 31813
rect 3789 31804 3801 31807
rect 3384 31776 3801 31804
rect 3384 31764 3390 31776
rect 3789 31773 3801 31776
rect 3835 31773 3847 31807
rect 3789 31767 3847 31773
rect 4798 31764 4804 31816
rect 4856 31764 4862 31816
rect 1912 31640 2636 31668
rect 1912 31628 1918 31640
rect 3326 31628 3332 31680
rect 3384 31668 3390 31680
rect 3973 31671 4031 31677
rect 3973 31668 3985 31671
rect 3384 31640 3985 31668
rect 3384 31628 3390 31640
rect 3973 31637 3985 31640
rect 4019 31637 4031 31671
rect 3973 31631 4031 31637
rect 4706 31628 4712 31680
rect 4764 31668 4770 31680
rect 4908 31668 4936 31968
rect 10042 31940 10048 31952
rect 10003 31912 10048 31940
rect 10042 31900 10048 31912
rect 10100 31900 10106 31952
rect 7926 31764 7932 31816
rect 7984 31804 7990 31816
rect 9861 31807 9919 31813
rect 9861 31804 9873 31807
rect 7984 31776 9873 31804
rect 7984 31764 7990 31776
rect 9861 31773 9873 31776
rect 9907 31773 9919 31807
rect 9861 31767 9919 31773
rect 4764 31640 4936 31668
rect 4764 31628 4770 31640
rect 1104 31578 10856 31600
rect 1104 31526 4214 31578
rect 4266 31526 4278 31578
rect 4330 31526 4342 31578
rect 4394 31526 4406 31578
rect 4458 31526 4470 31578
rect 4522 31526 7478 31578
rect 7530 31526 7542 31578
rect 7594 31526 7606 31578
rect 7658 31526 7670 31578
rect 7722 31526 7734 31578
rect 7786 31526 10856 31578
rect 1104 31504 10856 31526
rect 566 31424 572 31476
rect 624 31464 630 31476
rect 1026 31464 1032 31476
rect 624 31436 1032 31464
rect 624 31424 630 31436
rect 1026 31424 1032 31436
rect 1084 31424 1090 31476
rect 3050 31424 3056 31476
rect 3108 31464 3114 31476
rect 3234 31464 3240 31476
rect 3108 31436 3240 31464
rect 3108 31424 3114 31436
rect 3234 31424 3240 31436
rect 3292 31424 3298 31476
rect 5074 31424 5080 31476
rect 5132 31464 5138 31476
rect 5258 31464 5264 31476
rect 5132 31436 5264 31464
rect 5132 31424 5138 31436
rect 5258 31424 5264 31436
rect 5316 31424 5322 31476
rect 2225 31399 2283 31405
rect 2225 31365 2237 31399
rect 2271 31396 2283 31399
rect 6178 31396 6184 31408
rect 2271 31368 6184 31396
rect 2271 31365 2283 31368
rect 2225 31359 2283 31365
rect 6178 31356 6184 31368
rect 6236 31356 6242 31408
rect 2038 31328 2044 31340
rect 1999 31300 2044 31328
rect 2038 31288 2044 31300
rect 2096 31288 2102 31340
rect 2314 31288 2320 31340
rect 2372 31288 2378 31340
rect 2590 31288 2596 31340
rect 2648 31328 2654 31340
rect 2685 31331 2743 31337
rect 2685 31328 2697 31331
rect 2648 31300 2697 31328
rect 2648 31288 2654 31300
rect 2685 31297 2697 31300
rect 2731 31297 2743 31331
rect 2685 31291 2743 31297
rect 3421 31331 3479 31337
rect 3421 31297 3433 31331
rect 3467 31328 3479 31331
rect 3602 31328 3608 31340
rect 3467 31300 3608 31328
rect 3467 31297 3479 31300
rect 3421 31291 3479 31297
rect 3602 31288 3608 31300
rect 3660 31288 3666 31340
rect 5074 31288 5080 31340
rect 5132 31328 5138 31340
rect 9861 31331 9919 31337
rect 9861 31328 9873 31331
rect 5132 31300 9873 31328
rect 5132 31288 5138 31300
rect 9861 31297 9873 31300
rect 9907 31297 9919 31331
rect 9861 31291 9919 31297
rect 2222 31084 2228 31136
rect 2280 31124 2286 31136
rect 2332 31124 2360 31288
rect 3602 31192 3608 31204
rect 3563 31164 3608 31192
rect 3602 31152 3608 31164
rect 3660 31152 3666 31204
rect 2280 31096 2360 31124
rect 2869 31127 2927 31133
rect 2280 31084 2286 31096
rect 2869 31093 2881 31127
rect 2915 31124 2927 31127
rect 2958 31124 2964 31136
rect 2915 31096 2964 31124
rect 2915 31093 2927 31096
rect 2869 31087 2927 31093
rect 2958 31084 2964 31096
rect 3016 31084 3022 31136
rect 10042 31124 10048 31136
rect 10003 31096 10048 31124
rect 10042 31084 10048 31096
rect 10100 31084 10106 31136
rect 1104 31034 10856 31056
rect 1104 30982 2582 31034
rect 2634 30982 2646 31034
rect 2698 30982 2710 31034
rect 2762 30982 2774 31034
rect 2826 30982 2838 31034
rect 2890 30982 5846 31034
rect 5898 30982 5910 31034
rect 5962 30982 5974 31034
rect 6026 30982 6038 31034
rect 6090 30982 6102 31034
rect 6154 30982 9110 31034
rect 9162 30982 9174 31034
rect 9226 30982 9238 31034
rect 9290 30982 9302 31034
rect 9354 30982 9366 31034
rect 9418 30982 10856 31034
rect 1104 30960 10856 30982
rect 2038 30880 2044 30932
rect 2096 30920 2102 30932
rect 2501 30923 2559 30929
rect 2501 30920 2513 30923
rect 2096 30892 2513 30920
rect 2096 30880 2102 30892
rect 2501 30889 2513 30892
rect 2547 30889 2559 30923
rect 2501 30883 2559 30889
rect 1486 30744 1492 30796
rect 1544 30744 1550 30796
rect 1854 30744 1860 30796
rect 1912 30784 1918 30796
rect 2038 30784 2044 30796
rect 1912 30756 2044 30784
rect 1912 30744 1918 30756
rect 2038 30744 2044 30756
rect 2096 30784 2102 30796
rect 2133 30787 2191 30793
rect 2133 30784 2145 30787
rect 2096 30756 2145 30784
rect 2096 30744 2102 30756
rect 2133 30753 2145 30756
rect 2179 30753 2191 30787
rect 2133 30747 2191 30753
rect 750 30676 756 30728
rect 808 30716 814 30728
rect 1504 30716 1532 30744
rect 2317 30719 2375 30725
rect 2317 30716 2329 30719
rect 808 30688 2329 30716
rect 808 30676 814 30688
rect 2317 30685 2329 30688
rect 2363 30685 2375 30719
rect 2317 30679 2375 30685
rect 8386 30676 8392 30728
rect 8444 30716 8450 30728
rect 9861 30719 9919 30725
rect 9861 30716 9873 30719
rect 8444 30688 9873 30716
rect 8444 30676 8450 30688
rect 9861 30685 9873 30688
rect 9907 30685 9919 30719
rect 9861 30679 9919 30685
rect 1486 30648 1492 30660
rect 1447 30620 1492 30648
rect 1486 30608 1492 30620
rect 1544 30608 1550 30660
rect 1673 30651 1731 30657
rect 1673 30617 1685 30651
rect 1719 30648 1731 30651
rect 6454 30648 6460 30660
rect 1719 30620 6460 30648
rect 1719 30617 1731 30620
rect 1673 30611 1731 30617
rect 6454 30608 6460 30620
rect 6512 30608 6518 30660
rect 10042 30580 10048 30592
rect 10003 30552 10048 30580
rect 10042 30540 10048 30552
rect 10100 30540 10106 30592
rect 1104 30490 10856 30512
rect 1104 30438 4214 30490
rect 4266 30438 4278 30490
rect 4330 30438 4342 30490
rect 4394 30438 4406 30490
rect 4458 30438 4470 30490
rect 4522 30438 7478 30490
rect 7530 30438 7542 30490
rect 7594 30438 7606 30490
rect 7658 30438 7670 30490
rect 7722 30438 7734 30490
rect 7786 30438 10856 30490
rect 1104 30416 10856 30438
rect 1854 30240 1860 30252
rect 1815 30212 1860 30240
rect 1854 30200 1860 30212
rect 1912 30200 1918 30252
rect 2501 30243 2559 30249
rect 2501 30209 2513 30243
rect 2547 30240 2559 30243
rect 2590 30240 2596 30252
rect 2547 30212 2596 30240
rect 2547 30209 2559 30212
rect 2501 30203 2559 30209
rect 2590 30200 2596 30212
rect 2648 30200 2654 30252
rect 2041 30175 2099 30181
rect 2041 30141 2053 30175
rect 2087 30172 2099 30175
rect 8662 30172 8668 30184
rect 2087 30144 8668 30172
rect 2087 30141 2099 30144
rect 2041 30135 2099 30141
rect 8662 30132 8668 30144
rect 8720 30132 8726 30184
rect 2685 30107 2743 30113
rect 2685 30073 2697 30107
rect 2731 30104 2743 30107
rect 2774 30104 2780 30116
rect 2731 30076 2780 30104
rect 2731 30073 2743 30076
rect 2685 30067 2743 30073
rect 2774 30064 2780 30076
rect 2832 30064 2838 30116
rect 1104 29946 10856 29968
rect 1104 29894 2582 29946
rect 2634 29894 2646 29946
rect 2698 29894 2710 29946
rect 2762 29894 2774 29946
rect 2826 29894 2838 29946
rect 2890 29894 5846 29946
rect 5898 29894 5910 29946
rect 5962 29894 5974 29946
rect 6026 29894 6038 29946
rect 6090 29894 6102 29946
rect 6154 29894 9110 29946
rect 9162 29894 9174 29946
rect 9226 29894 9238 29946
rect 9290 29894 9302 29946
rect 9354 29894 9366 29946
rect 9418 29894 10856 29946
rect 1104 29872 10856 29894
rect 2869 29835 2927 29841
rect 2869 29801 2881 29835
rect 2915 29832 2927 29835
rect 8386 29832 8392 29844
rect 2915 29804 8392 29832
rect 2915 29801 2927 29804
rect 2869 29795 2927 29801
rect 8386 29792 8392 29804
rect 8444 29792 8450 29844
rect 2038 29764 2044 29776
rect 1999 29736 2044 29764
rect 2038 29724 2044 29736
rect 2096 29724 2102 29776
rect 1394 29588 1400 29640
rect 1452 29628 1458 29640
rect 2038 29628 2044 29640
rect 1452 29600 2044 29628
rect 1452 29588 1458 29600
rect 2038 29588 2044 29600
rect 2096 29588 2102 29640
rect 3053 29631 3111 29637
rect 3053 29597 3065 29631
rect 3099 29628 3111 29631
rect 3234 29628 3240 29640
rect 3099 29600 3240 29628
rect 3099 29597 3111 29600
rect 3053 29591 3111 29597
rect 3234 29588 3240 29600
rect 3292 29588 3298 29640
rect 10134 29628 10140 29640
rect 10095 29600 10140 29628
rect 10134 29588 10140 29600
rect 10192 29588 10198 29640
rect 1486 29520 1492 29572
rect 1544 29560 1550 29572
rect 1857 29563 1915 29569
rect 1857 29560 1869 29563
rect 1544 29532 1869 29560
rect 1544 29520 1550 29532
rect 1857 29529 1869 29532
rect 1903 29529 1915 29563
rect 1857 29523 1915 29529
rect 1104 29402 10856 29424
rect 1104 29350 4214 29402
rect 4266 29350 4278 29402
rect 4330 29350 4342 29402
rect 4394 29350 4406 29402
rect 4458 29350 4470 29402
rect 4522 29350 7478 29402
rect 7530 29350 7542 29402
rect 7594 29350 7606 29402
rect 7658 29350 7670 29402
rect 7722 29350 7734 29402
rect 7786 29350 10856 29402
rect 1104 29328 10856 29350
rect 658 29248 664 29300
rect 716 29288 722 29300
rect 1949 29291 2007 29297
rect 1949 29288 1961 29291
rect 716 29260 1961 29288
rect 716 29248 722 29260
rect 1949 29257 1961 29260
rect 1995 29257 2007 29291
rect 1949 29251 2007 29257
rect 2777 29223 2835 29229
rect 2777 29189 2789 29223
rect 2823 29220 2835 29223
rect 3878 29220 3884 29232
rect 2823 29192 3884 29220
rect 2823 29189 2835 29192
rect 2777 29183 2835 29189
rect 3878 29180 3884 29192
rect 3936 29180 3942 29232
rect 1394 29112 1400 29164
rect 1452 29152 1458 29164
rect 1857 29155 1915 29161
rect 1857 29152 1869 29155
rect 1452 29124 1869 29152
rect 1452 29112 1458 29124
rect 1857 29121 1869 29124
rect 1903 29121 1915 29155
rect 1857 29115 1915 29121
rect 2593 29155 2651 29161
rect 2593 29121 2605 29155
rect 2639 29152 2651 29155
rect 2958 29152 2964 29164
rect 2639 29124 2964 29152
rect 2639 29121 2651 29124
rect 2593 29115 2651 29121
rect 2958 29112 2964 29124
rect 3016 29112 3022 29164
rect 3329 29155 3387 29161
rect 3329 29121 3341 29155
rect 3375 29152 3387 29155
rect 3375 29124 4108 29152
rect 3375 29121 3387 29124
rect 3329 29115 3387 29121
rect 4080 29096 4108 29124
rect 1762 29044 1768 29096
rect 1820 29084 1826 29096
rect 3513 29087 3571 29093
rect 3513 29084 3525 29087
rect 1820 29056 3525 29084
rect 1820 29044 1826 29056
rect 3513 29053 3525 29056
rect 3559 29053 3571 29087
rect 3513 29047 3571 29053
rect 4062 29044 4068 29096
rect 4120 29044 4126 29096
rect 2866 28976 2872 29028
rect 2924 29016 2930 29028
rect 3878 29016 3884 29028
rect 2924 28988 3884 29016
rect 2924 28976 2930 28988
rect 3878 28976 3884 28988
rect 3936 28976 3942 29028
rect 10134 29016 10140 29028
rect 10095 28988 10140 29016
rect 10134 28976 10140 28988
rect 10192 28976 10198 29028
rect 2498 28948 2504 28960
rect 1044 28920 2504 28948
rect 1044 28744 1072 28920
rect 2498 28908 2504 28920
rect 2556 28908 2562 28960
rect 1104 28858 10856 28880
rect 1104 28806 2582 28858
rect 2634 28806 2646 28858
rect 2698 28806 2710 28858
rect 2762 28806 2774 28858
rect 2826 28806 2838 28858
rect 2890 28806 5846 28858
rect 5898 28806 5910 28858
rect 5962 28806 5974 28858
rect 6026 28806 6038 28858
rect 6090 28806 6102 28858
rect 6154 28806 9110 28858
rect 9162 28806 9174 28858
rect 9226 28806 9238 28858
rect 9290 28806 9302 28858
rect 9354 28806 9366 28858
rect 9418 28806 10856 28858
rect 1104 28784 10856 28806
rect 2498 28744 2504 28756
rect 1044 28716 2504 28744
rect 2498 28704 2504 28716
rect 2556 28704 2562 28756
rect 3789 28747 3847 28753
rect 3789 28713 3801 28747
rect 3835 28744 3847 28747
rect 9858 28744 9864 28756
rect 3835 28716 9864 28744
rect 3835 28713 3847 28716
rect 3789 28707 3847 28713
rect 9858 28704 9864 28716
rect 9916 28704 9922 28756
rect 1762 28636 1768 28688
rect 1820 28676 1826 28688
rect 2958 28676 2964 28688
rect 1820 28648 2964 28676
rect 1820 28636 1826 28648
rect 2958 28636 2964 28648
rect 3016 28636 3022 28688
rect 2406 28540 2412 28552
rect 2367 28512 2412 28540
rect 2406 28500 2412 28512
rect 2464 28500 2470 28552
rect 2590 28500 2596 28552
rect 2648 28540 2654 28552
rect 2777 28543 2835 28549
rect 2648 28512 2741 28540
rect 2648 28500 2654 28512
rect 2777 28509 2789 28543
rect 2823 28540 2835 28543
rect 3973 28543 4031 28549
rect 3973 28540 3985 28543
rect 2823 28512 3985 28540
rect 2823 28509 2835 28512
rect 2777 28503 2835 28509
rect 3973 28509 3985 28512
rect 4019 28509 4031 28543
rect 3973 28503 4031 28509
rect 1762 28472 1768 28484
rect 1723 28444 1768 28472
rect 1762 28432 1768 28444
rect 1820 28432 1826 28484
rect 1946 28472 1952 28484
rect 1907 28444 1952 28472
rect 1946 28432 1952 28444
rect 2004 28432 2010 28484
rect 2314 28432 2320 28484
rect 2372 28472 2378 28484
rect 2608 28472 2636 28500
rect 2372 28444 2636 28472
rect 2372 28432 2378 28444
rect 1104 28314 10856 28336
rect 1104 28262 4214 28314
rect 4266 28262 4278 28314
rect 4330 28262 4342 28314
rect 4394 28262 4406 28314
rect 4458 28262 4470 28314
rect 4522 28262 7478 28314
rect 7530 28262 7542 28314
rect 7594 28262 7606 28314
rect 7658 28262 7670 28314
rect 7722 28262 7734 28314
rect 7786 28262 10856 28314
rect 1104 28240 10856 28262
rect 1762 28160 1768 28212
rect 1820 28200 1826 28212
rect 2133 28203 2191 28209
rect 2133 28200 2145 28203
rect 1820 28172 2145 28200
rect 1820 28160 1826 28172
rect 2133 28169 2145 28172
rect 2179 28169 2191 28203
rect 2133 28163 2191 28169
rect 2869 28135 2927 28141
rect 2869 28101 2881 28135
rect 2915 28132 2927 28135
rect 3050 28132 3056 28144
rect 2915 28104 3056 28132
rect 2915 28101 2927 28104
rect 2869 28095 2927 28101
rect 3050 28092 3056 28104
rect 3108 28092 3114 28144
rect 750 28024 756 28076
rect 808 28064 814 28076
rect 1949 28067 2007 28073
rect 1949 28064 1961 28067
rect 808 28036 1961 28064
rect 808 28024 814 28036
rect 1949 28033 1961 28036
rect 1995 28033 2007 28067
rect 1949 28027 2007 28033
rect 2685 28067 2743 28073
rect 2685 28033 2697 28067
rect 2731 28064 2743 28067
rect 2958 28064 2964 28076
rect 2731 28036 2964 28064
rect 2731 28033 2743 28036
rect 2685 28027 2743 28033
rect 2958 28024 2964 28036
rect 3016 28024 3022 28076
rect 1765 27999 1823 28005
rect 1765 27965 1777 27999
rect 1811 27996 1823 27999
rect 3050 27996 3056 28008
rect 1811 27968 3056 27996
rect 1811 27965 1823 27968
rect 1765 27959 1823 27965
rect 3050 27956 3056 27968
rect 3108 27956 3114 28008
rect 9950 27996 9956 28008
rect 9911 27968 9956 27996
rect 9950 27956 9956 27968
rect 10008 27956 10014 28008
rect 1104 27770 10856 27792
rect 1104 27718 2582 27770
rect 2634 27718 2646 27770
rect 2698 27718 2710 27770
rect 2762 27718 2774 27770
rect 2826 27718 2838 27770
rect 2890 27718 5846 27770
rect 5898 27718 5910 27770
rect 5962 27718 5974 27770
rect 6026 27718 6038 27770
rect 6090 27718 6102 27770
rect 6154 27718 9110 27770
rect 9162 27718 9174 27770
rect 9226 27718 9238 27770
rect 9290 27718 9302 27770
rect 9354 27718 9366 27770
rect 9418 27718 10856 27770
rect 1104 27696 10856 27718
rect 1026 27548 1032 27600
rect 1084 27588 1090 27600
rect 2961 27591 3019 27597
rect 2961 27588 2973 27591
rect 1084 27560 2973 27588
rect 1084 27548 1090 27560
rect 2961 27557 2973 27560
rect 3007 27557 3019 27591
rect 2961 27551 3019 27557
rect 1673 27523 1731 27529
rect 1673 27489 1685 27523
rect 1719 27520 1731 27523
rect 3326 27520 3332 27532
rect 1719 27492 3332 27520
rect 1719 27489 1731 27492
rect 1673 27483 1731 27489
rect 3326 27480 3332 27492
rect 3384 27480 3390 27532
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27412 1458 27464
rect 2777 27387 2835 27393
rect 2777 27353 2789 27387
rect 2823 27384 2835 27387
rect 3050 27384 3056 27396
rect 2823 27356 3056 27384
rect 2823 27353 2835 27356
rect 2777 27347 2835 27353
rect 3050 27344 3056 27356
rect 3108 27344 3114 27396
rect 9950 27316 9956 27328
rect 9911 27288 9956 27316
rect 9950 27276 9956 27288
rect 10008 27276 10014 27328
rect 1104 27226 10856 27248
rect 1104 27174 4214 27226
rect 4266 27174 4278 27226
rect 4330 27174 4342 27226
rect 4394 27174 4406 27226
rect 4458 27174 4470 27226
rect 4522 27174 7478 27226
rect 7530 27174 7542 27226
rect 7594 27174 7606 27226
rect 7658 27174 7670 27226
rect 7722 27174 7734 27226
rect 7786 27174 10856 27226
rect 1104 27152 10856 27174
rect 750 27004 756 27056
rect 808 27044 814 27056
rect 3237 27047 3295 27053
rect 808 27016 2360 27044
rect 808 27004 814 27016
rect 1489 26979 1547 26985
rect 1489 26945 1501 26979
rect 1535 26976 1547 26979
rect 2038 26976 2044 26988
rect 1535 26948 2044 26976
rect 1535 26945 1547 26948
rect 1489 26939 1547 26945
rect 2038 26936 2044 26948
rect 2096 26936 2102 26988
rect 2332 26985 2360 27016
rect 3237 27013 3249 27047
rect 3283 27044 3295 27047
rect 4522 27044 4528 27056
rect 3283 27016 4528 27044
rect 3283 27013 3295 27016
rect 3237 27007 3295 27013
rect 4522 27004 4528 27016
rect 4580 27004 4586 27056
rect 2317 26979 2375 26985
rect 2317 26945 2329 26979
rect 2363 26945 2375 26979
rect 2317 26939 2375 26945
rect 2501 26979 2559 26985
rect 2501 26945 2513 26979
rect 2547 26976 2559 26979
rect 3053 26979 3111 26985
rect 3053 26976 3065 26979
rect 2547 26948 3065 26976
rect 2547 26945 2559 26948
rect 2501 26939 2559 26945
rect 3053 26945 3065 26948
rect 3099 26945 3111 26979
rect 3053 26939 3111 26945
rect 2130 26908 2136 26920
rect 2091 26880 2136 26908
rect 2130 26868 2136 26880
rect 2188 26868 2194 26920
rect 1670 26840 1676 26852
rect 1631 26812 1676 26840
rect 1670 26800 1676 26812
rect 1728 26800 1734 26852
rect 10134 26772 10140 26784
rect 10095 26744 10140 26772
rect 10134 26732 10140 26744
rect 10192 26732 10198 26784
rect 1104 26682 10856 26704
rect 1104 26630 2582 26682
rect 2634 26630 2646 26682
rect 2698 26630 2710 26682
rect 2762 26630 2774 26682
rect 2826 26630 2838 26682
rect 2890 26630 5846 26682
rect 5898 26630 5910 26682
rect 5962 26630 5974 26682
rect 6026 26630 6038 26682
rect 6090 26630 6102 26682
rect 6154 26630 9110 26682
rect 9162 26630 9174 26682
rect 9226 26630 9238 26682
rect 9290 26630 9302 26682
rect 9354 26630 9366 26682
rect 9418 26630 10856 26682
rect 1104 26608 10856 26630
rect 2038 26568 2044 26580
rect 1999 26540 2044 26568
rect 2038 26528 2044 26540
rect 2096 26528 2102 26580
rect 1670 26460 1676 26512
rect 1728 26500 1734 26512
rect 2130 26500 2136 26512
rect 1728 26472 2136 26500
rect 1728 26460 1734 26472
rect 2130 26460 2136 26472
rect 2188 26460 2194 26512
rect 2777 26503 2835 26509
rect 2777 26469 2789 26503
rect 2823 26500 2835 26503
rect 3142 26500 3148 26512
rect 2823 26472 3148 26500
rect 2823 26469 2835 26472
rect 2777 26463 2835 26469
rect 3142 26460 3148 26472
rect 3200 26460 3206 26512
rect 750 26392 756 26444
rect 808 26432 814 26444
rect 808 26404 1900 26432
rect 808 26392 814 26404
rect 934 26324 940 26376
rect 992 26364 998 26376
rect 1486 26364 1492 26376
rect 992 26336 1492 26364
rect 992 26324 998 26336
rect 1486 26324 1492 26336
rect 1544 26364 1550 26376
rect 1872 26373 1900 26404
rect 1673 26367 1731 26373
rect 1673 26364 1685 26367
rect 1544 26336 1685 26364
rect 1544 26324 1550 26336
rect 1673 26333 1685 26336
rect 1719 26333 1731 26367
rect 1673 26327 1731 26333
rect 1857 26367 1915 26373
rect 1857 26333 1869 26367
rect 1903 26333 1915 26367
rect 1857 26327 1915 26333
rect 2590 26296 2596 26308
rect 2551 26268 2596 26296
rect 2590 26256 2596 26268
rect 2648 26256 2654 26308
rect 3050 26188 3056 26240
rect 3108 26228 3114 26240
rect 3326 26228 3332 26240
rect 3108 26200 3332 26228
rect 3108 26188 3114 26200
rect 3326 26188 3332 26200
rect 3384 26188 3390 26240
rect 1104 26138 10856 26160
rect 1104 26086 4214 26138
rect 4266 26086 4278 26138
rect 4330 26086 4342 26138
rect 4394 26086 4406 26138
rect 4458 26086 4470 26138
rect 4522 26086 7478 26138
rect 7530 26086 7542 26138
rect 7594 26086 7606 26138
rect 7658 26086 7670 26138
rect 7722 26086 7734 26138
rect 7786 26086 10856 26138
rect 1104 26064 10856 26086
rect 14 25984 20 26036
rect 72 26024 78 26036
rect 1949 26027 2007 26033
rect 1949 26024 1961 26027
rect 72 25996 1961 26024
rect 72 25984 78 25996
rect 1949 25993 1961 25996
rect 1995 25993 2007 26027
rect 3418 26024 3424 26036
rect 3379 25996 3424 26024
rect 1949 25987 2007 25993
rect 3418 25984 3424 25996
rect 3476 25984 3482 26036
rect 2777 25959 2835 25965
rect 2777 25925 2789 25959
rect 2823 25956 2835 25959
rect 3602 25956 3608 25968
rect 2823 25928 3608 25956
rect 2823 25925 2835 25928
rect 2777 25919 2835 25925
rect 3602 25916 3608 25928
rect 3660 25916 3666 25968
rect 1857 25891 1915 25897
rect 1857 25857 1869 25891
rect 1903 25888 1915 25891
rect 2038 25888 2044 25900
rect 1903 25860 2044 25888
rect 1903 25857 1915 25860
rect 1857 25851 1915 25857
rect 2038 25848 2044 25860
rect 2096 25848 2102 25900
rect 2593 25891 2651 25897
rect 2593 25857 2605 25891
rect 2639 25888 2651 25891
rect 2958 25888 2964 25900
rect 2639 25860 2964 25888
rect 2639 25857 2651 25860
rect 2593 25851 2651 25857
rect 2958 25848 2964 25860
rect 3016 25848 3022 25900
rect 3326 25888 3332 25900
rect 3287 25860 3332 25888
rect 3326 25848 3332 25860
rect 3384 25848 3390 25900
rect 10134 25684 10140 25696
rect 10095 25656 10140 25684
rect 10134 25644 10140 25656
rect 10192 25644 10198 25696
rect 1104 25594 10856 25616
rect 1104 25542 2582 25594
rect 2634 25542 2646 25594
rect 2698 25542 2710 25594
rect 2762 25542 2774 25594
rect 2826 25542 2838 25594
rect 2890 25542 5846 25594
rect 5898 25542 5910 25594
rect 5962 25542 5974 25594
rect 6026 25542 6038 25594
rect 6090 25542 6102 25594
rect 6154 25542 9110 25594
rect 9162 25542 9174 25594
rect 9226 25542 9238 25594
rect 9290 25542 9302 25594
rect 9354 25542 9366 25594
rect 9418 25542 10856 25594
rect 1104 25520 10856 25542
rect 1854 25440 1860 25492
rect 1912 25480 1918 25492
rect 1949 25483 2007 25489
rect 1949 25480 1961 25483
rect 1912 25452 1961 25480
rect 1912 25440 1918 25452
rect 1949 25449 1961 25452
rect 1995 25449 2007 25483
rect 1949 25443 2007 25449
rect 3786 25440 3792 25492
rect 3844 25480 3850 25492
rect 3973 25483 4031 25489
rect 3973 25480 3985 25483
rect 3844 25452 3985 25480
rect 3844 25440 3850 25452
rect 3973 25449 3985 25452
rect 4019 25449 4031 25483
rect 3973 25443 4031 25449
rect 2777 25415 2835 25421
rect 2777 25381 2789 25415
rect 2823 25412 2835 25415
rect 3050 25412 3056 25424
rect 2823 25384 3056 25412
rect 2823 25381 2835 25384
rect 2777 25375 2835 25381
rect 3050 25372 3056 25384
rect 3108 25372 3114 25424
rect 10134 25276 10140 25288
rect 10095 25248 10140 25276
rect 10134 25236 10140 25248
rect 10192 25236 10198 25288
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 2593 25211 2651 25217
rect 2593 25177 2605 25211
rect 2639 25208 2651 25211
rect 3878 25208 3884 25220
rect 2639 25180 2774 25208
rect 3839 25180 3884 25208
rect 2639 25177 2651 25180
rect 2593 25171 2651 25177
rect 2746 25140 2774 25180
rect 3878 25168 3884 25180
rect 3936 25168 3942 25220
rect 2866 25140 2872 25152
rect 2746 25112 2872 25140
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 1104 25050 10856 25072
rect 1104 24998 4214 25050
rect 4266 24998 4278 25050
rect 4330 24998 4342 25050
rect 4394 24998 4406 25050
rect 4458 24998 4470 25050
rect 4522 24998 7478 25050
rect 7530 24998 7542 25050
rect 7594 24998 7606 25050
rect 7658 24998 7670 25050
rect 7722 24998 7734 25050
rect 7786 24998 10856 25050
rect 1104 24976 10856 24998
rect 2314 24828 2320 24880
rect 2372 24868 2378 24880
rect 2372 24840 2636 24868
rect 2372 24828 2378 24840
rect 2608 24809 2636 24840
rect 1765 24803 1823 24809
rect 1765 24769 1777 24803
rect 1811 24800 1823 24803
rect 2593 24803 2651 24809
rect 1811 24772 2544 24800
rect 1811 24769 1823 24772
rect 1765 24763 1823 24769
rect 1118 24692 1124 24744
rect 1176 24732 1182 24744
rect 1949 24735 2007 24741
rect 1949 24732 1961 24735
rect 1176 24704 1961 24732
rect 1176 24692 1182 24704
rect 1949 24701 1961 24704
rect 1995 24701 2007 24735
rect 1949 24695 2007 24701
rect 2130 24692 2136 24744
rect 2188 24732 2194 24744
rect 2409 24735 2467 24741
rect 2409 24732 2421 24735
rect 2188 24704 2421 24732
rect 2188 24692 2194 24704
rect 2409 24701 2421 24704
rect 2455 24701 2467 24735
rect 2516 24732 2544 24772
rect 2593 24769 2605 24803
rect 2639 24800 2651 24803
rect 2958 24800 2964 24812
rect 2639 24772 2964 24800
rect 2639 24769 2651 24772
rect 2593 24763 2651 24769
rect 2958 24760 2964 24772
rect 3016 24760 3022 24812
rect 3234 24732 3240 24744
rect 2516 24704 3240 24732
rect 2409 24695 2467 24701
rect 3234 24692 3240 24704
rect 3292 24692 3298 24744
rect 2777 24599 2835 24605
rect 2777 24565 2789 24599
rect 2823 24596 2835 24599
rect 3786 24596 3792 24608
rect 2823 24568 3792 24596
rect 2823 24565 2835 24568
rect 2777 24559 2835 24565
rect 3786 24556 3792 24568
rect 3844 24556 3850 24608
rect 1104 24506 10856 24528
rect 1104 24454 2582 24506
rect 2634 24454 2646 24506
rect 2698 24454 2710 24506
rect 2762 24454 2774 24506
rect 2826 24454 2838 24506
rect 2890 24454 5846 24506
rect 5898 24454 5910 24506
rect 5962 24454 5974 24506
rect 6026 24454 6038 24506
rect 6090 24454 6102 24506
rect 6154 24454 9110 24506
rect 9162 24454 9174 24506
rect 9226 24454 9238 24506
rect 9290 24454 9302 24506
rect 9354 24454 9366 24506
rect 9418 24454 10856 24506
rect 1104 24432 10856 24454
rect 2041 24327 2099 24333
rect 2041 24293 2053 24327
rect 2087 24324 2099 24327
rect 2222 24324 2228 24336
rect 2087 24296 2228 24324
rect 2087 24293 2099 24296
rect 2041 24287 2099 24293
rect 2222 24284 2228 24296
rect 2280 24284 2286 24336
rect 3786 24256 3792 24268
rect 3747 24228 3792 24256
rect 3786 24216 3792 24228
rect 3844 24216 3850 24268
rect 4065 24259 4123 24265
rect 4065 24225 4077 24259
rect 4111 24256 4123 24259
rect 7834 24256 7840 24268
rect 4111 24228 7840 24256
rect 4111 24225 4123 24228
rect 4065 24219 4123 24225
rect 7834 24216 7840 24228
rect 7892 24216 7898 24268
rect 2682 24188 2688 24200
rect 2643 24160 2688 24188
rect 2682 24148 2688 24160
rect 2740 24148 2746 24200
rect 2777 24191 2835 24197
rect 2777 24157 2789 24191
rect 2823 24188 2835 24191
rect 2958 24188 2964 24200
rect 2823 24160 2964 24188
rect 2823 24157 2835 24160
rect 2777 24151 2835 24157
rect 2958 24148 2964 24160
rect 3016 24148 3022 24200
rect 10134 24188 10140 24200
rect 10095 24160 10140 24188
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 1857 24123 1915 24129
rect 1857 24089 1869 24123
rect 1903 24120 1915 24123
rect 3050 24120 3056 24132
rect 1903 24092 3056 24120
rect 1903 24089 1915 24092
rect 1857 24083 1915 24089
rect 3050 24080 3056 24092
rect 3108 24080 3114 24132
rect 2961 24055 3019 24061
rect 2961 24021 2973 24055
rect 3007 24052 3019 24055
rect 3786 24052 3792 24064
rect 3007 24024 3792 24052
rect 3007 24021 3019 24024
rect 2961 24015 3019 24021
rect 3786 24012 3792 24024
rect 3844 24012 3850 24064
rect 1104 23962 10856 23984
rect 1104 23910 4214 23962
rect 4266 23910 4278 23962
rect 4330 23910 4342 23962
rect 4394 23910 4406 23962
rect 4458 23910 4470 23962
rect 4522 23910 7478 23962
rect 7530 23910 7542 23962
rect 7594 23910 7606 23962
rect 7658 23910 7670 23962
rect 7722 23910 7734 23962
rect 7786 23910 10856 23962
rect 1104 23888 10856 23910
rect 3050 23848 3056 23860
rect 3011 23820 3056 23848
rect 3050 23808 3056 23820
rect 3108 23808 3114 23860
rect 3970 23808 3976 23860
rect 4028 23808 4034 23860
rect 5074 23848 5080 23860
rect 5035 23820 5080 23848
rect 5074 23808 5080 23820
rect 5132 23808 5138 23860
rect 5258 23808 5264 23860
rect 5316 23808 5322 23860
rect 750 23740 756 23792
rect 808 23780 814 23792
rect 808 23752 2912 23780
rect 808 23740 814 23752
rect 1578 23672 1584 23724
rect 1636 23712 1642 23724
rect 2884 23721 2912 23752
rect 1673 23715 1731 23721
rect 1673 23712 1685 23715
rect 1636 23684 1685 23712
rect 1636 23672 1642 23684
rect 1673 23681 1685 23684
rect 1719 23681 1731 23715
rect 1673 23675 1731 23681
rect 2869 23715 2927 23721
rect 2869 23681 2881 23715
rect 2915 23712 2927 23715
rect 3050 23712 3056 23724
rect 2915 23684 3056 23712
rect 2915 23681 2927 23684
rect 2869 23675 2927 23681
rect 3050 23672 3056 23684
rect 3108 23672 3114 23724
rect 3786 23712 3792 23724
rect 3747 23684 3792 23712
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 1118 23604 1124 23656
rect 1176 23644 1182 23656
rect 1397 23647 1455 23653
rect 1397 23644 1409 23647
rect 1176 23616 1409 23644
rect 1176 23604 1182 23616
rect 1397 23613 1409 23616
rect 1443 23613 1455 23647
rect 1397 23607 1455 23613
rect 2685 23647 2743 23653
rect 2685 23613 2697 23647
rect 2731 23644 2743 23647
rect 2774 23644 2780 23656
rect 2731 23616 2780 23644
rect 2731 23613 2743 23616
rect 2685 23607 2743 23613
rect 2774 23604 2780 23616
rect 2832 23644 2838 23656
rect 3326 23644 3332 23656
rect 2832 23616 3332 23644
rect 2832 23604 2838 23616
rect 3326 23604 3332 23616
rect 3384 23604 3390 23656
rect 3786 23536 3792 23588
rect 3844 23576 3850 23588
rect 3988 23576 4016 23808
rect 4522 23740 4528 23792
rect 4580 23780 4586 23792
rect 5276 23780 5304 23808
rect 4580 23752 5304 23780
rect 4580 23740 4586 23752
rect 4890 23672 4896 23724
rect 4948 23712 4954 23724
rect 5074 23712 5080 23724
rect 4948 23684 5080 23712
rect 4948 23672 4954 23684
rect 5074 23672 5080 23684
rect 5132 23672 5138 23724
rect 5258 23712 5264 23724
rect 5219 23684 5264 23712
rect 5258 23672 5264 23684
rect 5316 23672 5322 23724
rect 4065 23647 4123 23653
rect 4065 23613 4077 23647
rect 4111 23644 4123 23647
rect 7926 23644 7932 23656
rect 4111 23616 7932 23644
rect 4111 23613 4123 23616
rect 4065 23607 4123 23613
rect 7926 23604 7932 23616
rect 7984 23604 7990 23656
rect 3844 23548 4016 23576
rect 3844 23536 3850 23548
rect 3234 23468 3240 23520
rect 3292 23508 3298 23520
rect 4062 23508 4068 23520
rect 3292 23480 4068 23508
rect 3292 23468 3298 23480
rect 4062 23468 4068 23480
rect 4120 23468 4126 23520
rect 10134 23508 10140 23520
rect 10095 23480 10140 23508
rect 10134 23468 10140 23480
rect 10192 23468 10198 23520
rect 1104 23418 10856 23440
rect 1104 23366 2582 23418
rect 2634 23366 2646 23418
rect 2698 23366 2710 23418
rect 2762 23366 2774 23418
rect 2826 23366 2838 23418
rect 2890 23366 5846 23418
rect 5898 23366 5910 23418
rect 5962 23366 5974 23418
rect 6026 23366 6038 23418
rect 6090 23366 6102 23418
rect 6154 23366 9110 23418
rect 9162 23366 9174 23418
rect 9226 23366 9238 23418
rect 9290 23366 9302 23418
rect 9354 23366 9366 23418
rect 9418 23366 10856 23418
rect 1104 23344 10856 23366
rect 4154 23264 4160 23316
rect 4212 23304 4218 23316
rect 4341 23307 4399 23313
rect 4341 23304 4353 23307
rect 4212 23276 4353 23304
rect 4212 23264 4218 23276
rect 4341 23273 4353 23276
rect 4387 23273 4399 23307
rect 4341 23267 4399 23273
rect 4982 23264 4988 23316
rect 5040 23304 5046 23316
rect 5077 23307 5135 23313
rect 5077 23304 5089 23307
rect 5040 23276 5089 23304
rect 5040 23264 5046 23276
rect 5077 23273 5089 23276
rect 5123 23273 5135 23307
rect 5077 23267 5135 23273
rect 5718 23236 5724 23248
rect 1688 23208 5724 23236
rect 1688 23177 1716 23208
rect 5718 23196 5724 23208
rect 5776 23196 5782 23248
rect 1673 23171 1731 23177
rect 1673 23137 1685 23171
rect 1719 23137 1731 23171
rect 1673 23131 1731 23137
rect 3050 23128 3056 23180
rect 3108 23128 3114 23180
rect 1394 23100 1400 23112
rect 1355 23072 1400 23100
rect 1394 23060 1400 23072
rect 1452 23060 1458 23112
rect 2130 23060 2136 23112
rect 2188 23100 2194 23112
rect 2685 23103 2743 23109
rect 2685 23100 2697 23103
rect 2188 23072 2697 23100
rect 2188 23060 2194 23072
rect 2685 23069 2697 23072
rect 2731 23069 2743 23103
rect 2685 23063 2743 23069
rect 2869 23103 2927 23109
rect 2869 23069 2881 23103
rect 2915 23100 2927 23103
rect 3068 23100 3096 23128
rect 2915 23072 3096 23100
rect 2915 23069 2927 23072
rect 2869 23063 2927 23069
rect 3878 23060 3884 23112
rect 3936 23100 3942 23112
rect 4985 23103 5043 23109
rect 4985 23100 4997 23103
rect 3936 23072 4997 23100
rect 3936 23060 3942 23072
rect 4985 23069 4997 23072
rect 5031 23069 5043 23103
rect 4985 23063 5043 23069
rect 3053 23035 3111 23041
rect 3053 23001 3065 23035
rect 3099 23032 3111 23035
rect 4249 23035 4307 23041
rect 4249 23032 4261 23035
rect 3099 23004 4261 23032
rect 3099 23001 3111 23004
rect 3053 22995 3111 23001
rect 4249 23001 4261 23004
rect 4295 23001 4307 23035
rect 4249 22995 4307 23001
rect 4522 22992 4528 23044
rect 4580 23032 4586 23044
rect 4580 23004 4752 23032
rect 4580 22992 4586 23004
rect 4724 22976 4752 23004
rect 1762 22924 1768 22976
rect 1820 22964 1826 22976
rect 2314 22964 2320 22976
rect 1820 22936 2320 22964
rect 1820 22924 1826 22936
rect 2314 22924 2320 22936
rect 2372 22924 2378 22976
rect 4706 22924 4712 22976
rect 4764 22924 4770 22976
rect 1104 22874 10856 22896
rect 1104 22822 4214 22874
rect 4266 22822 4278 22874
rect 4330 22822 4342 22874
rect 4394 22822 4406 22874
rect 4458 22822 4470 22874
rect 4522 22822 7478 22874
rect 7530 22822 7542 22874
rect 7594 22822 7606 22874
rect 7658 22822 7670 22874
rect 7722 22822 7734 22874
rect 7786 22822 10856 22874
rect 1104 22800 10856 22822
rect 3050 22760 3056 22772
rect 1872 22732 3056 22760
rect 1872 22633 1900 22732
rect 3050 22720 3056 22732
rect 3108 22760 3114 22772
rect 3234 22760 3240 22772
rect 3108 22732 3240 22760
rect 3108 22720 3114 22732
rect 3234 22720 3240 22732
rect 3292 22720 3298 22772
rect 3510 22720 3516 22772
rect 3568 22760 3574 22772
rect 3605 22763 3663 22769
rect 3605 22760 3617 22763
rect 3568 22732 3617 22760
rect 3568 22720 3574 22732
rect 3605 22729 3617 22732
rect 3651 22729 3663 22763
rect 3605 22723 3663 22729
rect 2961 22695 3019 22701
rect 2961 22661 2973 22695
rect 3007 22692 3019 22695
rect 5258 22692 5264 22704
rect 3007 22664 5264 22692
rect 3007 22661 3019 22664
rect 2961 22655 3019 22661
rect 5258 22652 5264 22664
rect 5316 22652 5322 22704
rect 1857 22627 1915 22633
rect 1857 22593 1869 22627
rect 1903 22593 1915 22627
rect 1857 22587 1915 22593
rect 2777 22627 2835 22633
rect 2777 22593 2789 22627
rect 2823 22593 2835 22627
rect 3510 22624 3516 22636
rect 3471 22596 3516 22624
rect 2777 22587 2835 22593
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22556 1731 22559
rect 2314 22556 2320 22568
rect 1719 22528 2320 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 2314 22516 2320 22528
rect 2372 22556 2378 22568
rect 2593 22559 2651 22565
rect 2593 22556 2605 22559
rect 2372 22528 2605 22556
rect 2372 22516 2378 22528
rect 2593 22525 2605 22528
rect 2639 22525 2651 22559
rect 2792 22556 2820 22587
rect 3510 22584 3516 22596
rect 3568 22584 3574 22636
rect 2958 22556 2964 22568
rect 2792 22528 2964 22556
rect 2593 22519 2651 22525
rect 2958 22516 2964 22528
rect 3016 22516 3022 22568
rect 2041 22491 2099 22497
rect 2041 22457 2053 22491
rect 2087 22488 2099 22491
rect 3050 22488 3056 22500
rect 2087 22460 3056 22488
rect 2087 22457 2099 22460
rect 2041 22451 2099 22457
rect 3050 22448 3056 22460
rect 3108 22448 3114 22500
rect 10134 22488 10140 22500
rect 10095 22460 10140 22488
rect 10134 22448 10140 22460
rect 10192 22448 10198 22500
rect 3142 22380 3148 22432
rect 3200 22420 3206 22432
rect 3970 22420 3976 22432
rect 3200 22392 3976 22420
rect 3200 22380 3206 22392
rect 3970 22380 3976 22392
rect 4028 22380 4034 22432
rect 1104 22330 10856 22352
rect 1104 22278 2582 22330
rect 2634 22278 2646 22330
rect 2698 22278 2710 22330
rect 2762 22278 2774 22330
rect 2826 22278 2838 22330
rect 2890 22278 5846 22330
rect 5898 22278 5910 22330
rect 5962 22278 5974 22330
rect 6026 22278 6038 22330
rect 6090 22278 6102 22330
rect 6154 22278 9110 22330
rect 9162 22278 9174 22330
rect 9226 22278 9238 22330
rect 9290 22278 9302 22330
rect 9354 22278 9366 22330
rect 9418 22278 10856 22330
rect 1104 22256 10856 22278
rect 2314 22216 2320 22228
rect 2240 22188 2320 22216
rect 2240 22160 2268 22188
rect 2314 22176 2320 22188
rect 2372 22176 2378 22228
rect 3142 22176 3148 22228
rect 3200 22216 3206 22228
rect 3602 22216 3608 22228
rect 3200 22188 3608 22216
rect 3200 22176 3206 22188
rect 3602 22176 3608 22188
rect 3660 22176 3666 22228
rect 2222 22108 2228 22160
rect 2280 22108 2286 22160
rect 10134 22148 10140 22160
rect 10095 22120 10140 22148
rect 10134 22108 10140 22120
rect 10192 22108 10198 22160
rect 1673 22083 1731 22089
rect 1673 22049 1685 22083
rect 1719 22080 1731 22083
rect 1946 22080 1952 22092
rect 1719 22052 1952 22080
rect 1719 22049 1731 22052
rect 1673 22043 1731 22049
rect 1946 22040 1952 22052
rect 2004 22040 2010 22092
rect 2130 22040 2136 22092
rect 2188 22080 2194 22092
rect 2314 22080 2320 22092
rect 2188 22052 2320 22080
rect 2188 22040 2194 22052
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 2961 22083 3019 22089
rect 2961 22049 2973 22083
rect 3007 22080 3019 22083
rect 5074 22080 5080 22092
rect 3007 22052 5080 22080
rect 3007 22049 3019 22052
rect 2961 22043 3019 22049
rect 5074 22040 5080 22052
rect 5132 22040 5138 22092
rect 1394 22012 1400 22024
rect 1355 21984 1400 22012
rect 1394 21972 1400 21984
rect 1452 21972 1458 22024
rect 2777 22015 2835 22021
rect 2777 21981 2789 22015
rect 2823 22012 2835 22015
rect 3050 22012 3056 22024
rect 2823 21984 3056 22012
rect 2823 21981 2835 21984
rect 2777 21975 2835 21981
rect 3050 21972 3056 21984
rect 3108 21972 3114 22024
rect 1104 21786 10856 21808
rect 1104 21734 4214 21786
rect 4266 21734 4278 21786
rect 4330 21734 4342 21786
rect 4394 21734 4406 21786
rect 4458 21734 4470 21786
rect 4522 21734 7478 21786
rect 7530 21734 7542 21786
rect 7594 21734 7606 21786
rect 7658 21734 7670 21786
rect 7722 21734 7734 21786
rect 7786 21734 10856 21786
rect 1104 21712 10856 21734
rect 2869 21675 2927 21681
rect 2869 21641 2881 21675
rect 2915 21672 2927 21675
rect 4798 21672 4804 21684
rect 2915 21644 4804 21672
rect 2915 21641 2927 21644
rect 2869 21635 2927 21641
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 3697 21607 3755 21613
rect 3697 21573 3709 21607
rect 3743 21604 3755 21607
rect 5442 21604 5448 21616
rect 3743 21576 5448 21604
rect 3743 21573 3755 21576
rect 3697 21567 3755 21573
rect 5442 21564 5448 21576
rect 5500 21564 5506 21616
rect 2777 21539 2835 21545
rect 2777 21505 2789 21539
rect 2823 21536 2835 21539
rect 3050 21536 3056 21548
rect 2823 21508 3056 21536
rect 2823 21505 2835 21508
rect 2777 21499 2835 21505
rect 3050 21496 3056 21508
rect 3108 21496 3114 21548
rect 3513 21539 3571 21545
rect 3513 21505 3525 21539
rect 3559 21536 3571 21539
rect 4798 21536 4804 21548
rect 3559 21508 4804 21536
rect 3559 21505 3571 21508
rect 3513 21499 3571 21505
rect 4798 21496 4804 21508
rect 4856 21496 4862 21548
rect 1394 21468 1400 21480
rect 1355 21440 1400 21468
rect 1394 21428 1400 21440
rect 1452 21428 1458 21480
rect 1673 21471 1731 21477
rect 1673 21437 1685 21471
rect 1719 21468 1731 21471
rect 3970 21468 3976 21480
rect 1719 21440 3976 21468
rect 1719 21437 1731 21440
rect 1673 21431 1731 21437
rect 3970 21428 3976 21440
rect 4028 21428 4034 21480
rect 10134 21332 10140 21344
rect 10095 21304 10140 21332
rect 10134 21292 10140 21304
rect 10192 21292 10198 21344
rect 1104 21242 10856 21264
rect 1104 21190 2582 21242
rect 2634 21190 2646 21242
rect 2698 21190 2710 21242
rect 2762 21190 2774 21242
rect 2826 21190 2838 21242
rect 2890 21190 5846 21242
rect 5898 21190 5910 21242
rect 5962 21190 5974 21242
rect 6026 21190 6038 21242
rect 6090 21190 6102 21242
rect 6154 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 9238 21242
rect 9290 21190 9302 21242
rect 9354 21190 9366 21242
rect 9418 21190 10856 21242
rect 1104 21168 10856 21190
rect 3053 21131 3111 21137
rect 3053 21097 3065 21131
rect 3099 21128 3111 21131
rect 3418 21128 3424 21140
rect 3099 21100 3424 21128
rect 3099 21097 3111 21100
rect 3053 21091 3111 21097
rect 3418 21088 3424 21100
rect 3476 21088 3482 21140
rect 1026 21020 1032 21072
rect 1084 21060 1090 21072
rect 1084 21032 1716 21060
rect 1084 21020 1090 21032
rect 1210 20952 1216 21004
rect 1268 20992 1274 21004
rect 1688 21001 1716 21032
rect 1397 20995 1455 21001
rect 1397 20992 1409 20995
rect 1268 20964 1409 20992
rect 1268 20952 1274 20964
rect 1397 20961 1409 20964
rect 1443 20961 1455 20995
rect 1397 20955 1455 20961
rect 1673 20995 1731 21001
rect 1673 20961 1685 20995
rect 1719 20961 1731 20995
rect 1673 20955 1731 20961
rect 1946 20884 1952 20936
rect 2004 20924 2010 20936
rect 2685 20927 2743 20933
rect 2685 20924 2697 20927
rect 2004 20896 2697 20924
rect 2004 20884 2010 20896
rect 2685 20893 2697 20896
rect 2731 20893 2743 20927
rect 2685 20887 2743 20893
rect 2869 20927 2927 20933
rect 2869 20893 2881 20927
rect 2915 20924 2927 20927
rect 2958 20924 2964 20936
rect 2915 20896 2964 20924
rect 2915 20893 2927 20896
rect 2869 20887 2927 20893
rect 2958 20884 2964 20896
rect 3016 20924 3022 20936
rect 3418 20924 3424 20936
rect 3016 20896 3424 20924
rect 3016 20884 3022 20896
rect 3418 20884 3424 20896
rect 3476 20884 3482 20936
rect 1104 20698 10856 20720
rect 1104 20646 4214 20698
rect 4266 20646 4278 20698
rect 4330 20646 4342 20698
rect 4394 20646 4406 20698
rect 4458 20646 4470 20698
rect 4522 20646 7478 20698
rect 7530 20646 7542 20698
rect 7594 20646 7606 20698
rect 7658 20646 7670 20698
rect 7722 20646 7734 20698
rect 7786 20646 10856 20698
rect 1104 20624 10856 20646
rect 1670 20448 1676 20460
rect 1631 20420 1676 20448
rect 1670 20408 1676 20420
rect 1728 20408 1734 20460
rect 2685 20451 2743 20457
rect 2685 20417 2697 20451
rect 2731 20448 2743 20451
rect 2774 20448 2780 20460
rect 2731 20420 2780 20448
rect 2731 20417 2743 20420
rect 2685 20411 2743 20417
rect 2774 20408 2780 20420
rect 2832 20408 2838 20460
rect 2961 20451 3019 20457
rect 2961 20417 2973 20451
rect 3007 20448 3019 20451
rect 3142 20448 3148 20460
rect 3007 20420 3148 20448
rect 3007 20417 3019 20420
rect 2961 20411 3019 20417
rect 3142 20408 3148 20420
rect 3200 20408 3206 20460
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20448 9919 20451
rect 10134 20448 10140 20460
rect 9907 20420 10140 20448
rect 9907 20417 9919 20420
rect 9861 20411 9919 20417
rect 10134 20408 10140 20420
rect 10192 20408 10198 20460
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 10042 20312 10048 20324
rect 10003 20284 10048 20312
rect 10042 20272 10048 20284
rect 10100 20272 10106 20324
rect 1104 20154 10856 20176
rect 1104 20102 2582 20154
rect 2634 20102 2646 20154
rect 2698 20102 2710 20154
rect 2762 20102 2774 20154
rect 2826 20102 2838 20154
rect 2890 20102 5846 20154
rect 5898 20102 5910 20154
rect 5962 20102 5974 20154
rect 6026 20102 6038 20154
rect 6090 20102 6102 20154
rect 6154 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 9238 20154
rect 9290 20102 9302 20154
rect 9354 20102 9366 20154
rect 9418 20102 10856 20154
rect 1104 20080 10856 20102
rect 3050 20040 3056 20052
rect 3011 20012 3056 20040
rect 3050 20000 3056 20012
rect 3108 20000 3114 20052
rect 1578 19864 1584 19916
rect 1636 19904 1642 19916
rect 1673 19907 1731 19913
rect 1673 19904 1685 19907
rect 1636 19876 1685 19904
rect 1636 19864 1642 19876
rect 1673 19873 1685 19876
rect 1719 19873 1731 19907
rect 1673 19867 1731 19873
rect 1762 19864 1768 19916
rect 1820 19904 1826 19916
rect 2130 19904 2136 19916
rect 1820 19876 2136 19904
rect 1820 19864 1826 19876
rect 2130 19864 2136 19876
rect 2188 19904 2194 19916
rect 2685 19907 2743 19913
rect 2685 19904 2697 19907
rect 2188 19876 2697 19904
rect 2188 19864 2194 19876
rect 2685 19873 2697 19876
rect 2731 19873 2743 19907
rect 2685 19867 2743 19873
rect 1394 19836 1400 19848
rect 1355 19808 1400 19836
rect 1394 19796 1400 19808
rect 1452 19796 1458 19848
rect 2869 19839 2927 19845
rect 2869 19805 2881 19839
rect 2915 19836 2927 19839
rect 3234 19836 3240 19848
rect 2915 19808 3240 19836
rect 2915 19805 2927 19808
rect 2869 19799 2927 19805
rect 3234 19796 3240 19808
rect 3292 19796 3298 19848
rect 9214 19796 9220 19848
rect 9272 19836 9278 19848
rect 9861 19839 9919 19845
rect 9861 19836 9873 19839
rect 9272 19808 9873 19836
rect 9272 19796 9278 19808
rect 9861 19805 9873 19808
rect 9907 19805 9919 19839
rect 9861 19799 9919 19805
rect 10042 19700 10048 19712
rect 10003 19672 10048 19700
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 1104 19610 10856 19632
rect 1104 19558 4214 19610
rect 4266 19558 4278 19610
rect 4330 19558 4342 19610
rect 4394 19558 4406 19610
rect 4458 19558 4470 19610
rect 4522 19558 7478 19610
rect 7530 19558 7542 19610
rect 7594 19558 7606 19610
rect 7658 19558 7670 19610
rect 7722 19558 7734 19610
rect 7786 19558 10856 19610
rect 1104 19536 10856 19558
rect 9214 19496 9220 19508
rect 9175 19468 9220 19496
rect 9214 19456 9220 19468
rect 9272 19456 9278 19508
rect 3602 19388 3608 19440
rect 3660 19428 3666 19440
rect 3660 19400 10088 19428
rect 3660 19388 3666 19400
rect 1486 19320 1492 19372
rect 1544 19360 1550 19372
rect 1673 19363 1731 19369
rect 1673 19360 1685 19363
rect 1544 19332 1685 19360
rect 1544 19320 1550 19332
rect 1673 19329 1685 19332
rect 1719 19329 1731 19363
rect 1673 19323 1731 19329
rect 2777 19363 2835 19369
rect 2777 19329 2789 19363
rect 2823 19360 2835 19363
rect 2958 19360 2964 19372
rect 2823 19332 2964 19360
rect 2823 19329 2835 19332
rect 2777 19323 2835 19329
rect 2958 19320 2964 19332
rect 3016 19320 3022 19372
rect 3510 19320 3516 19372
rect 3568 19360 3574 19372
rect 10060 19369 10088 19400
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 3568 19332 9413 19360
rect 3568 19320 3574 19332
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 9401 19323 9459 19329
rect 10045 19363 10103 19369
rect 10045 19329 10057 19363
rect 10091 19329 10103 19363
rect 10045 19323 10103 19329
rect 1394 19292 1400 19304
rect 1355 19264 1400 19292
rect 1394 19252 1400 19264
rect 1452 19252 1458 19304
rect 2961 19227 3019 19233
rect 2961 19193 2973 19227
rect 3007 19224 3019 19227
rect 5166 19224 5172 19236
rect 3007 19196 5172 19224
rect 3007 19193 3019 19196
rect 2961 19187 3019 19193
rect 5166 19184 5172 19196
rect 5224 19184 5230 19236
rect 9858 19156 9864 19168
rect 9819 19128 9864 19156
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 1104 19066 10856 19088
rect 1104 19014 2582 19066
rect 2634 19014 2646 19066
rect 2698 19014 2710 19066
rect 2762 19014 2774 19066
rect 2826 19014 2838 19066
rect 2890 19014 5846 19066
rect 5898 19014 5910 19066
rect 5962 19014 5974 19066
rect 6026 19014 6038 19066
rect 6090 19014 6102 19066
rect 6154 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 9238 19066
rect 9290 19014 9302 19066
rect 9354 19014 9366 19066
rect 9418 19014 10856 19066
rect 1104 18992 10856 19014
rect 2130 18912 2136 18964
rect 2188 18952 2194 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 2188 18924 3801 18952
rect 2188 18912 2194 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 3789 18915 3847 18921
rect 1210 18776 1216 18828
rect 1268 18816 1274 18828
rect 1397 18819 1455 18825
rect 1397 18816 1409 18819
rect 1268 18788 1409 18816
rect 1268 18776 1274 18788
rect 1397 18785 1409 18788
rect 1443 18785 1455 18819
rect 1397 18779 1455 18785
rect 1673 18819 1731 18825
rect 1673 18785 1685 18819
rect 1719 18816 1731 18819
rect 2498 18816 2504 18828
rect 1719 18788 2504 18816
rect 1719 18785 1731 18788
rect 1673 18779 1731 18785
rect 2498 18776 2504 18788
rect 2556 18776 2562 18828
rect 2774 18776 2780 18828
rect 2832 18816 2838 18828
rect 2961 18819 3019 18825
rect 2961 18816 2973 18819
rect 2832 18788 2973 18816
rect 2832 18776 2838 18788
rect 2961 18785 2973 18788
rect 3007 18816 3019 18819
rect 3234 18816 3240 18828
rect 3007 18788 3240 18816
rect 3007 18785 3019 18788
rect 2961 18779 3019 18785
rect 3234 18776 3240 18788
rect 3292 18776 3298 18828
rect 2685 18751 2743 18757
rect 2685 18717 2697 18751
rect 2731 18717 2743 18751
rect 3970 18748 3976 18760
rect 3931 18720 3976 18748
rect 2685 18711 2743 18717
rect 2700 18680 2728 18711
rect 3970 18708 3976 18720
rect 4028 18708 4034 18760
rect 9858 18748 9864 18760
rect 9819 18720 9864 18748
rect 9858 18708 9864 18720
rect 9916 18708 9922 18760
rect 3234 18680 3240 18692
rect 2700 18652 3240 18680
rect 3234 18640 3240 18652
rect 3292 18680 3298 18692
rect 3878 18680 3884 18692
rect 3292 18652 3884 18680
rect 3292 18640 3298 18652
rect 3878 18640 3884 18652
rect 3936 18640 3942 18692
rect 10042 18612 10048 18624
rect 10003 18584 10048 18612
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 1104 18522 10856 18544
rect 1104 18470 4214 18522
rect 4266 18470 4278 18522
rect 4330 18470 4342 18522
rect 4394 18470 4406 18522
rect 4458 18470 4470 18522
rect 4522 18470 7478 18522
rect 7530 18470 7542 18522
rect 7594 18470 7606 18522
rect 7658 18470 7670 18522
rect 7722 18470 7734 18522
rect 7786 18470 10856 18522
rect 1104 18448 10856 18470
rect 2041 18411 2099 18417
rect 2041 18377 2053 18411
rect 2087 18408 2099 18411
rect 2958 18408 2964 18420
rect 2087 18380 2964 18408
rect 2087 18377 2099 18380
rect 2041 18371 2099 18377
rect 2958 18368 2964 18380
rect 3016 18368 3022 18420
rect 3513 18411 3571 18417
rect 3513 18377 3525 18411
rect 3559 18377 3571 18411
rect 3513 18371 3571 18377
rect 1946 18340 1952 18352
rect 1780 18312 1952 18340
rect 1780 18281 1808 18312
rect 1946 18300 1952 18312
rect 2004 18300 2010 18352
rect 2869 18343 2927 18349
rect 2869 18309 2881 18343
rect 2915 18340 2927 18343
rect 3142 18340 3148 18352
rect 2915 18312 3148 18340
rect 2915 18309 2927 18312
rect 2869 18303 2927 18309
rect 3142 18300 3148 18312
rect 3200 18300 3206 18352
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18241 1823 18275
rect 1765 18235 1823 18241
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18272 1915 18275
rect 2682 18272 2688 18284
rect 1903 18244 2688 18272
rect 1903 18241 1915 18244
rect 1857 18235 1915 18241
rect 2682 18232 2688 18244
rect 2740 18232 2746 18284
rect 3528 18272 3556 18371
rect 3694 18272 3700 18284
rect 2792 18244 3556 18272
rect 3655 18244 3700 18272
rect 2314 18164 2320 18216
rect 2372 18204 2378 18216
rect 2792 18204 2820 18244
rect 3694 18232 3700 18244
rect 3752 18232 3758 18284
rect 9858 18272 9864 18284
rect 9819 18244 9864 18272
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 3050 18204 3056 18216
rect 2372 18176 2820 18204
rect 2884 18176 3056 18204
rect 2372 18164 2378 18176
rect 2498 18136 2504 18148
rect 2459 18108 2504 18136
rect 2498 18096 2504 18108
rect 2556 18096 2562 18148
rect 2884 18077 2912 18176
rect 3050 18164 3056 18176
rect 3108 18164 3114 18216
rect 2869 18071 2927 18077
rect 2869 18037 2881 18071
rect 2915 18037 2927 18071
rect 2869 18031 2927 18037
rect 2958 18028 2964 18080
rect 3016 18068 3022 18080
rect 3053 18071 3111 18077
rect 3053 18068 3065 18071
rect 3016 18040 3065 18068
rect 3016 18028 3022 18040
rect 3053 18037 3065 18040
rect 3099 18037 3111 18071
rect 10042 18068 10048 18080
rect 10003 18040 10048 18068
rect 3053 18031 3111 18037
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 1104 17978 10856 18000
rect 1104 17926 2582 17978
rect 2634 17926 2646 17978
rect 2698 17926 2710 17978
rect 2762 17926 2774 17978
rect 2826 17926 2838 17978
rect 2890 17926 5846 17978
rect 5898 17926 5910 17978
rect 5962 17926 5974 17978
rect 6026 17926 6038 17978
rect 6090 17926 6102 17978
rect 6154 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 9238 17978
rect 9290 17926 9302 17978
rect 9354 17926 9366 17978
rect 9418 17926 10856 17978
rect 1104 17904 10856 17926
rect 1397 17867 1455 17873
rect 1397 17833 1409 17867
rect 1443 17864 1455 17867
rect 1946 17864 1952 17876
rect 1443 17836 1952 17864
rect 1443 17833 1455 17836
rect 1397 17827 1455 17833
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 3602 17824 3608 17876
rect 3660 17864 3666 17876
rect 3973 17867 4031 17873
rect 3973 17864 3985 17867
rect 3660 17836 3985 17864
rect 3660 17824 3666 17836
rect 3973 17833 3985 17836
rect 4019 17833 4031 17867
rect 3973 17827 4031 17833
rect 2409 17799 2467 17805
rect 2409 17765 2421 17799
rect 2455 17796 2467 17799
rect 3878 17796 3884 17808
rect 2455 17768 3884 17796
rect 2455 17765 2467 17768
rect 2409 17759 2467 17765
rect 3878 17756 3884 17768
rect 3936 17756 3942 17808
rect 4157 17799 4215 17805
rect 4157 17765 4169 17799
rect 4203 17765 4215 17799
rect 4157 17759 4215 17765
rect 3050 17728 3056 17740
rect 2884 17700 3056 17728
rect 1578 17660 1584 17672
rect 1539 17632 1584 17660
rect 1578 17620 1584 17632
rect 1636 17620 1642 17672
rect 2317 17663 2375 17669
rect 2317 17629 2329 17663
rect 2363 17660 2375 17663
rect 2498 17660 2504 17672
rect 2363 17632 2504 17660
rect 2363 17629 2375 17632
rect 2317 17623 2375 17629
rect 2498 17620 2504 17632
rect 2556 17620 2562 17672
rect 2884 17669 2912 17700
rect 3050 17688 3056 17700
rect 3108 17728 3114 17740
rect 4172 17728 4200 17759
rect 3108 17700 4200 17728
rect 3108 17688 3114 17700
rect 2869 17663 2927 17669
rect 2869 17629 2881 17663
rect 2915 17629 2927 17663
rect 3142 17660 3148 17672
rect 3103 17632 3148 17660
rect 2869 17623 2927 17629
rect 3142 17620 3148 17632
rect 3200 17620 3206 17672
rect 9030 17620 9036 17672
rect 9088 17660 9094 17672
rect 9861 17663 9919 17669
rect 9861 17660 9873 17663
rect 9088 17632 9873 17660
rect 9088 17620 9094 17632
rect 9861 17629 9873 17632
rect 9907 17629 9919 17663
rect 9861 17623 9919 17629
rect 1670 17552 1676 17604
rect 1728 17592 1734 17604
rect 1728 17564 2774 17592
rect 1728 17552 1734 17564
rect 2746 17524 2774 17564
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 3789 17595 3847 17601
rect 3789 17592 3801 17595
rect 3568 17564 3801 17592
rect 3568 17552 3574 17564
rect 3789 17561 3801 17564
rect 3835 17561 3847 17595
rect 3789 17555 3847 17561
rect 3970 17524 3976 17536
rect 4028 17533 4034 17536
rect 4028 17527 4047 17533
rect 2746 17496 3976 17524
rect 3970 17484 3976 17496
rect 4035 17493 4047 17527
rect 10042 17524 10048 17536
rect 10003 17496 10048 17524
rect 4028 17487 4047 17493
rect 4028 17484 4034 17487
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 1104 17434 10856 17456
rect 1104 17382 4214 17434
rect 4266 17382 4278 17434
rect 4330 17382 4342 17434
rect 4394 17382 4406 17434
rect 4458 17382 4470 17434
rect 4522 17382 7478 17434
rect 7530 17382 7542 17434
rect 7594 17382 7606 17434
rect 7658 17382 7670 17434
rect 7722 17382 7734 17434
rect 7786 17382 10856 17434
rect 1104 17360 10856 17382
rect 1118 17280 1124 17332
rect 1176 17320 1182 17332
rect 1949 17323 2007 17329
rect 1949 17320 1961 17323
rect 1176 17292 1961 17320
rect 1176 17280 1182 17292
rect 1949 17289 1961 17292
rect 1995 17289 2007 17323
rect 1949 17283 2007 17289
rect 4706 17280 4712 17332
rect 4764 17320 4770 17332
rect 4982 17320 4988 17332
rect 4764 17292 4988 17320
rect 4764 17280 4770 17292
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 9953 17323 10011 17329
rect 9953 17320 9965 17323
rect 9916 17292 9965 17320
rect 9916 17280 9922 17292
rect 9953 17289 9965 17292
rect 9999 17289 10011 17323
rect 9953 17283 10011 17289
rect 1857 17255 1915 17261
rect 1857 17221 1869 17255
rect 1903 17252 1915 17255
rect 3878 17252 3884 17264
rect 1903 17224 3884 17252
rect 1903 17221 1915 17224
rect 1857 17215 1915 17221
rect 3878 17212 3884 17224
rect 3936 17212 3942 17264
rect 2958 17184 2964 17196
rect 2919 17156 2964 17184
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 3970 17144 3976 17196
rect 4028 17184 4034 17196
rect 10137 17187 10195 17193
rect 10137 17184 10149 17187
rect 4028 17156 10149 17184
rect 4028 17144 4034 17156
rect 10137 17153 10149 17156
rect 10183 17153 10195 17187
rect 10137 17147 10195 17153
rect 3234 17116 3240 17128
rect 3195 17088 3240 17116
rect 3234 17076 3240 17088
rect 3292 17076 3298 17128
rect 4614 16940 4620 16992
rect 4672 16980 4678 16992
rect 4798 16980 4804 16992
rect 4672 16952 4804 16980
rect 4672 16940 4678 16952
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 1104 16890 10856 16912
rect 1104 16838 2582 16890
rect 2634 16838 2646 16890
rect 2698 16838 2710 16890
rect 2762 16838 2774 16890
rect 2826 16838 2838 16890
rect 2890 16838 5846 16890
rect 5898 16838 5910 16890
rect 5962 16838 5974 16890
rect 6026 16838 6038 16890
rect 6090 16838 6102 16890
rect 6154 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 9238 16890
rect 9290 16838 9302 16890
rect 9354 16838 9366 16890
rect 9418 16838 10856 16890
rect 1104 16816 10856 16838
rect 1210 16532 1216 16584
rect 1268 16572 1274 16584
rect 1581 16575 1639 16581
rect 1581 16572 1593 16575
rect 1268 16544 1593 16572
rect 1268 16532 1274 16544
rect 1581 16541 1593 16544
rect 1627 16541 1639 16575
rect 2406 16572 2412 16584
rect 2367 16544 2412 16572
rect 1581 16535 1639 16541
rect 2406 16532 2412 16544
rect 2464 16532 2470 16584
rect 3050 16572 3056 16584
rect 3011 16544 3056 16572
rect 3050 16532 3056 16544
rect 3108 16532 3114 16584
rect 3970 16572 3976 16584
rect 3931 16544 3976 16572
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 9214 16532 9220 16584
rect 9272 16572 9278 16584
rect 9861 16575 9919 16581
rect 9861 16572 9873 16575
rect 9272 16544 9873 16572
rect 9272 16532 9278 16544
rect 9861 16541 9873 16544
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 3326 16504 3332 16516
rect 2884 16476 3332 16504
rect 1397 16439 1455 16445
rect 1397 16405 1409 16439
rect 1443 16436 1455 16439
rect 1578 16436 1584 16448
rect 1443 16408 1584 16436
rect 1443 16405 1455 16408
rect 1397 16399 1455 16405
rect 1578 16396 1584 16408
rect 1636 16396 1642 16448
rect 2222 16436 2228 16448
rect 2183 16408 2228 16436
rect 2222 16396 2228 16408
rect 2280 16396 2286 16448
rect 2884 16445 2912 16476
rect 3326 16464 3332 16476
rect 3384 16464 3390 16516
rect 2869 16439 2927 16445
rect 2869 16405 2881 16439
rect 2915 16405 2927 16439
rect 2869 16399 2927 16405
rect 3234 16396 3240 16448
rect 3292 16436 3298 16448
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 3292 16408 3801 16436
rect 3292 16396 3298 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 10042 16436 10048 16448
rect 10003 16408 10048 16436
rect 3789 16399 3847 16405
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 1104 16346 10856 16368
rect 1104 16294 4214 16346
rect 4266 16294 4278 16346
rect 4330 16294 4342 16346
rect 4394 16294 4406 16346
rect 4458 16294 4470 16346
rect 4522 16294 7478 16346
rect 7530 16294 7542 16346
rect 7594 16294 7606 16346
rect 7658 16294 7670 16346
rect 7722 16294 7734 16346
rect 7786 16294 10856 16346
rect 1104 16272 10856 16294
rect 9214 16232 9220 16244
rect 9175 16204 9220 16232
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 1394 16056 1400 16108
rect 1452 16096 1458 16108
rect 1581 16099 1639 16105
rect 1581 16096 1593 16099
rect 1452 16068 1593 16096
rect 1452 16056 1458 16068
rect 1581 16065 1593 16068
rect 1627 16065 1639 16099
rect 2222 16096 2228 16108
rect 2183 16068 2228 16096
rect 1581 16059 1639 16065
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 2866 16096 2872 16108
rect 2827 16068 2872 16096
rect 2866 16056 2872 16068
rect 2924 16056 2930 16108
rect 3694 16056 3700 16108
rect 3752 16096 3758 16108
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 3752 16068 9413 16096
rect 3752 16056 3758 16068
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 9950 16096 9956 16108
rect 9907 16068 9956 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 9950 16056 9956 16068
rect 10008 16056 10014 16108
rect 1397 15895 1455 15901
rect 1397 15861 1409 15895
rect 1443 15892 1455 15895
rect 1486 15892 1492 15904
rect 1443 15864 1492 15892
rect 1443 15861 1455 15864
rect 1397 15855 1455 15861
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 2038 15892 2044 15904
rect 1999 15864 2044 15892
rect 2038 15852 2044 15864
rect 2096 15852 2102 15904
rect 2130 15852 2136 15904
rect 2188 15892 2194 15904
rect 2685 15895 2743 15901
rect 2685 15892 2697 15895
rect 2188 15864 2697 15892
rect 2188 15852 2194 15864
rect 2685 15861 2697 15864
rect 2731 15861 2743 15895
rect 10042 15892 10048 15904
rect 10003 15864 10048 15892
rect 2685 15855 2743 15861
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 1104 15802 10856 15824
rect 1104 15750 2582 15802
rect 2634 15750 2646 15802
rect 2698 15750 2710 15802
rect 2762 15750 2774 15802
rect 2826 15750 2838 15802
rect 2890 15750 5846 15802
rect 5898 15750 5910 15802
rect 5962 15750 5974 15802
rect 6026 15750 6038 15802
rect 6090 15750 6102 15802
rect 6154 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 9238 15802
rect 9290 15750 9302 15802
rect 9354 15750 9366 15802
rect 9418 15750 10856 15802
rect 1104 15728 10856 15750
rect 1949 15691 2007 15697
rect 1949 15657 1961 15691
rect 1995 15688 2007 15691
rect 2130 15688 2136 15700
rect 1995 15660 2136 15688
rect 1995 15657 2007 15660
rect 1949 15651 2007 15657
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 9950 15688 9956 15700
rect 9911 15660 9956 15688
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 2869 15623 2927 15629
rect 2869 15589 2881 15623
rect 2915 15620 2927 15623
rect 4982 15620 4988 15632
rect 2915 15592 4988 15620
rect 2915 15589 2927 15592
rect 2869 15583 2927 15589
rect 4982 15580 4988 15592
rect 5040 15580 5046 15632
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15552 1547 15555
rect 2038 15552 2044 15564
rect 1535 15524 2044 15552
rect 1535 15521 1547 15524
rect 1489 15515 1547 15521
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 1578 15444 1584 15496
rect 1636 15484 1642 15496
rect 1949 15487 2007 15493
rect 1636 15456 1681 15484
rect 1636 15444 1642 15456
rect 1949 15453 1961 15487
rect 1995 15484 2007 15487
rect 3234 15484 3240 15496
rect 1995 15456 3240 15484
rect 1995 15453 2007 15456
rect 1949 15447 2007 15453
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 10137 15487 10195 15493
rect 10137 15453 10149 15487
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 2685 15419 2743 15425
rect 2685 15385 2697 15419
rect 2731 15416 2743 15419
rect 3510 15416 3516 15428
rect 2731 15388 3516 15416
rect 2731 15385 2743 15388
rect 2685 15379 2743 15385
rect 3510 15376 3516 15388
rect 3568 15376 3574 15428
rect 2130 15348 2136 15360
rect 2091 15320 2136 15348
rect 2130 15308 2136 15320
rect 2188 15308 2194 15360
rect 2406 15308 2412 15360
rect 2464 15348 2470 15360
rect 10152 15348 10180 15447
rect 2464 15320 10180 15348
rect 2464 15308 2470 15320
rect 1104 15258 10856 15280
rect 1104 15206 4214 15258
rect 4266 15206 4278 15258
rect 4330 15206 4342 15258
rect 4394 15206 4406 15258
rect 4458 15206 4470 15258
rect 4522 15206 7478 15258
rect 7530 15206 7542 15258
rect 7594 15206 7606 15258
rect 7658 15206 7670 15258
rect 7722 15206 7734 15258
rect 7786 15206 10856 15258
rect 1104 15184 10856 15206
rect 2041 15147 2099 15153
rect 2041 15113 2053 15147
rect 2087 15144 2099 15147
rect 8570 15144 8576 15156
rect 2087 15116 8576 15144
rect 2087 15113 2099 15116
rect 2041 15107 2099 15113
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 1949 15079 2007 15085
rect 1949 15045 1961 15079
rect 1995 15076 2007 15079
rect 3050 15076 3056 15088
rect 1995 15048 3056 15076
rect 1995 15045 2007 15048
rect 1949 15039 2007 15045
rect 3050 15036 3056 15048
rect 3108 15036 3114 15088
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 15008 2835 15011
rect 2958 15008 2964 15020
rect 2823 14980 2964 15008
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 2958 14968 2964 14980
rect 3016 14968 3022 15020
rect 9490 14968 9496 15020
rect 9548 15008 9554 15020
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 9548 14980 9873 15008
rect 9548 14968 9554 14980
rect 9861 14977 9873 14980
rect 9907 14977 9919 15011
rect 9861 14971 9919 14977
rect 10042 14872 10048 14884
rect 10003 14844 10048 14872
rect 10042 14832 10048 14844
rect 10100 14832 10106 14884
rect 1670 14764 1676 14816
rect 1728 14804 1734 14816
rect 2593 14807 2651 14813
rect 2593 14804 2605 14807
rect 1728 14776 2605 14804
rect 1728 14764 1734 14776
rect 2593 14773 2605 14776
rect 2639 14773 2651 14807
rect 2593 14767 2651 14773
rect 1104 14714 10856 14736
rect 1104 14662 2582 14714
rect 2634 14662 2646 14714
rect 2698 14662 2710 14714
rect 2762 14662 2774 14714
rect 2826 14662 2838 14714
rect 2890 14662 5846 14714
rect 5898 14662 5910 14714
rect 5962 14662 5974 14714
rect 6026 14662 6038 14714
rect 6090 14662 6102 14714
rect 6154 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 9238 14714
rect 9290 14662 9302 14714
rect 9354 14662 9366 14714
rect 9418 14662 10856 14714
rect 1104 14640 10856 14662
rect 1673 14603 1731 14609
rect 1673 14569 1685 14603
rect 1719 14600 1731 14603
rect 1762 14600 1768 14612
rect 1719 14572 1768 14600
rect 1719 14569 1731 14572
rect 1673 14563 1731 14569
rect 1762 14560 1768 14572
rect 1820 14560 1826 14612
rect 1857 14603 1915 14609
rect 1857 14569 1869 14603
rect 1903 14600 1915 14603
rect 2317 14603 2375 14609
rect 2317 14600 2329 14603
rect 1903 14572 2329 14600
rect 1903 14569 1915 14572
rect 1857 14563 1915 14569
rect 2317 14569 2329 14572
rect 2363 14569 2375 14603
rect 2317 14563 2375 14569
rect 2498 14560 2504 14612
rect 2556 14600 2562 14612
rect 2685 14603 2743 14609
rect 2685 14600 2697 14603
rect 2556 14572 2697 14600
rect 2556 14560 2562 14572
rect 2685 14569 2697 14572
rect 2731 14569 2743 14603
rect 2685 14563 2743 14569
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 2130 14424 2136 14476
rect 2188 14464 2194 14476
rect 2409 14467 2467 14473
rect 2409 14464 2421 14467
rect 2188 14436 2421 14464
rect 2188 14424 2194 14436
rect 2409 14433 2421 14436
rect 2455 14433 2467 14467
rect 2409 14427 2467 14433
rect 1670 14396 1676 14408
rect 1631 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 2314 14396 2320 14408
rect 2275 14368 2320 14396
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 3970 14396 3976 14408
rect 3931 14368 3976 14396
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 9858 14396 9864 14408
rect 9819 14368 9864 14396
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 1397 14331 1455 14337
rect 1397 14297 1409 14331
rect 1443 14328 1455 14331
rect 1443 14300 2774 14328
rect 1443 14297 1455 14300
rect 1397 14291 1455 14297
rect 1578 14220 1584 14272
rect 1636 14260 1642 14272
rect 1946 14260 1952 14272
rect 1636 14232 1952 14260
rect 1636 14220 1642 14232
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 2746 14260 2774 14300
rect 3789 14263 3847 14269
rect 3789 14260 3801 14263
rect 2746 14232 3801 14260
rect 3789 14229 3801 14232
rect 3835 14229 3847 14263
rect 10042 14260 10048 14272
rect 10003 14232 10048 14260
rect 3789 14223 3847 14229
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 1104 14170 10856 14192
rect 1104 14118 4214 14170
rect 4266 14118 4278 14170
rect 4330 14118 4342 14170
rect 4394 14118 4406 14170
rect 4458 14118 4470 14170
rect 4522 14118 7478 14170
rect 7530 14118 7542 14170
rect 7594 14118 7606 14170
rect 7658 14118 7670 14170
rect 7722 14118 7734 14170
rect 7786 14118 10856 14170
rect 1104 14096 10856 14118
rect 2593 14059 2651 14065
rect 2593 14025 2605 14059
rect 2639 14056 2651 14059
rect 9217 14059 9275 14065
rect 2639 14028 6316 14056
rect 2639 14025 2651 14028
rect 2593 14019 2651 14025
rect 2222 13948 2228 14000
rect 2280 13988 2286 14000
rect 3602 13988 3608 14000
rect 2280 13960 3608 13988
rect 2280 13948 2286 13960
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 2792 13929 2820 13960
rect 3602 13948 3608 13960
rect 3660 13948 3666 14000
rect 6288 13988 6316 14028
rect 9217 14025 9229 14059
rect 9263 14056 9275 14059
rect 9490 14056 9496 14068
rect 9263 14028 9496 14056
rect 9263 14025 9275 14028
rect 9217 14019 9275 14025
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 9582 14016 9588 14068
rect 9640 14056 9646 14068
rect 10045 14059 10103 14065
rect 10045 14056 10057 14059
rect 9640 14028 10057 14056
rect 9640 14016 9646 14028
rect 10045 14025 10057 14028
rect 10091 14025 10103 14059
rect 10045 14019 10103 14025
rect 6288 13960 9904 13988
rect 1581 13923 1639 13929
rect 1581 13920 1593 13923
rect 1544 13892 1593 13920
rect 1544 13880 1550 13892
rect 1581 13889 1593 13892
rect 1627 13889 1639 13923
rect 1581 13883 1639 13889
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13920 2835 13923
rect 3418 13920 3424 13932
rect 2823 13892 2857 13920
rect 3379 13892 3424 13920
rect 2823 13889 2835 13892
rect 2777 13883 2835 13889
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 9876 13929 9904 13960
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13889 9459 13923
rect 9401 13883 9459 13889
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 1762 13812 1768 13864
rect 1820 13852 1826 13864
rect 9416 13852 9444 13883
rect 1820 13824 3280 13852
rect 1820 13812 1826 13824
rect 3252 13793 3280 13824
rect 3344 13824 9444 13852
rect 3237 13787 3295 13793
rect 3237 13753 3249 13787
rect 3283 13753 3295 13787
rect 3237 13747 3295 13753
rect 1394 13716 1400 13728
rect 1355 13688 1400 13716
rect 1394 13676 1400 13688
rect 1452 13676 1458 13728
rect 2406 13676 2412 13728
rect 2464 13716 2470 13728
rect 3344 13716 3372 13824
rect 2464 13688 3372 13716
rect 2464 13676 2470 13688
rect 1104 13626 10856 13648
rect 1104 13574 2582 13626
rect 2634 13574 2646 13626
rect 2698 13574 2710 13626
rect 2762 13574 2774 13626
rect 2826 13574 2838 13626
rect 2890 13574 5846 13626
rect 5898 13574 5910 13626
rect 5962 13574 5974 13626
rect 6026 13574 6038 13626
rect 6090 13574 6102 13626
rect 6154 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 9238 13626
rect 9290 13574 9302 13626
rect 9354 13574 9366 13626
rect 9418 13574 10856 13626
rect 1104 13552 10856 13574
rect 3050 13512 3056 13524
rect 2608 13484 2774 13512
rect 3011 13484 3056 13512
rect 2038 13404 2044 13456
rect 2096 13444 2102 13456
rect 2498 13444 2504 13456
rect 2096 13416 2504 13444
rect 2096 13404 2102 13416
rect 2498 13404 2504 13416
rect 2556 13404 2562 13456
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 2222 13268 2228 13320
rect 2280 13308 2286 13320
rect 2608 13308 2636 13484
rect 2746 13444 2774 13484
rect 3050 13472 3056 13484
rect 3108 13472 3114 13524
rect 9030 13472 9036 13524
rect 9088 13512 9094 13524
rect 9309 13515 9367 13521
rect 9309 13512 9321 13515
rect 9088 13484 9321 13512
rect 9088 13472 9094 13484
rect 9309 13481 9321 13484
rect 9355 13481 9367 13515
rect 9309 13475 9367 13481
rect 9858 13472 9864 13524
rect 9916 13512 9922 13524
rect 9953 13515 10011 13521
rect 9953 13512 9965 13515
rect 9916 13484 9965 13512
rect 9916 13472 9922 13484
rect 9953 13481 9965 13484
rect 9999 13481 10011 13515
rect 9953 13475 10011 13481
rect 2746 13416 10180 13444
rect 2777 13311 2835 13317
rect 2777 13308 2789 13311
rect 2280 13280 2789 13308
rect 2280 13268 2286 13280
rect 2777 13277 2789 13280
rect 2823 13277 2835 13311
rect 2777 13271 2835 13277
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 3970 13308 3976 13320
rect 2915 13280 3832 13308
rect 3931 13280 3976 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 3804 13240 3832 13280
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 9490 13308 9496 13320
rect 9451 13280 9496 13308
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 10152 13317 10180 13416
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 3878 13240 3884 13252
rect 3804 13212 3884 13240
rect 3878 13200 3884 13212
rect 3936 13200 3942 13252
rect 1397 13175 1455 13181
rect 1397 13141 1409 13175
rect 1443 13172 1455 13175
rect 1670 13172 1676 13184
rect 1443 13144 1676 13172
rect 1443 13141 1455 13144
rect 1397 13135 1455 13141
rect 1670 13132 1676 13144
rect 1728 13132 1734 13184
rect 2406 13132 2412 13184
rect 2464 13172 2470 13184
rect 2685 13175 2743 13181
rect 2685 13172 2697 13175
rect 2464 13144 2697 13172
rect 2464 13132 2470 13144
rect 2685 13141 2697 13144
rect 2731 13141 2743 13175
rect 2685 13135 2743 13141
rect 3234 13132 3240 13184
rect 3292 13172 3298 13184
rect 3789 13175 3847 13181
rect 3789 13172 3801 13175
rect 3292 13144 3801 13172
rect 3292 13132 3298 13144
rect 3789 13141 3801 13144
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 1104 13082 10856 13104
rect 1104 13030 4214 13082
rect 4266 13030 4278 13082
rect 4330 13030 4342 13082
rect 4394 13030 4406 13082
rect 4458 13030 4470 13082
rect 4522 13030 7478 13082
rect 7530 13030 7542 13082
rect 7594 13030 7606 13082
rect 7658 13030 7670 13082
rect 7722 13030 7734 13082
rect 7786 13030 10856 13082
rect 1104 13008 10856 13030
rect 1857 12971 1915 12977
rect 1857 12937 1869 12971
rect 1903 12968 1915 12971
rect 2314 12968 2320 12980
rect 1903 12940 2320 12968
rect 1903 12937 1915 12940
rect 1857 12931 1915 12937
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 2895 12971 2953 12977
rect 2895 12937 2907 12971
rect 2941 12968 2953 12971
rect 3050 12968 3056 12980
rect 2941 12940 3056 12968
rect 2941 12937 2953 12940
rect 2895 12931 2953 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 3513 12971 3571 12977
rect 3513 12937 3525 12971
rect 3559 12937 3571 12971
rect 3513 12931 3571 12937
rect 1394 12900 1400 12912
rect 1355 12872 1400 12900
rect 1394 12860 1400 12872
rect 1452 12860 1458 12912
rect 1762 12860 1768 12912
rect 1820 12900 1826 12912
rect 2685 12903 2743 12909
rect 2685 12900 2697 12903
rect 1820 12872 2697 12900
rect 1820 12860 1826 12872
rect 2685 12869 2697 12872
rect 2731 12900 2743 12903
rect 3528 12900 3556 12931
rect 2731 12872 3464 12900
rect 3528 12872 9904 12900
rect 2731 12869 2743 12872
rect 2685 12863 2743 12869
rect 1670 12832 1676 12844
rect 1631 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 3234 12832 3240 12844
rect 2746 12804 3240 12832
rect 1581 12767 1639 12773
rect 1581 12733 1593 12767
rect 1627 12764 1639 12767
rect 2746 12764 2774 12804
rect 3234 12792 3240 12804
rect 3292 12792 3298 12844
rect 1627 12736 2774 12764
rect 3436 12764 3464 12872
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 3786 12832 3792 12844
rect 3743 12804 3792 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 9876 12841 9904 12872
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 9490 12764 9496 12776
rect 3436 12736 9496 12764
rect 1627 12733 1639 12736
rect 1581 12727 1639 12733
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 2958 12696 2964 12708
rect 1688 12668 2964 12696
rect 1688 12637 1716 12668
rect 2958 12656 2964 12668
rect 3016 12656 3022 12708
rect 3053 12699 3111 12705
rect 3053 12665 3065 12699
rect 3099 12696 3111 12699
rect 3142 12696 3148 12708
rect 3099 12668 3148 12696
rect 3099 12665 3111 12668
rect 3053 12659 3111 12665
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 3694 12656 3700 12708
rect 3752 12696 3758 12708
rect 3970 12696 3976 12708
rect 3752 12668 3976 12696
rect 3752 12656 3758 12668
rect 3970 12656 3976 12668
rect 4028 12656 4034 12708
rect 1673 12631 1731 12637
rect 1673 12597 1685 12631
rect 1719 12597 1731 12631
rect 1673 12591 1731 12597
rect 2869 12631 2927 12637
rect 2869 12597 2881 12631
rect 2915 12628 2927 12631
rect 3712 12628 3740 12656
rect 10042 12628 10048 12640
rect 2915 12600 3740 12628
rect 10003 12600 10048 12628
rect 2915 12597 2927 12600
rect 2869 12591 2927 12597
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 1104 12538 10856 12560
rect 1104 12486 2582 12538
rect 2634 12486 2646 12538
rect 2698 12486 2710 12538
rect 2762 12486 2774 12538
rect 2826 12486 2838 12538
rect 2890 12486 5846 12538
rect 5898 12486 5910 12538
rect 5962 12486 5974 12538
rect 6026 12486 6038 12538
rect 6090 12486 6102 12538
rect 6154 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 9238 12538
rect 9290 12486 9302 12538
rect 9354 12486 9366 12538
rect 9418 12486 10856 12538
rect 1104 12464 10856 12486
rect 4706 12384 4712 12436
rect 4764 12384 4770 12436
rect 1673 12291 1731 12297
rect 1673 12257 1685 12291
rect 1719 12288 1731 12291
rect 3878 12288 3884 12300
rect 1719 12260 3884 12288
rect 1719 12257 1731 12260
rect 1673 12251 1731 12257
rect 3878 12248 3884 12260
rect 3936 12248 3942 12300
rect 4724 12232 4752 12384
rect 1210 12180 1216 12232
rect 1268 12220 1274 12232
rect 1397 12223 1455 12229
rect 1397 12220 1409 12223
rect 1268 12192 1409 12220
rect 1268 12180 1274 12192
rect 1397 12189 1409 12192
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 2130 12180 2136 12232
rect 2188 12220 2194 12232
rect 2869 12223 2927 12229
rect 2869 12220 2881 12223
rect 2188 12192 2881 12220
rect 2188 12180 2194 12192
rect 2869 12189 2881 12192
rect 2915 12220 2927 12223
rect 4614 12220 4620 12232
rect 2915 12192 4620 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 4706 12180 4712 12232
rect 4764 12180 4770 12232
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 2685 12087 2743 12093
rect 2685 12053 2697 12087
rect 2731 12084 2743 12087
rect 9876 12084 9904 12183
rect 10042 12084 10048 12096
rect 2731 12056 9904 12084
rect 10003 12056 10048 12084
rect 2731 12053 2743 12056
rect 2685 12047 2743 12053
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 1104 11994 10856 12016
rect 1104 11942 4214 11994
rect 4266 11942 4278 11994
rect 4330 11942 4342 11994
rect 4394 11942 4406 11994
rect 4458 11942 4470 11994
rect 4522 11942 7478 11994
rect 7530 11942 7542 11994
rect 7594 11942 7606 11994
rect 7658 11942 7670 11994
rect 7722 11942 7734 11994
rect 7786 11942 10856 11994
rect 1104 11920 10856 11942
rect 3050 11880 3056 11892
rect 3011 11852 3056 11880
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 9953 11883 10011 11889
rect 9953 11849 9965 11883
rect 9999 11880 10011 11883
rect 10134 11880 10140 11892
rect 9999 11852 10140 11880
rect 9999 11849 10011 11852
rect 9953 11843 10011 11849
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 3234 11812 3240 11824
rect 1688 11784 3240 11812
rect 1688 11753 1716 11784
rect 3234 11772 3240 11784
rect 3292 11772 3298 11824
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 3050 11744 3056 11756
rect 2915 11716 3056 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 3694 11744 3700 11756
rect 3655 11716 3700 11744
rect 3694 11704 3700 11716
rect 3752 11704 3758 11756
rect 3878 11704 3884 11756
rect 3936 11744 3942 11756
rect 10137 11747 10195 11753
rect 10137 11744 10149 11747
rect 3936 11716 10149 11744
rect 3936 11704 3942 11716
rect 10137 11713 10149 11716
rect 10183 11713 10195 11747
rect 10137 11707 10195 11713
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 2731 11648 3740 11676
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 2958 11568 2964 11620
rect 3016 11608 3022 11620
rect 3513 11611 3571 11617
rect 3513 11608 3525 11611
rect 3016 11580 3525 11608
rect 3016 11568 3022 11580
rect 3513 11577 3525 11580
rect 3559 11577 3571 11611
rect 3513 11571 3571 11577
rect 3712 11552 3740 11648
rect 3694 11500 3700 11552
rect 3752 11500 3758 11552
rect 1104 11450 10856 11472
rect 1104 11398 2582 11450
rect 2634 11398 2646 11450
rect 2698 11398 2710 11450
rect 2762 11398 2774 11450
rect 2826 11398 2838 11450
rect 2890 11398 5846 11450
rect 5898 11398 5910 11450
rect 5962 11398 5974 11450
rect 6026 11398 6038 11450
rect 6090 11398 6102 11450
rect 6154 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 9238 11450
rect 9290 11398 9302 11450
rect 9354 11398 9366 11450
rect 9418 11398 10856 11450
rect 1104 11376 10856 11398
rect 3053 11339 3111 11345
rect 3053 11305 3065 11339
rect 3099 11336 3111 11339
rect 3326 11336 3332 11348
rect 3099 11308 3332 11336
rect 3099 11305 3111 11308
rect 3053 11299 3111 11305
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 3418 11268 3424 11280
rect 1688 11240 3424 11268
rect 1688 11209 1716 11240
rect 3418 11228 3424 11240
rect 3476 11228 3482 11280
rect 10042 11268 10048 11280
rect 10003 11240 10048 11268
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11169 1731 11203
rect 1673 11163 1731 11169
rect 2130 11160 2136 11212
rect 2188 11200 2194 11212
rect 3050 11200 3056 11212
rect 2188 11172 3056 11200
rect 2188 11160 2194 11172
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 1486 11132 1492 11144
rect 1443 11104 1492 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 2884 11141 2912 11172
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11101 2835 11135
rect 2777 11095 2835 11101
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 9858 11132 9864 11144
rect 9819 11104 9864 11132
rect 2869 11095 2927 11101
rect 2792 11064 2820 11095
rect 9858 11092 9864 11104
rect 9916 11092 9922 11144
rect 3326 11064 3332 11076
rect 2792 11036 3332 11064
rect 3326 11024 3332 11036
rect 3384 11024 3390 11076
rect 1104 10906 10856 10928
rect 1104 10854 4214 10906
rect 4266 10854 4278 10906
rect 4330 10854 4342 10906
rect 4394 10854 4406 10906
rect 4458 10854 4470 10906
rect 4522 10854 7478 10906
rect 7530 10854 7542 10906
rect 7594 10854 7606 10906
rect 7658 10854 7670 10906
rect 7722 10854 7734 10906
rect 7786 10854 10856 10906
rect 1104 10832 10856 10854
rect 3421 10795 3479 10801
rect 3421 10761 3433 10795
rect 3467 10792 3479 10795
rect 9858 10792 9864 10804
rect 3467 10764 9864 10792
rect 3467 10761 3479 10764
rect 3421 10755 3479 10761
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 1946 10656 1952 10668
rect 1719 10628 1952 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 3234 10656 3240 10668
rect 2731 10628 3240 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 3234 10616 3240 10628
rect 3292 10616 3298 10668
rect 3510 10616 3516 10668
rect 3568 10656 3574 10668
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 3568 10628 3617 10656
rect 3568 10616 3574 10628
rect 3605 10625 3617 10628
rect 3651 10656 3663 10659
rect 4062 10656 4068 10668
rect 3651 10628 4068 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 9858 10656 9864 10668
rect 9819 10628 9864 10656
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 2869 10523 2927 10529
rect 2869 10489 2881 10523
rect 2915 10520 2927 10523
rect 4890 10520 4896 10532
rect 2915 10492 4896 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 4890 10480 4896 10492
rect 4948 10480 4954 10532
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 1104 10362 10856 10384
rect 1104 10310 2582 10362
rect 2634 10310 2646 10362
rect 2698 10310 2710 10362
rect 2762 10310 2774 10362
rect 2826 10310 2838 10362
rect 2890 10310 5846 10362
rect 5898 10310 5910 10362
rect 5962 10310 5974 10362
rect 6026 10310 6038 10362
rect 6090 10310 6102 10362
rect 6154 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 9238 10362
rect 9290 10310 9302 10362
rect 9354 10310 9366 10362
rect 9418 10310 10856 10362
rect 1104 10288 10856 10310
rect 3970 10248 3976 10260
rect 3931 10220 3976 10248
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 2869 10183 2927 10189
rect 2869 10149 2881 10183
rect 2915 10180 2927 10183
rect 4706 10180 4712 10192
rect 2915 10152 4712 10180
rect 2915 10149 2927 10152
rect 2869 10143 2927 10149
rect 4706 10140 4712 10152
rect 4764 10140 4770 10192
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 1762 10112 1768 10124
rect 1719 10084 1768 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 1762 10072 1768 10084
rect 1820 10072 1826 10124
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 1486 10044 1492 10056
rect 1443 10016 1492 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10044 2743 10047
rect 3142 10044 3148 10056
rect 2731 10016 3148 10044
rect 2731 10013 2743 10016
rect 2685 10007 2743 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10044 3847 10047
rect 3970 10044 3976 10056
rect 3835 10016 3976 10044
rect 3835 10013 3847 10016
rect 3789 10007 3847 10013
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 1104 9818 10856 9840
rect 1104 9766 4214 9818
rect 4266 9766 4278 9818
rect 4330 9766 4342 9818
rect 4394 9766 4406 9818
rect 4458 9766 4470 9818
rect 4522 9766 7478 9818
rect 7530 9766 7542 9818
rect 7594 9766 7606 9818
rect 7658 9766 7670 9818
rect 7722 9766 7734 9818
rect 7786 9766 10856 9818
rect 1104 9744 10856 9766
rect 3878 9636 3884 9648
rect 1688 9608 3884 9636
rect 1688 9577 1716 9608
rect 3878 9596 3884 9608
rect 3936 9596 3942 9648
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 2700 9364 2728 9531
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 3476 9540 3617 9568
rect 3476 9528 3482 9540
rect 3605 9537 3617 9540
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9568 4307 9571
rect 4706 9568 4712 9580
rect 4295 9540 4712 9568
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 9876 9500 9904 9531
rect 3436 9472 9904 9500
rect 3050 9432 3056 9444
rect 2792 9404 3056 9432
rect 2792 9364 2820 9404
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 3436 9441 3464 9472
rect 3421 9435 3479 9441
rect 3421 9401 3433 9435
rect 3467 9401 3479 9435
rect 3421 9395 3479 9401
rect 4065 9435 4123 9441
rect 4065 9401 4077 9435
rect 4111 9432 4123 9435
rect 9858 9432 9864 9444
rect 4111 9404 9864 9432
rect 4111 9401 4123 9404
rect 4065 9395 4123 9401
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 10042 9432 10048 9444
rect 10003 9404 10048 9432
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 2700 9336 2820 9364
rect 2869 9367 2927 9373
rect 2869 9333 2881 9367
rect 2915 9364 2927 9367
rect 8294 9364 8300 9376
rect 2915 9336 8300 9364
rect 2915 9333 2927 9336
rect 2869 9327 2927 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 1104 9274 10856 9296
rect 1104 9222 2582 9274
rect 2634 9222 2646 9274
rect 2698 9222 2710 9274
rect 2762 9222 2774 9274
rect 2826 9222 2838 9274
rect 2890 9222 5846 9274
rect 5898 9222 5910 9274
rect 5962 9222 5974 9274
rect 6026 9222 6038 9274
rect 6090 9222 6102 9274
rect 6154 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 9238 9274
rect 9290 9222 9302 9274
rect 9354 9222 9366 9274
rect 9418 9222 10856 9274
rect 1104 9200 10856 9222
rect 3050 9120 3056 9172
rect 3108 9160 3114 9172
rect 3878 9160 3884 9172
rect 3108 9132 3884 9160
rect 3108 9120 3114 9132
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 9024 1731 9027
rect 2038 9024 2044 9036
rect 1719 8996 2044 9024
rect 1719 8993 1731 8996
rect 1673 8987 1731 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 3234 8956 3240 8968
rect 3195 8928 3240 8956
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3970 8956 3976 8968
rect 3931 8928 3976 8956
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 9876 8888 9904 8919
rect 3804 8860 9904 8888
rect 3050 8820 3056 8832
rect 3011 8792 3056 8820
rect 3050 8780 3056 8792
rect 3108 8780 3114 8832
rect 3804 8829 3832 8860
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8789 3847 8823
rect 10042 8820 10048 8832
rect 10003 8792 10048 8820
rect 3789 8783 3847 8789
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 1104 8730 10856 8752
rect 1104 8678 4214 8730
rect 4266 8678 4278 8730
rect 4330 8678 4342 8730
rect 4394 8678 4406 8730
rect 4458 8678 4470 8730
rect 4522 8678 7478 8730
rect 7530 8678 7542 8730
rect 7594 8678 7606 8730
rect 7658 8678 7670 8730
rect 7722 8678 7734 8730
rect 7786 8678 10856 8730
rect 1104 8656 10856 8678
rect 2869 8619 2927 8625
rect 2869 8585 2881 8619
rect 2915 8616 2927 8619
rect 3602 8616 3608 8628
rect 2915 8588 3608 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2406 8480 2412 8492
rect 1719 8452 2412 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8480 2743 8483
rect 2958 8480 2964 8492
rect 2731 8452 2964 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 3050 8440 3056 8492
rect 3108 8480 3114 8492
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 3108 8452 9873 8480
rect 3108 8440 3114 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 2866 8304 2872 8356
rect 2924 8344 2930 8356
rect 3050 8344 3056 8356
rect 2924 8316 3056 8344
rect 2924 8304 2930 8316
rect 3050 8304 3056 8316
rect 3108 8304 3114 8356
rect 10042 8344 10048 8356
rect 10003 8316 10048 8344
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 1104 8186 10856 8208
rect 1104 8134 2582 8186
rect 2634 8134 2646 8186
rect 2698 8134 2710 8186
rect 2762 8134 2774 8186
rect 2826 8134 2838 8186
rect 2890 8134 5846 8186
rect 5898 8134 5910 8186
rect 5962 8134 5974 8186
rect 6026 8134 6038 8186
rect 6090 8134 6102 8186
rect 6154 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 9238 8186
rect 9290 8134 9302 8186
rect 9354 8134 9366 8186
rect 9418 8134 10856 8186
rect 1104 8112 10856 8134
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 5350 8072 5356 8084
rect 2915 8044 5356 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 2222 7936 2228 7948
rect 1719 7908 2228 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 2682 7868 2688 7880
rect 1636 7840 2688 7868
rect 1636 7828 1642 7840
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 3878 7828 3884 7880
rect 3936 7868 3942 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3936 7840 3985 7868
rect 3936 7828 3942 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 3789 7735 3847 7741
rect 3789 7701 3801 7735
rect 3835 7732 3847 7735
rect 9858 7732 9864 7744
rect 3835 7704 9864 7732
rect 3835 7701 3847 7704
rect 3789 7695 3847 7701
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 1104 7642 10856 7664
rect 1104 7590 4214 7642
rect 4266 7590 4278 7642
rect 4330 7590 4342 7642
rect 4394 7590 4406 7642
rect 4458 7590 4470 7642
rect 4522 7590 7478 7642
rect 7530 7590 7542 7642
rect 7594 7590 7606 7642
rect 7658 7590 7670 7642
rect 7722 7590 7734 7642
rect 7786 7590 10856 7642
rect 1104 7568 10856 7590
rect 2961 7531 3019 7537
rect 2961 7497 2973 7531
rect 3007 7528 3019 7531
rect 3510 7528 3516 7540
rect 3007 7500 3516 7528
rect 3007 7497 3019 7500
rect 2961 7491 3019 7497
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 3697 7531 3755 7537
rect 3697 7497 3709 7531
rect 3743 7528 3755 7531
rect 3786 7528 3792 7540
rect 3743 7500 3792 7528
rect 3743 7497 3755 7500
rect 3697 7491 3755 7497
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 2682 7420 2688 7472
rect 2740 7460 2746 7472
rect 2740 7432 4476 7460
rect 2740 7420 2746 7432
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2130 7352 2136 7404
rect 2188 7392 2194 7404
rect 2869 7395 2927 7401
rect 2188 7364 2233 7392
rect 2188 7352 2194 7364
rect 2869 7361 2881 7395
rect 2915 7361 2927 7395
rect 3602 7392 3608 7404
rect 3563 7364 3608 7392
rect 2869 7355 2927 7361
rect 2884 7324 2912 7355
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 4448 7401 4476 7432
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 9858 7392 9864 7404
rect 9819 7364 9864 7392
rect 4433 7355 4491 7361
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 2958 7324 2964 7336
rect 2884 7296 2964 7324
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 2406 7188 2412 7200
rect 2363 7160 2412 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 4249 7191 4307 7197
rect 4249 7157 4261 7191
rect 4295 7188 4307 7191
rect 9858 7188 9864 7200
rect 4295 7160 9864 7188
rect 4295 7157 4307 7160
rect 4249 7151 4307 7157
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10042 7188 10048 7200
rect 10003 7160 10048 7188
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 1104 7098 10856 7120
rect 1104 7046 2582 7098
rect 2634 7046 2646 7098
rect 2698 7046 2710 7098
rect 2762 7046 2774 7098
rect 2826 7046 2838 7098
rect 2890 7046 5846 7098
rect 5898 7046 5910 7098
rect 5962 7046 5974 7098
rect 6026 7046 6038 7098
rect 6090 7046 6102 7098
rect 6154 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 9238 7098
rect 9290 7046 9302 7098
rect 9354 7046 9366 7098
rect 9418 7046 10856 7098
rect 1104 7024 10856 7046
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6848 3019 6851
rect 3142 6848 3148 6860
rect 3007 6820 3148 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6848 4491 6851
rect 4614 6848 4620 6860
rect 4479 6820 4620 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 1762 6780 1768 6792
rect 1723 6752 1768 6780
rect 1762 6740 1768 6752
rect 1820 6740 1826 6792
rect 1946 6780 1952 6792
rect 1907 6752 1952 6780
rect 1946 6740 1952 6752
rect 2004 6780 2010 6792
rect 2130 6780 2136 6792
rect 2004 6752 2136 6780
rect 2004 6740 2010 6752
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2498 6740 2504 6792
rect 2556 6780 2562 6792
rect 2593 6783 2651 6789
rect 2593 6780 2605 6783
rect 2556 6752 2605 6780
rect 2556 6740 2562 6752
rect 2593 6749 2605 6752
rect 2639 6749 2651 6783
rect 2593 6743 2651 6749
rect 2777 6783 2835 6789
rect 2777 6749 2789 6783
rect 2823 6749 2835 6783
rect 9858 6780 9864 6792
rect 9819 6752 9864 6780
rect 2777 6743 2835 6749
rect 2148 6712 2176 6740
rect 2792 6712 2820 6743
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 2148 6684 2820 6712
rect 3142 6672 3148 6724
rect 3200 6712 3206 6724
rect 4249 6715 4307 6721
rect 4249 6712 4261 6715
rect 3200 6684 4261 6712
rect 3200 6672 3206 6684
rect 4249 6681 4261 6684
rect 4295 6681 4307 6715
rect 4249 6675 4307 6681
rect 1670 6604 1676 6656
rect 1728 6644 1734 6656
rect 2133 6647 2191 6653
rect 2133 6644 2145 6647
rect 1728 6616 2145 6644
rect 1728 6604 1734 6616
rect 2133 6613 2145 6616
rect 2179 6613 2191 6647
rect 10042 6644 10048 6656
rect 10003 6616 10048 6644
rect 2133 6607 2191 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 1104 6554 10856 6576
rect 1104 6502 4214 6554
rect 4266 6502 4278 6554
rect 4330 6502 4342 6554
rect 4394 6502 4406 6554
rect 4458 6502 4470 6554
rect 4522 6502 7478 6554
rect 7530 6502 7542 6554
rect 7594 6502 7606 6554
rect 7658 6502 7670 6554
rect 7722 6502 7734 6554
rect 7786 6502 10856 6554
rect 1104 6480 10856 6502
rect 1854 6440 1860 6452
rect 1815 6412 1860 6440
rect 1854 6400 1860 6412
rect 1912 6400 1918 6452
rect 2590 6440 2596 6452
rect 2551 6412 2596 6440
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 3050 6332 3056 6384
rect 3108 6372 3114 6384
rect 3108 6344 3556 6372
rect 3108 6332 3114 6344
rect 1670 6304 1676 6316
rect 1631 6276 1676 6304
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 2406 6304 2412 6316
rect 2367 6276 2412 6304
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 3326 6304 3332 6316
rect 3287 6276 3332 6304
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 3528 6313 3556 6344
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 3697 6103 3755 6109
rect 3697 6069 3709 6103
rect 3743 6100 3755 6103
rect 9030 6100 9036 6112
rect 3743 6072 9036 6100
rect 3743 6069 3755 6072
rect 3697 6063 3755 6069
rect 9030 6060 9036 6072
rect 9088 6060 9094 6112
rect 1104 6010 10856 6032
rect 1104 5958 2582 6010
rect 2634 5958 2646 6010
rect 2698 5958 2710 6010
rect 2762 5958 2774 6010
rect 2826 5958 2838 6010
rect 2890 5958 5846 6010
rect 5898 5958 5910 6010
rect 5962 5958 5974 6010
rect 6026 5958 6038 6010
rect 6090 5958 6102 6010
rect 6154 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 9238 6010
rect 9290 5958 9302 6010
rect 9354 5958 9366 6010
rect 9418 5958 10856 6010
rect 1104 5936 10856 5958
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 2958 5896 2964 5908
rect 2915 5868 2964 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 4028 5868 4445 5896
rect 4028 5856 4034 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 3789 5831 3847 5837
rect 3789 5797 3801 5831
rect 3835 5797 3847 5831
rect 3789 5791 3847 5797
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5760 1731 5763
rect 3418 5760 3424 5772
rect 1719 5732 3424 5760
rect 1719 5729 1731 5732
rect 1673 5723 1731 5729
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 3804 5760 3832 5791
rect 3804 5732 9904 5760
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 2222 5652 2228 5704
rect 2280 5692 2286 5704
rect 2685 5695 2743 5701
rect 2685 5692 2697 5695
rect 2280 5664 2697 5692
rect 2280 5652 2286 5664
rect 2685 5661 2697 5664
rect 2731 5692 2743 5695
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 2731 5664 3985 5692
rect 2731 5661 2743 5664
rect 2685 5655 2743 5661
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 9876 5701 9904 5732
rect 4617 5695 4675 5701
rect 4617 5692 4629 5695
rect 4212 5664 4629 5692
rect 4212 5652 4218 5664
rect 4617 5661 4629 5664
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 10042 5556 10048 5568
rect 10003 5528 10048 5556
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 1104 5466 10856 5488
rect 1104 5414 4214 5466
rect 4266 5414 4278 5466
rect 4330 5414 4342 5466
rect 4394 5414 4406 5466
rect 4458 5414 4470 5466
rect 4522 5414 7478 5466
rect 7530 5414 7542 5466
rect 7594 5414 7606 5466
rect 7658 5414 7670 5466
rect 7722 5414 7734 5466
rect 7786 5414 10856 5466
rect 1104 5392 10856 5414
rect 2866 5352 2872 5364
rect 2827 5324 2872 5352
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 3421 5355 3479 5361
rect 3421 5352 3433 5355
rect 3292 5324 3433 5352
rect 3292 5312 3298 5324
rect 3421 5321 3433 5324
rect 3467 5321 3479 5355
rect 3421 5315 3479 5321
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 1360 5188 1409 5216
rect 1360 5176 1366 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1946 5176 1952 5228
rect 2004 5216 2010 5228
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 2004 5188 2697 5216
rect 2004 5176 2010 5188
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 3602 5216 3608 5228
rect 3563 5188 3608 5216
rect 2685 5179 2743 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4522 5216 4528 5228
rect 4483 5188 4528 5216
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 9030 5176 9036 5228
rect 9088 5216 9094 5228
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 9088 5188 9413 5216
rect 9088 5176 9094 5188
rect 9401 5185 9413 5188
rect 9447 5185 9459 5219
rect 9401 5179 9459 5185
rect 9861 5219 9919 5225
rect 9861 5185 9873 5219
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5148 1731 5151
rect 4706 5148 4712 5160
rect 1719 5120 4712 5148
rect 1719 5117 1731 5120
rect 1673 5111 1731 5117
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 9876 5148 9904 5179
rect 9232 5120 9904 5148
rect 9232 5089 9260 5120
rect 9217 5083 9275 5089
rect 9217 5049 9229 5083
rect 9263 5049 9275 5083
rect 9217 5043 9275 5049
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 9858 5012 9864 5024
rect 4387 4984 9864 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 10042 5012 10048 5024
rect 10003 4984 10048 5012
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 1104 4922 10856 4944
rect 1104 4870 2582 4922
rect 2634 4870 2646 4922
rect 2698 4870 2710 4922
rect 2762 4870 2774 4922
rect 2826 4870 2838 4922
rect 2890 4870 5846 4922
rect 5898 4870 5910 4922
rect 5962 4870 5974 4922
rect 6026 4870 6038 4922
rect 6090 4870 6102 4922
rect 6154 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 9238 4922
rect 9290 4870 9302 4922
rect 9354 4870 9366 4922
rect 9418 4870 10856 4922
rect 1104 4848 10856 4870
rect 1946 4808 1952 4820
rect 1907 4780 1952 4808
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 4522 4808 4528 4820
rect 2823 4780 4528 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 3694 4632 3700 4684
rect 3752 4672 3758 4684
rect 3789 4675 3847 4681
rect 3789 4672 3801 4675
rect 3752 4644 3801 4672
rect 3752 4632 3758 4644
rect 3789 4641 3801 4644
rect 3835 4672 3847 4675
rect 3878 4672 3884 4684
rect 3835 4644 3884 4672
rect 3835 4641 3847 4644
rect 3789 4635 3847 4641
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 1854 4604 1860 4616
rect 1811 4576 1860 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 1688 4536 1716 4567
rect 1854 4564 1860 4576
rect 1912 4564 1918 4616
rect 2498 4604 2504 4616
rect 2459 4576 2504 4604
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 2774 4604 2780 4616
rect 2639 4576 2780 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 2774 4564 2780 4576
rect 2832 4604 2838 4616
rect 3050 4604 3056 4616
rect 2832 4576 3056 4604
rect 2832 4564 2838 4576
rect 3050 4564 3056 4576
rect 3108 4604 3114 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3108 4576 3985 4604
rect 3108 4564 3114 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 4798 4604 4804 4616
rect 4759 4576 4804 4604
rect 3973 4567 4031 4573
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 9858 4604 9864 4616
rect 9819 4576 9864 4604
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 2314 4536 2320 4548
rect 1688 4508 2320 4536
rect 2314 4496 2320 4508
rect 2372 4536 2378 4548
rect 2682 4536 2688 4548
rect 2372 4508 2688 4536
rect 2372 4496 2378 4508
rect 2682 4496 2688 4508
rect 2740 4496 2746 4548
rect 4154 4536 4160 4548
rect 4115 4508 4160 4536
rect 4154 4496 4160 4508
rect 4212 4496 4218 4548
rect 4617 4471 4675 4477
rect 4617 4437 4629 4471
rect 4663 4468 4675 4471
rect 9858 4468 9864 4480
rect 4663 4440 9864 4468
rect 4663 4437 4675 4440
rect 4617 4431 4675 4437
rect 9858 4428 9864 4440
rect 9916 4428 9922 4480
rect 10042 4468 10048 4480
rect 10003 4440 10048 4468
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 1104 4378 10856 4400
rect 1104 4326 4214 4378
rect 4266 4326 4278 4378
rect 4330 4326 4342 4378
rect 4394 4326 4406 4378
rect 4458 4326 4470 4378
rect 4522 4326 7478 4378
rect 7530 4326 7542 4378
rect 7594 4326 7606 4378
rect 7658 4326 7670 4378
rect 7722 4326 7734 4378
rect 7786 4326 10856 4378
rect 1104 4304 10856 4326
rect 4617 4267 4675 4273
rect 4617 4233 4629 4267
rect 4663 4264 4675 4267
rect 4798 4264 4804 4276
rect 4663 4236 4804 4264
rect 4663 4233 4675 4236
rect 4617 4227 4675 4233
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 2792 4168 4476 4196
rect 2792 4140 2820 4168
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 2406 4128 2412 4140
rect 1443 4100 2412 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 3620 4137 3648 4168
rect 4448 4137 4476 4168
rect 2961 4131 3019 4137
rect 2832 4100 2877 4128
rect 2832 4088 2838 4100
rect 2961 4097 2973 4131
rect 3007 4128 3019 4131
rect 3605 4131 3663 4137
rect 3007 4100 3556 4128
rect 3007 4097 3019 4100
rect 2961 4091 3019 4097
rect 1762 4020 1768 4072
rect 1820 4060 1826 4072
rect 2593 4063 2651 4069
rect 2593 4060 2605 4063
rect 1820 4032 2605 4060
rect 1820 4020 1826 4032
rect 2593 4029 2605 4032
rect 2639 4029 2651 4063
rect 2593 4023 2651 4029
rect 2682 4020 2688 4072
rect 2740 4060 2746 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 2740 4032 3433 4060
rect 2740 4020 2746 4032
rect 3421 4029 3433 4032
rect 3467 4029 3479 4063
rect 3528 4060 3556 4100
rect 3605 4097 3617 4131
rect 3651 4097 3663 4131
rect 4433 4131 4491 4137
rect 3605 4091 3663 4097
rect 4172 4100 4384 4128
rect 4172 4060 4200 4100
rect 3528 4032 4200 4060
rect 4249 4063 4307 4069
rect 3421 4023 3479 4029
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 4356 4060 4384 4100
rect 4433 4097 4445 4131
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 5276 4060 5304 4091
rect 4356 4032 5304 4060
rect 4249 4023 4307 4029
rect 1210 3952 1216 4004
rect 1268 3992 1274 4004
rect 1581 3995 1639 4001
rect 1581 3992 1593 3995
rect 1268 3964 1593 3992
rect 1268 3952 1274 3964
rect 1581 3961 1593 3964
rect 1627 3961 1639 3995
rect 4264 3992 4292 4023
rect 1581 3955 1639 3961
rect 2746 3964 4292 3992
rect 2038 3884 2044 3936
rect 2096 3924 2102 3936
rect 2746 3924 2774 3964
rect 2096 3896 2774 3924
rect 3789 3927 3847 3933
rect 2096 3884 2102 3896
rect 3789 3893 3801 3927
rect 3835 3924 3847 3927
rect 4614 3924 4620 3936
rect 3835 3896 4620 3924
rect 3835 3893 3847 3896
rect 3789 3887 3847 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5074 3924 5080 3936
rect 5035 3896 5080 3924
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 1104 3834 10856 3856
rect 1104 3782 2582 3834
rect 2634 3782 2646 3834
rect 2698 3782 2710 3834
rect 2762 3782 2774 3834
rect 2826 3782 2838 3834
rect 2890 3782 5846 3834
rect 5898 3782 5910 3834
rect 5962 3782 5974 3834
rect 6026 3782 6038 3834
rect 6090 3782 6102 3834
rect 6154 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 9238 3834
rect 9290 3782 9302 3834
rect 9354 3782 9366 3834
rect 9418 3782 10856 3834
rect 1104 3760 10856 3782
rect 1397 3723 1455 3729
rect 1397 3689 1409 3723
rect 1443 3720 1455 3723
rect 2222 3720 2228 3732
rect 1443 3692 2228 3720
rect 1443 3689 1455 3692
rect 1397 3683 1455 3689
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 3789 3655 3847 3661
rect 3789 3621 3801 3655
rect 3835 3652 3847 3655
rect 5534 3652 5540 3664
rect 3835 3624 5540 3652
rect 3835 3621 3847 3624
rect 3789 3615 3847 3621
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 2406 3476 2412 3528
rect 2464 3516 2470 3528
rect 2501 3519 2559 3525
rect 2501 3516 2513 3519
rect 2464 3488 2513 3516
rect 2464 3476 2470 3488
rect 2501 3485 2513 3488
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3516 4031 3519
rect 4154 3516 4160 3528
rect 4019 3488 4160 3516
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4614 3516 4620 3528
rect 4575 3488 4620 3516
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 9858 3516 9864 3528
rect 9819 3488 9864 3516
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 9674 3448 9680 3460
rect 2746 3420 9680 3448
rect 2317 3383 2375 3389
rect 2317 3349 2329 3383
rect 2363 3380 2375 3383
rect 2746 3380 2774 3420
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 2363 3352 2774 3380
rect 4433 3383 4491 3389
rect 2363 3349 2375 3352
rect 2317 3343 2375 3349
rect 4433 3349 4445 3383
rect 4479 3380 4491 3383
rect 9858 3380 9864 3392
rect 4479 3352 9864 3380
rect 4479 3349 4491 3352
rect 4433 3343 4491 3349
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 10042 3380 10048 3392
rect 10003 3352 10048 3380
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 1104 3290 10856 3312
rect 1104 3238 4214 3290
rect 4266 3238 4278 3290
rect 4330 3238 4342 3290
rect 4394 3238 4406 3290
rect 4458 3238 4470 3290
rect 4522 3238 7478 3290
rect 7530 3238 7542 3290
rect 7594 3238 7606 3290
rect 7658 3238 7670 3290
rect 7722 3238 7734 3290
rect 7786 3238 10856 3290
rect 1104 3216 10856 3238
rect 1397 3179 1455 3185
rect 1397 3145 1409 3179
rect 1443 3176 1455 3179
rect 1670 3176 1676 3188
rect 1443 3148 1676 3176
rect 1443 3145 1455 3148
rect 1397 3139 1455 3145
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 2498 3136 2504 3188
rect 2556 3176 2562 3188
rect 2685 3179 2743 3185
rect 2685 3176 2697 3179
rect 2556 3148 2697 3176
rect 2556 3136 2562 3148
rect 2685 3145 2697 3148
rect 2731 3145 2743 3179
rect 3326 3176 3332 3188
rect 3287 3148 3332 3176
rect 2685 3139 2743 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1452 3012 1593 3040
rect 1452 3000 1458 3012
rect 1581 3009 1593 3012
rect 1627 3009 1639 3043
rect 2222 3040 2228 3052
rect 2183 3012 2228 3040
rect 1581 3003 1639 3009
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 2958 3040 2964 3052
rect 2915 3012 2964 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 3510 3040 3516 3052
rect 3471 3012 3516 3040
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 5074 3000 5080 3052
rect 5132 3040 5138 3052
rect 9125 3043 9183 3049
rect 9125 3040 9137 3043
rect 5132 3012 9137 3040
rect 5132 3000 5138 3012
rect 9125 3009 9137 3012
rect 9171 3009 9183 3043
rect 9858 3040 9864 3052
rect 9819 3012 9864 3040
rect 9125 3003 9183 3009
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 9309 2839 9367 2845
rect 9309 2805 9321 2839
rect 9355 2836 9367 2839
rect 9490 2836 9496 2848
rect 9355 2808 9496 2836
rect 9355 2805 9367 2808
rect 9309 2799 9367 2805
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 10042 2836 10048 2848
rect 10003 2808 10048 2836
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 1104 2746 10856 2768
rect 1104 2694 2582 2746
rect 2634 2694 2646 2746
rect 2698 2694 2710 2746
rect 2762 2694 2774 2746
rect 2826 2694 2838 2746
rect 2890 2694 5846 2746
rect 5898 2694 5910 2746
rect 5962 2694 5974 2746
rect 6026 2694 6038 2746
rect 6090 2694 6102 2746
rect 6154 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 9238 2746
rect 9290 2694 9302 2746
rect 9354 2694 9366 2746
rect 9418 2694 10856 2746
rect 1104 2672 10856 2694
rect 2041 2635 2099 2641
rect 2041 2601 2053 2635
rect 2087 2632 2099 2635
rect 2406 2632 2412 2644
rect 2087 2604 2412 2632
rect 2087 2601 2099 2604
rect 2041 2595 2099 2601
rect 2406 2592 2412 2604
rect 2464 2592 2470 2644
rect 3789 2635 3847 2641
rect 3789 2601 3801 2635
rect 3835 2632 3847 2635
rect 3878 2632 3884 2644
rect 3835 2604 3884 2632
rect 3835 2601 3847 2604
rect 3789 2595 3847 2601
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 1397 2567 1455 2573
rect 1397 2533 1409 2567
rect 1443 2533 1455 2567
rect 1397 2527 1455 2533
rect 1412 2496 1440 2527
rect 2314 2524 2320 2576
rect 2372 2564 2378 2576
rect 2685 2567 2743 2573
rect 2685 2564 2697 2567
rect 2372 2536 2697 2564
rect 2372 2524 2378 2536
rect 2685 2533 2697 2536
rect 2731 2533 2743 2567
rect 2685 2527 2743 2533
rect 3970 2524 3976 2576
rect 4028 2524 4034 2576
rect 3988 2496 4016 2524
rect 1412 2468 4016 2496
rect 1486 2388 1492 2440
rect 1544 2428 1550 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1544 2400 1593 2428
rect 1544 2388 1550 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2866 2428 2872 2440
rect 2271 2400 2728 2428
rect 2827 2400 2872 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2700 2360 2728 2400
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3970 2428 3976 2440
rect 3931 2400 3976 2428
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 4614 2428 4620 2440
rect 4575 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 5592 2400 9137 2428
rect 5592 2388 5598 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9732 2400 9873 2428
rect 9732 2388 9738 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 2774 2360 2780 2372
rect 2700 2332 2780 2360
rect 2774 2320 2780 2332
rect 2832 2320 2838 2372
rect 1762 2252 1768 2304
rect 1820 2292 1826 2304
rect 4433 2295 4491 2301
rect 4433 2292 4445 2295
rect 1820 2264 4445 2292
rect 1820 2252 1826 2264
rect 4433 2261 4445 2264
rect 4479 2261 4491 2295
rect 9306 2292 9312 2304
rect 9267 2264 9312 2292
rect 4433 2255 4491 2261
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 9582 2252 9588 2304
rect 9640 2292 9646 2304
rect 10045 2295 10103 2301
rect 10045 2292 10057 2295
rect 9640 2264 10057 2292
rect 9640 2252 9646 2264
rect 10045 2261 10057 2264
rect 10091 2261 10103 2295
rect 10045 2255 10103 2261
rect 1104 2202 10856 2224
rect 1104 2150 4214 2202
rect 4266 2150 4278 2202
rect 4330 2150 4342 2202
rect 4394 2150 4406 2202
rect 4458 2150 4470 2202
rect 4522 2150 7478 2202
rect 7530 2150 7542 2202
rect 7594 2150 7606 2202
rect 7658 2150 7670 2202
rect 7722 2150 7734 2202
rect 7786 2150 10856 2202
rect 1104 2128 10856 2150
rect 2866 1028 2872 1080
rect 2924 1068 2930 1080
rect 4614 1068 4620 1080
rect 2924 1040 4620 1068
rect 2924 1028 2930 1040
rect 4614 1028 4620 1040
rect 4672 1028 4678 1080
<< via1 >>
rect 2582 77766 2634 77818
rect 2646 77766 2698 77818
rect 2710 77766 2762 77818
rect 2774 77766 2826 77818
rect 2838 77766 2890 77818
rect 5846 77766 5898 77818
rect 5910 77766 5962 77818
rect 5974 77766 6026 77818
rect 6038 77766 6090 77818
rect 6102 77766 6154 77818
rect 9110 77766 9162 77818
rect 9174 77766 9226 77818
rect 9238 77766 9290 77818
rect 9302 77766 9354 77818
rect 9366 77766 9418 77818
rect 1400 77571 1452 77580
rect 1400 77537 1409 77571
rect 1409 77537 1443 77571
rect 1443 77537 1452 77571
rect 1400 77528 1452 77537
rect 3792 77528 3844 77580
rect 1768 77460 1820 77512
rect 2872 77503 2924 77512
rect 2872 77469 2881 77503
rect 2881 77469 2915 77503
rect 2915 77469 2924 77503
rect 2872 77460 2924 77469
rect 3976 77503 4028 77512
rect 3976 77469 3985 77503
rect 3985 77469 4019 77503
rect 4019 77469 4028 77503
rect 3976 77460 4028 77469
rect 4068 77460 4120 77512
rect 9404 77503 9456 77512
rect 9404 77469 9413 77503
rect 9413 77469 9447 77503
rect 9447 77469 9456 77503
rect 9404 77460 9456 77469
rect 9956 77503 10008 77512
rect 9956 77469 9965 77503
rect 9965 77469 9999 77503
rect 9999 77469 10008 77503
rect 9956 77460 10008 77469
rect 2228 77324 2280 77376
rect 3056 77324 3108 77376
rect 4068 77324 4120 77376
rect 8300 77324 8352 77376
rect 4214 77222 4266 77274
rect 4278 77222 4330 77274
rect 4342 77222 4394 77274
rect 4406 77222 4458 77274
rect 4470 77222 4522 77274
rect 7478 77222 7530 77274
rect 7542 77222 7594 77274
rect 7606 77222 7658 77274
rect 7670 77222 7722 77274
rect 7734 77222 7786 77274
rect 1308 76984 1360 77036
rect 1492 76984 1544 77036
rect 2964 77027 3016 77036
rect 2964 76993 2973 77027
rect 2973 76993 3007 77027
rect 3007 76993 3016 77027
rect 2964 76984 3016 76993
rect 3608 77027 3660 77036
rect 3608 76993 3617 77027
rect 3617 76993 3651 77027
rect 3651 76993 3660 77027
rect 3608 76984 3660 76993
rect 3884 76984 3936 77036
rect 9496 76984 9548 77036
rect 9588 76984 9640 77036
rect 2504 76848 2556 76900
rect 1400 76780 1452 76832
rect 2320 76780 2372 76832
rect 3148 76780 3200 76832
rect 3424 76823 3476 76832
rect 3424 76789 3433 76823
rect 3433 76789 3467 76823
rect 3467 76789 3476 76823
rect 3424 76780 3476 76789
rect 4068 76823 4120 76832
rect 4068 76789 4077 76823
rect 4077 76789 4111 76823
rect 4111 76789 4120 76823
rect 4068 76780 4120 76789
rect 9772 76780 9824 76832
rect 2582 76678 2634 76730
rect 2646 76678 2698 76730
rect 2710 76678 2762 76730
rect 2774 76678 2826 76730
rect 2838 76678 2890 76730
rect 5846 76678 5898 76730
rect 5910 76678 5962 76730
rect 5974 76678 6026 76730
rect 6038 76678 6090 76730
rect 6102 76678 6154 76730
rect 9110 76678 9162 76730
rect 9174 76678 9226 76730
rect 9238 76678 9290 76730
rect 9302 76678 9354 76730
rect 9366 76678 9418 76730
rect 1952 76551 2004 76560
rect 1952 76517 1961 76551
rect 1961 76517 1995 76551
rect 1995 76517 2004 76551
rect 1952 76508 2004 76517
rect 3792 76508 3844 76560
rect 2136 76440 2188 76492
rect 2044 76372 2096 76424
rect 2504 76415 2556 76424
rect 2504 76381 2513 76415
rect 2513 76381 2547 76415
rect 2547 76381 2556 76415
rect 2504 76372 2556 76381
rect 10140 76415 10192 76424
rect 10140 76381 10149 76415
rect 10149 76381 10183 76415
rect 10183 76381 10192 76415
rect 10140 76372 10192 76381
rect 2136 76304 2188 76356
rect 4068 76304 4120 76356
rect 3424 76236 3476 76288
rect 4214 76134 4266 76186
rect 4278 76134 4330 76186
rect 4342 76134 4394 76186
rect 4406 76134 4458 76186
rect 4470 76134 4522 76186
rect 7478 76134 7530 76186
rect 7542 76134 7594 76186
rect 7606 76134 7658 76186
rect 7670 76134 7722 76186
rect 7734 76134 7786 76186
rect 1676 76032 1728 76084
rect 1584 75939 1636 75948
rect 1584 75905 1593 75939
rect 1593 75905 1627 75939
rect 1627 75905 1636 75939
rect 1584 75896 1636 75905
rect 2596 76007 2648 76016
rect 2596 75973 2605 76007
rect 2605 75973 2639 76007
rect 2639 75973 2648 76007
rect 2596 75964 2648 75973
rect 3516 75964 3568 76016
rect 2504 75939 2556 75948
rect 2504 75905 2513 75939
rect 2513 75905 2547 75939
rect 2547 75905 2556 75939
rect 2504 75896 2556 75905
rect 3608 75939 3660 75948
rect 2044 75828 2096 75880
rect 3608 75905 3617 75939
rect 3617 75905 3651 75939
rect 3651 75905 3660 75939
rect 3608 75896 3660 75905
rect 10140 75939 10192 75948
rect 10140 75905 10149 75939
rect 10149 75905 10183 75939
rect 10183 75905 10192 75939
rect 10140 75896 10192 75905
rect 2136 75760 2188 75812
rect 2504 75760 2556 75812
rect 3424 75735 3476 75744
rect 3424 75701 3433 75735
rect 3433 75701 3467 75735
rect 3467 75701 3476 75735
rect 3424 75692 3476 75701
rect 2582 75590 2634 75642
rect 2646 75590 2698 75642
rect 2710 75590 2762 75642
rect 2774 75590 2826 75642
rect 2838 75590 2890 75642
rect 5846 75590 5898 75642
rect 5910 75590 5962 75642
rect 5974 75590 6026 75642
rect 6038 75590 6090 75642
rect 6102 75590 6154 75642
rect 9110 75590 9162 75642
rect 9174 75590 9226 75642
rect 9238 75590 9290 75642
rect 9302 75590 9354 75642
rect 9366 75590 9418 75642
rect 1860 75488 1912 75540
rect 2504 75463 2556 75472
rect 2504 75429 2513 75463
rect 2513 75429 2547 75463
rect 2547 75429 2556 75463
rect 2504 75420 2556 75429
rect 2228 75327 2280 75336
rect 2228 75293 2237 75327
rect 2237 75293 2271 75327
rect 2271 75293 2280 75327
rect 2228 75284 2280 75293
rect 3240 75327 3292 75336
rect 2136 75259 2188 75268
rect 2136 75225 2145 75259
rect 2145 75225 2179 75259
rect 2179 75225 2188 75259
rect 2136 75216 2188 75225
rect 2044 75148 2096 75200
rect 3240 75293 3249 75327
rect 3249 75293 3283 75327
rect 3283 75293 3292 75327
rect 3240 75284 3292 75293
rect 10140 75327 10192 75336
rect 10140 75293 10149 75327
rect 10149 75293 10183 75327
rect 10183 75293 10192 75327
rect 10140 75284 10192 75293
rect 4214 75046 4266 75098
rect 4278 75046 4330 75098
rect 4342 75046 4394 75098
rect 4406 75046 4458 75098
rect 4470 75046 4522 75098
rect 7478 75046 7530 75098
rect 7542 75046 7594 75098
rect 7606 75046 7658 75098
rect 7670 75046 7722 75098
rect 7734 75046 7786 75098
rect 2136 74944 2188 74996
rect 3976 74876 4028 74928
rect 2044 74808 2096 74860
rect 2964 74808 3016 74860
rect 8300 74740 8352 74792
rect 1492 74672 1544 74724
rect 1952 74647 2004 74656
rect 1952 74613 1961 74647
rect 1961 74613 1995 74647
rect 1995 74613 2004 74647
rect 1952 74604 2004 74613
rect 2582 74502 2634 74554
rect 2646 74502 2698 74554
rect 2710 74502 2762 74554
rect 2774 74502 2826 74554
rect 2838 74502 2890 74554
rect 5846 74502 5898 74554
rect 5910 74502 5962 74554
rect 5974 74502 6026 74554
rect 6038 74502 6090 74554
rect 6102 74502 6154 74554
rect 9110 74502 9162 74554
rect 9174 74502 9226 74554
rect 9238 74502 9290 74554
rect 9302 74502 9354 74554
rect 9366 74502 9418 74554
rect 2412 74332 2464 74384
rect 2044 74196 2096 74248
rect 2872 74196 2924 74248
rect 3240 74239 3292 74248
rect 3240 74205 3249 74239
rect 3249 74205 3283 74239
rect 3283 74205 3292 74239
rect 3240 74196 3292 74205
rect 10140 74239 10192 74248
rect 10140 74205 10149 74239
rect 10149 74205 10183 74239
rect 10183 74205 10192 74239
rect 10140 74196 10192 74205
rect 2136 74171 2188 74180
rect 2136 74137 2145 74171
rect 2145 74137 2179 74171
rect 2179 74137 2188 74171
rect 2136 74128 2188 74137
rect 3148 74128 3200 74180
rect 3240 74060 3292 74112
rect 4214 73958 4266 74010
rect 4278 73958 4330 74010
rect 4342 73958 4394 74010
rect 4406 73958 4458 74010
rect 4470 73958 4522 74010
rect 7478 73958 7530 74010
rect 7542 73958 7594 74010
rect 7606 73958 7658 74010
rect 7670 73958 7722 74010
rect 7734 73958 7786 74010
rect 1584 73763 1636 73772
rect 1584 73729 1593 73763
rect 1593 73729 1627 73763
rect 1627 73729 1636 73763
rect 1584 73720 1636 73729
rect 2228 73763 2280 73772
rect 2228 73729 2237 73763
rect 2237 73729 2271 73763
rect 2271 73729 2280 73763
rect 2228 73720 2280 73729
rect 10140 73763 10192 73772
rect 10140 73729 10149 73763
rect 10149 73729 10183 73763
rect 10183 73729 10192 73763
rect 10140 73720 10192 73729
rect 1216 73652 1268 73704
rect 3148 73584 3200 73636
rect 2044 73559 2096 73568
rect 2044 73525 2053 73559
rect 2053 73525 2087 73559
rect 2087 73525 2096 73559
rect 2044 73516 2096 73525
rect 2582 73414 2634 73466
rect 2646 73414 2698 73466
rect 2710 73414 2762 73466
rect 2774 73414 2826 73466
rect 2838 73414 2890 73466
rect 5846 73414 5898 73466
rect 5910 73414 5962 73466
rect 5974 73414 6026 73466
rect 6038 73414 6090 73466
rect 6102 73414 6154 73466
rect 9110 73414 9162 73466
rect 9174 73414 9226 73466
rect 9238 73414 9290 73466
rect 9302 73414 9354 73466
rect 9366 73414 9418 73466
rect 2136 73176 2188 73228
rect 2964 73108 3016 73160
rect 9956 73108 10008 73160
rect 1860 72972 1912 73024
rect 4712 72972 4764 73024
rect 4214 72870 4266 72922
rect 4278 72870 4330 72922
rect 4342 72870 4394 72922
rect 4406 72870 4458 72922
rect 4470 72870 4522 72922
rect 7478 72870 7530 72922
rect 7542 72870 7594 72922
rect 7606 72870 7658 72922
rect 7670 72870 7722 72922
rect 7734 72870 7786 72922
rect 1400 72632 1452 72684
rect 2228 72675 2280 72684
rect 2228 72641 2237 72675
rect 2237 72641 2271 72675
rect 2271 72641 2280 72675
rect 2228 72632 2280 72641
rect 2872 72675 2924 72684
rect 2872 72641 2881 72675
rect 2881 72641 2915 72675
rect 2915 72641 2924 72675
rect 2872 72632 2924 72641
rect 10140 72675 10192 72684
rect 10140 72641 10149 72675
rect 10149 72641 10183 72675
rect 10183 72641 10192 72675
rect 10140 72632 10192 72641
rect 3332 72496 3384 72548
rect 1492 72428 1544 72480
rect 2504 72428 2556 72480
rect 8300 72428 8352 72480
rect 2582 72326 2634 72378
rect 2646 72326 2698 72378
rect 2710 72326 2762 72378
rect 2774 72326 2826 72378
rect 2838 72326 2890 72378
rect 5846 72326 5898 72378
rect 5910 72326 5962 72378
rect 5974 72326 6026 72378
rect 6038 72326 6090 72378
rect 6102 72326 6154 72378
rect 9110 72326 9162 72378
rect 9174 72326 9226 72378
rect 9238 72326 9290 72378
rect 9302 72326 9354 72378
rect 9366 72326 9418 72378
rect 9956 72267 10008 72276
rect 9956 72233 9965 72267
rect 9965 72233 9999 72267
rect 9999 72233 10008 72267
rect 9956 72224 10008 72233
rect 664 72156 716 72208
rect 1216 72088 1268 72140
rect 1584 72063 1636 72072
rect 1584 72029 1593 72063
rect 1593 72029 1627 72063
rect 1627 72029 1636 72063
rect 1584 72020 1636 72029
rect 2136 72088 2188 72140
rect 2320 72063 2372 72072
rect 2320 72029 2329 72063
rect 2329 72029 2363 72063
rect 2363 72029 2372 72063
rect 2320 72020 2372 72029
rect 2872 72020 2924 72072
rect 10140 72063 10192 72072
rect 10140 72029 10149 72063
rect 10149 72029 10183 72063
rect 10183 72029 10192 72063
rect 10140 72020 10192 72029
rect 1860 71884 1912 71936
rect 4214 71782 4266 71834
rect 4278 71782 4330 71834
rect 4342 71782 4394 71834
rect 4406 71782 4458 71834
rect 4470 71782 4522 71834
rect 7478 71782 7530 71834
rect 7542 71782 7594 71834
rect 7606 71782 7658 71834
rect 7670 71782 7722 71834
rect 7734 71782 7786 71834
rect 1676 71655 1728 71664
rect 1676 71621 1685 71655
rect 1685 71621 1719 71655
rect 1719 71621 1728 71655
rect 1676 71612 1728 71621
rect 2228 71680 2280 71732
rect 2872 71680 2924 71732
rect 1676 71476 1728 71528
rect 2136 71612 2188 71664
rect 3424 71612 3476 71664
rect 2872 71587 2924 71596
rect 2872 71553 2886 71587
rect 2886 71553 2920 71587
rect 2920 71553 2924 71587
rect 10140 71587 10192 71596
rect 2872 71544 2924 71553
rect 10140 71553 10149 71587
rect 10149 71553 10183 71587
rect 10183 71553 10192 71587
rect 10140 71544 10192 71553
rect 8300 71476 8352 71528
rect 2964 71340 3016 71392
rect 3976 71340 4028 71392
rect 2582 71238 2634 71290
rect 2646 71238 2698 71290
rect 2710 71238 2762 71290
rect 2774 71238 2826 71290
rect 2838 71238 2890 71290
rect 5846 71238 5898 71290
rect 5910 71238 5962 71290
rect 5974 71238 6026 71290
rect 6038 71238 6090 71290
rect 6102 71238 6154 71290
rect 9110 71238 9162 71290
rect 9174 71238 9226 71290
rect 9238 71238 9290 71290
rect 9302 71238 9354 71290
rect 9366 71238 9418 71290
rect 2688 71068 2740 71120
rect 940 70932 992 70984
rect 2228 70975 2280 70984
rect 2228 70941 2237 70975
rect 2237 70941 2271 70975
rect 2271 70941 2280 70975
rect 2228 70932 2280 70941
rect 2964 70864 3016 70916
rect 3608 70864 3660 70916
rect 1124 70796 1176 70848
rect 1492 70796 1544 70848
rect 2320 70796 2372 70848
rect 4214 70694 4266 70746
rect 4278 70694 4330 70746
rect 4342 70694 4394 70746
rect 4406 70694 4458 70746
rect 4470 70694 4522 70746
rect 7478 70694 7530 70746
rect 7542 70694 7594 70746
rect 7606 70694 7658 70746
rect 7670 70694 7722 70746
rect 7734 70694 7786 70746
rect 3240 70524 3292 70576
rect 1584 70499 1636 70508
rect 1584 70465 1593 70499
rect 1593 70465 1627 70499
rect 1627 70465 1636 70499
rect 1584 70456 1636 70465
rect 2136 70456 2188 70508
rect 10140 70499 10192 70508
rect 10140 70465 10149 70499
rect 10149 70465 10183 70499
rect 10183 70465 10192 70499
rect 10140 70456 10192 70465
rect 1216 70388 1268 70440
rect 3240 70388 3292 70440
rect 2582 70150 2634 70202
rect 2646 70150 2698 70202
rect 2710 70150 2762 70202
rect 2774 70150 2826 70202
rect 2838 70150 2890 70202
rect 5846 70150 5898 70202
rect 5910 70150 5962 70202
rect 5974 70150 6026 70202
rect 6038 70150 6090 70202
rect 6102 70150 6154 70202
rect 9110 70150 9162 70202
rect 9174 70150 9226 70202
rect 9238 70150 9290 70202
rect 9302 70150 9354 70202
rect 9366 70150 9418 70202
rect 1308 70048 1360 70100
rect 1584 70048 1636 70100
rect 1584 69887 1636 69896
rect 1584 69853 1593 69887
rect 1593 69853 1627 69887
rect 1627 69853 1636 69887
rect 1584 69844 1636 69853
rect 1676 69844 1728 69896
rect 10140 69887 10192 69896
rect 10140 69853 10149 69887
rect 10149 69853 10183 69887
rect 10183 69853 10192 69887
rect 10140 69844 10192 69853
rect 1400 69751 1452 69760
rect 1400 69717 1409 69751
rect 1409 69717 1443 69751
rect 1443 69717 1452 69751
rect 1400 69708 1452 69717
rect 1768 69708 1820 69760
rect 9956 69751 10008 69760
rect 9956 69717 9965 69751
rect 9965 69717 9999 69751
rect 9999 69717 10008 69751
rect 9956 69708 10008 69717
rect 4214 69606 4266 69658
rect 4278 69606 4330 69658
rect 4342 69606 4394 69658
rect 4406 69606 4458 69658
rect 4470 69606 4522 69658
rect 7478 69606 7530 69658
rect 7542 69606 7594 69658
rect 7606 69606 7658 69658
rect 7670 69606 7722 69658
rect 7734 69606 7786 69658
rect 572 69436 624 69488
rect 1860 69436 1912 69488
rect 1584 69411 1636 69420
rect 1584 69377 1593 69411
rect 1593 69377 1627 69411
rect 1627 69377 1636 69411
rect 1584 69368 1636 69377
rect 2228 69411 2280 69420
rect 2228 69377 2237 69411
rect 2237 69377 2271 69411
rect 2271 69377 2280 69411
rect 2228 69368 2280 69377
rect 1400 69300 1452 69352
rect 1676 69300 1728 69352
rect 1400 69207 1452 69216
rect 1400 69173 1409 69207
rect 1409 69173 1443 69207
rect 1443 69173 1452 69207
rect 1400 69164 1452 69173
rect 1860 69164 1912 69216
rect 2582 69062 2634 69114
rect 2646 69062 2698 69114
rect 2710 69062 2762 69114
rect 2774 69062 2826 69114
rect 2838 69062 2890 69114
rect 5846 69062 5898 69114
rect 5910 69062 5962 69114
rect 5974 69062 6026 69114
rect 6038 69062 6090 69114
rect 6102 69062 6154 69114
rect 9110 69062 9162 69114
rect 9174 69062 9226 69114
rect 9238 69062 9290 69114
rect 9302 69062 9354 69114
rect 9366 69062 9418 69114
rect 4896 68960 4948 69012
rect 9956 68824 10008 68876
rect 1492 68756 1544 68808
rect 1308 68688 1360 68740
rect 1952 68756 2004 68808
rect 2228 68756 2280 68808
rect 2780 68756 2832 68808
rect 10140 68799 10192 68808
rect 10140 68765 10149 68799
rect 10149 68765 10183 68799
rect 10183 68765 10192 68799
rect 10140 68756 10192 68765
rect 2596 68688 2648 68740
rect 1492 68620 1544 68672
rect 9956 68663 10008 68672
rect 9956 68629 9965 68663
rect 9965 68629 9999 68663
rect 9999 68629 10008 68663
rect 9956 68620 10008 68629
rect 4214 68518 4266 68570
rect 4278 68518 4330 68570
rect 4342 68518 4394 68570
rect 4406 68518 4458 68570
rect 4470 68518 4522 68570
rect 7478 68518 7530 68570
rect 7542 68518 7594 68570
rect 7606 68518 7658 68570
rect 7670 68518 7722 68570
rect 7734 68518 7786 68570
rect 1308 68348 1360 68400
rect 2044 68416 2096 68468
rect 2596 68348 2648 68400
rect 3240 68348 3292 68400
rect 1952 68280 2004 68332
rect 2412 68280 2464 68332
rect 2964 68280 3016 68332
rect 10140 68323 10192 68332
rect 10140 68289 10149 68323
rect 10149 68289 10183 68323
rect 10183 68289 10192 68323
rect 10140 68280 10192 68289
rect 9956 68212 10008 68264
rect 4620 68144 4672 68196
rect 2412 68076 2464 68128
rect 9864 68076 9916 68128
rect 2582 67974 2634 68026
rect 2646 67974 2698 68026
rect 2710 67974 2762 68026
rect 2774 67974 2826 68026
rect 2838 67974 2890 68026
rect 5846 67974 5898 68026
rect 5910 67974 5962 68026
rect 5974 67974 6026 68026
rect 6038 67974 6090 68026
rect 6102 67974 6154 68026
rect 9110 67974 9162 68026
rect 9174 67974 9226 68026
rect 9238 67974 9290 68026
rect 9302 67974 9354 68026
rect 9366 67974 9418 68026
rect 2044 67804 2096 67856
rect 3700 67804 3752 67856
rect 1308 67736 1360 67788
rect 1584 67711 1636 67720
rect 1584 67677 1593 67711
rect 1593 67677 1627 67711
rect 1627 67677 1636 67711
rect 1584 67668 1636 67677
rect 940 67600 992 67652
rect 1492 67600 1544 67652
rect 9956 67736 10008 67788
rect 2504 67711 2556 67720
rect 2504 67677 2513 67711
rect 2513 67677 2547 67711
rect 2547 67677 2556 67711
rect 2504 67668 2556 67677
rect 3240 67668 3292 67720
rect 2872 67600 2924 67652
rect 4214 67430 4266 67482
rect 4278 67430 4330 67482
rect 4342 67430 4394 67482
rect 4406 67430 4458 67482
rect 4470 67430 4522 67482
rect 7478 67430 7530 67482
rect 7542 67430 7594 67482
rect 7606 67430 7658 67482
rect 7670 67430 7722 67482
rect 7734 67430 7786 67482
rect 9680 67328 9732 67380
rect 9956 67371 10008 67380
rect 9956 67337 9965 67371
rect 9965 67337 9999 67371
rect 9999 67337 10008 67371
rect 9956 67328 10008 67337
rect 2872 67303 2924 67312
rect 2872 67269 2881 67303
rect 2881 67269 2915 67303
rect 2915 67269 2924 67303
rect 2872 67260 2924 67269
rect 2780 67192 2832 67244
rect 3240 67192 3292 67244
rect 10140 67235 10192 67244
rect 10140 67201 10149 67235
rect 10149 67201 10183 67235
rect 10183 67201 10192 67235
rect 10140 67192 10192 67201
rect 1400 67167 1452 67176
rect 1400 67133 1409 67167
rect 1409 67133 1443 67167
rect 1443 67133 1452 67167
rect 1400 67124 1452 67133
rect 1676 67167 1728 67176
rect 1676 67133 1685 67167
rect 1685 67133 1719 67167
rect 1719 67133 1728 67167
rect 1676 67124 1728 67133
rect 8484 66988 8536 67040
rect 2582 66886 2634 66938
rect 2646 66886 2698 66938
rect 2710 66886 2762 66938
rect 2774 66886 2826 66938
rect 2838 66886 2890 66938
rect 5846 66886 5898 66938
rect 5910 66886 5962 66938
rect 5974 66886 6026 66938
rect 6038 66886 6090 66938
rect 6102 66886 6154 66938
rect 9110 66886 9162 66938
rect 9174 66886 9226 66938
rect 9238 66886 9290 66938
rect 9302 66886 9354 66938
rect 9366 66886 9418 66938
rect 9680 66784 9732 66836
rect 2964 66716 3016 66768
rect 848 66648 900 66700
rect 1400 66623 1452 66632
rect 1400 66589 1409 66623
rect 1409 66589 1443 66623
rect 1443 66589 1452 66623
rect 1400 66580 1452 66589
rect 2780 66623 2832 66632
rect 2780 66589 2789 66623
rect 2789 66589 2823 66623
rect 2823 66589 2832 66623
rect 2780 66580 2832 66589
rect 10140 66623 10192 66632
rect 10140 66589 10149 66623
rect 10149 66589 10183 66623
rect 10183 66589 10192 66623
rect 10140 66580 10192 66589
rect 4214 66342 4266 66394
rect 4278 66342 4330 66394
rect 4342 66342 4394 66394
rect 4406 66342 4458 66394
rect 4470 66342 4522 66394
rect 7478 66342 7530 66394
rect 7542 66342 7594 66394
rect 7606 66342 7658 66394
rect 7670 66342 7722 66394
rect 7734 66342 7786 66394
rect 3148 66240 3200 66292
rect 2872 66215 2924 66224
rect 2872 66181 2881 66215
rect 2881 66181 2915 66215
rect 2915 66181 2924 66215
rect 2872 66172 2924 66181
rect 204 66104 256 66156
rect 1400 66079 1452 66088
rect 1400 66045 1409 66079
rect 1409 66045 1443 66079
rect 1443 66045 1452 66079
rect 1400 66036 1452 66045
rect 3240 66104 3292 66156
rect 10140 66147 10192 66156
rect 10140 66113 10149 66147
rect 10149 66113 10183 66147
rect 10183 66113 10192 66147
rect 10140 66104 10192 66113
rect 9864 66036 9916 66088
rect 3240 65943 3292 65952
rect 3240 65909 3249 65943
rect 3249 65909 3283 65943
rect 3283 65909 3292 65943
rect 3240 65900 3292 65909
rect 8300 65900 8352 65952
rect 2582 65798 2634 65850
rect 2646 65798 2698 65850
rect 2710 65798 2762 65850
rect 2774 65798 2826 65850
rect 2838 65798 2890 65850
rect 5846 65798 5898 65850
rect 5910 65798 5962 65850
rect 5974 65798 6026 65850
rect 6038 65798 6090 65850
rect 6102 65798 6154 65850
rect 9110 65798 9162 65850
rect 9174 65798 9226 65850
rect 9238 65798 9290 65850
rect 9302 65798 9354 65850
rect 9366 65798 9418 65850
rect 3884 65628 3936 65680
rect 4988 65628 5040 65680
rect 664 65560 716 65612
rect 1124 65560 1176 65612
rect 1308 65560 1360 65612
rect 3148 65560 3200 65612
rect 480 65492 532 65544
rect 1216 65492 1268 65544
rect 1676 65535 1728 65544
rect 1676 65501 1685 65535
rect 1685 65501 1719 65535
rect 1719 65501 1728 65535
rect 1676 65492 1728 65501
rect 2504 65492 2556 65544
rect 4068 65492 4120 65544
rect 3976 65399 4028 65408
rect 3976 65365 3985 65399
rect 3985 65365 4019 65399
rect 4019 65365 4028 65399
rect 3976 65356 4028 65365
rect 4214 65254 4266 65306
rect 4278 65254 4330 65306
rect 4342 65254 4394 65306
rect 4406 65254 4458 65306
rect 4470 65254 4522 65306
rect 7478 65254 7530 65306
rect 7542 65254 7594 65306
rect 7606 65254 7658 65306
rect 7670 65254 7722 65306
rect 7734 65254 7786 65306
rect 1216 65152 1268 65204
rect 2044 65152 2096 65204
rect 3700 65084 3752 65136
rect 3976 65084 4028 65136
rect 2044 65016 2096 65068
rect 1584 64923 1636 64932
rect 1584 64889 1593 64923
rect 1593 64889 1627 64923
rect 1627 64889 1636 64923
rect 1584 64880 1636 64889
rect 3148 64948 3200 65000
rect 3424 65016 3476 65068
rect 10140 65059 10192 65068
rect 10140 65025 10149 65059
rect 10149 65025 10183 65059
rect 10183 65025 10192 65059
rect 10140 65016 10192 65025
rect 3700 64948 3752 65000
rect 3056 64923 3108 64932
rect 3056 64889 3065 64923
rect 3065 64889 3099 64923
rect 3099 64889 3108 64923
rect 3056 64880 3108 64889
rect 8392 64880 8444 64932
rect 1676 64812 1728 64864
rect 3332 64812 3384 64864
rect 2582 64710 2634 64762
rect 2646 64710 2698 64762
rect 2710 64710 2762 64762
rect 2774 64710 2826 64762
rect 2838 64710 2890 64762
rect 5846 64710 5898 64762
rect 5910 64710 5962 64762
rect 5974 64710 6026 64762
rect 6038 64710 6090 64762
rect 6102 64710 6154 64762
rect 9110 64710 9162 64762
rect 9174 64710 9226 64762
rect 9238 64710 9290 64762
rect 9302 64710 9354 64762
rect 9366 64710 9418 64762
rect 8300 64608 8352 64660
rect 4804 64540 4856 64592
rect 1032 64336 1084 64388
rect 10140 64447 10192 64456
rect 2964 64336 3016 64388
rect 10140 64413 10149 64447
rect 10149 64413 10183 64447
rect 10183 64413 10192 64447
rect 10140 64404 10192 64413
rect 3056 64268 3108 64320
rect 8300 64268 8352 64320
rect 4214 64166 4266 64218
rect 4278 64166 4330 64218
rect 4342 64166 4394 64218
rect 4406 64166 4458 64218
rect 4470 64166 4522 64218
rect 7478 64166 7530 64218
rect 7542 64166 7594 64218
rect 7606 64166 7658 64218
rect 7670 64166 7722 64218
rect 7734 64166 7786 64218
rect 2320 64064 2372 64116
rect 3056 63928 3108 63980
rect 2228 63860 2280 63912
rect 8392 63860 8444 63912
rect 5172 63724 5224 63776
rect 2582 63622 2634 63674
rect 2646 63622 2698 63674
rect 2710 63622 2762 63674
rect 2774 63622 2826 63674
rect 2838 63622 2890 63674
rect 5846 63622 5898 63674
rect 5910 63622 5962 63674
rect 5974 63622 6026 63674
rect 6038 63622 6090 63674
rect 6102 63622 6154 63674
rect 9110 63622 9162 63674
rect 9174 63622 9226 63674
rect 9238 63622 9290 63674
rect 9302 63622 9354 63674
rect 9366 63622 9418 63674
rect 1584 63248 1636 63300
rect 2228 63452 2280 63504
rect 3056 63452 3108 63504
rect 3148 63452 3200 63504
rect 3424 63452 3476 63504
rect 8300 63452 8352 63504
rect 2228 63359 2280 63368
rect 2228 63325 2237 63359
rect 2237 63325 2271 63359
rect 2271 63325 2280 63359
rect 2228 63316 2280 63325
rect 2412 63359 2464 63368
rect 2412 63325 2415 63359
rect 2415 63325 2464 63359
rect 2412 63316 2464 63325
rect 2872 63316 2924 63368
rect 3424 63316 3476 63368
rect 9312 63359 9364 63368
rect 9312 63325 9321 63359
rect 9321 63325 9355 63359
rect 9355 63325 9364 63359
rect 9312 63316 9364 63325
rect 9588 63359 9640 63368
rect 9588 63325 9597 63359
rect 9597 63325 9631 63359
rect 9631 63325 9640 63359
rect 9588 63316 9640 63325
rect 2688 63248 2740 63300
rect 2964 63248 3016 63300
rect 3332 63180 3384 63232
rect 4214 63078 4266 63130
rect 4278 63078 4330 63130
rect 4342 63078 4394 63130
rect 4406 63078 4458 63130
rect 4470 63078 4522 63130
rect 7478 63078 7530 63130
rect 7542 63078 7594 63130
rect 7606 63078 7658 63130
rect 7670 63078 7722 63130
rect 7734 63078 7786 63130
rect 1400 62976 1452 63028
rect 1584 62883 1636 62892
rect 1584 62849 1593 62883
rect 1593 62849 1627 62883
rect 1627 62849 1636 62883
rect 1584 62840 1636 62849
rect 2412 62840 2464 62892
rect 4988 62976 5040 63028
rect 2596 62908 2648 62960
rect 3332 62908 3384 62960
rect 3700 62908 3752 62960
rect 2688 62883 2740 62892
rect 2688 62849 2697 62883
rect 2697 62849 2731 62883
rect 2731 62849 2740 62883
rect 2688 62840 2740 62849
rect 2872 62883 2924 62892
rect 2872 62849 2881 62883
rect 2881 62849 2915 62883
rect 2915 62849 2924 62883
rect 2872 62840 2924 62849
rect 5356 62840 5408 62892
rect 10140 62883 10192 62892
rect 10140 62849 10149 62883
rect 10149 62849 10183 62883
rect 10183 62849 10192 62883
rect 10140 62840 10192 62849
rect 1400 62704 1452 62756
rect 1584 62704 1636 62756
rect 3700 62747 3752 62756
rect 3700 62713 3709 62747
rect 3709 62713 3743 62747
rect 3743 62713 3752 62747
rect 3700 62704 3752 62713
rect 1952 62679 2004 62688
rect 1952 62645 1961 62679
rect 1961 62645 1995 62679
rect 1995 62645 2004 62679
rect 1952 62636 2004 62645
rect 5264 62636 5316 62688
rect 2582 62534 2634 62586
rect 2646 62534 2698 62586
rect 2710 62534 2762 62586
rect 2774 62534 2826 62586
rect 2838 62534 2890 62586
rect 5846 62534 5898 62586
rect 5910 62534 5962 62586
rect 5974 62534 6026 62586
rect 6038 62534 6090 62586
rect 6102 62534 6154 62586
rect 9110 62534 9162 62586
rect 9174 62534 9226 62586
rect 9238 62534 9290 62586
rect 9302 62534 9354 62586
rect 9366 62534 9418 62586
rect 1952 62432 2004 62484
rect 3976 62432 4028 62484
rect 2412 62364 2464 62416
rect 2596 62364 2648 62416
rect 1952 62296 2004 62348
rect 2320 62296 2372 62348
rect 20 62228 72 62280
rect 572 62160 624 62212
rect 2412 62228 2464 62280
rect 10140 62271 10192 62280
rect 10140 62237 10149 62271
rect 10149 62237 10183 62271
rect 10183 62237 10192 62271
rect 10140 62228 10192 62237
rect 1584 62135 1636 62144
rect 1584 62101 1593 62135
rect 1593 62101 1627 62135
rect 1627 62101 1636 62135
rect 1584 62092 1636 62101
rect 2320 62135 2372 62144
rect 2320 62101 2329 62135
rect 2329 62101 2363 62135
rect 2363 62101 2372 62135
rect 2320 62092 2372 62101
rect 2780 62092 2832 62144
rect 8300 62092 8352 62144
rect 4214 61990 4266 62042
rect 4278 61990 4330 62042
rect 4342 61990 4394 62042
rect 4406 61990 4458 62042
rect 4470 61990 4522 62042
rect 7478 61990 7530 62042
rect 7542 61990 7594 62042
rect 7606 61990 7658 62042
rect 7670 61990 7722 62042
rect 7734 61990 7786 62042
rect 8300 61820 8352 61872
rect 1400 61616 1452 61668
rect 1676 61795 1728 61804
rect 1676 61761 1685 61795
rect 1685 61761 1719 61795
rect 1719 61761 1728 61795
rect 1676 61752 1728 61761
rect 2596 61752 2648 61804
rect 940 61548 992 61600
rect 1676 61548 1728 61600
rect 2044 61548 2096 61600
rect 2582 61446 2634 61498
rect 2646 61446 2698 61498
rect 2710 61446 2762 61498
rect 2774 61446 2826 61498
rect 2838 61446 2890 61498
rect 5846 61446 5898 61498
rect 5910 61446 5962 61498
rect 5974 61446 6026 61498
rect 6038 61446 6090 61498
rect 6102 61446 6154 61498
rect 9110 61446 9162 61498
rect 9174 61446 9226 61498
rect 9238 61446 9290 61498
rect 9302 61446 9354 61498
rect 9366 61446 9418 61498
rect 1216 61344 1268 61396
rect 1768 61344 1820 61396
rect 1032 61140 1084 61192
rect 10140 61183 10192 61192
rect 940 61072 992 61124
rect 10140 61149 10149 61183
rect 10149 61149 10183 61183
rect 10183 61149 10192 61183
rect 10140 61140 10192 61149
rect 1584 61047 1636 61056
rect 1584 61013 1593 61047
rect 1593 61013 1627 61047
rect 1627 61013 1636 61047
rect 1584 61004 1636 61013
rect 1952 61004 2004 61056
rect 2136 61004 2188 61056
rect 2320 61047 2372 61056
rect 2320 61013 2329 61047
rect 2329 61013 2363 61047
rect 2363 61013 2372 61047
rect 2320 61004 2372 61013
rect 2780 61004 2832 61056
rect 4214 60902 4266 60954
rect 4278 60902 4330 60954
rect 4342 60902 4394 60954
rect 4406 60902 4458 60954
rect 4470 60902 4522 60954
rect 7478 60902 7530 60954
rect 7542 60902 7594 60954
rect 7606 60902 7658 60954
rect 7670 60902 7722 60954
rect 7734 60902 7786 60954
rect 2780 60800 2832 60852
rect 2320 60732 2372 60784
rect 3056 60664 3108 60716
rect 3976 60664 4028 60716
rect 10140 60707 10192 60716
rect 10140 60673 10149 60707
rect 10149 60673 10183 60707
rect 10183 60673 10192 60707
rect 10140 60664 10192 60673
rect 1860 60596 1912 60648
rect 2964 60596 3016 60648
rect 1400 60528 1452 60580
rect 2780 60528 2832 60580
rect 1860 60460 1912 60512
rect 6920 60460 6972 60512
rect 2582 60358 2634 60410
rect 2646 60358 2698 60410
rect 2710 60358 2762 60410
rect 2774 60358 2826 60410
rect 2838 60358 2890 60410
rect 5846 60358 5898 60410
rect 5910 60358 5962 60410
rect 5974 60358 6026 60410
rect 6038 60358 6090 60410
rect 6102 60358 6154 60410
rect 9110 60358 9162 60410
rect 9174 60358 9226 60410
rect 9238 60358 9290 60410
rect 9302 60358 9354 60410
rect 9366 60358 9418 60410
rect 3148 60256 3200 60308
rect 2964 60188 3016 60240
rect 3148 60120 3200 60172
rect 756 60052 808 60104
rect 112 59984 164 60036
rect 2964 60052 3016 60104
rect 1584 59959 1636 59968
rect 1584 59925 1593 59959
rect 1593 59925 1627 59959
rect 1627 59925 1636 59959
rect 1584 59916 1636 59925
rect 2320 59959 2372 59968
rect 2320 59925 2329 59959
rect 2329 59925 2363 59959
rect 2363 59925 2372 59959
rect 2320 59916 2372 59925
rect 4214 59814 4266 59866
rect 4278 59814 4330 59866
rect 4342 59814 4394 59866
rect 4406 59814 4458 59866
rect 4470 59814 4522 59866
rect 7478 59814 7530 59866
rect 7542 59814 7594 59866
rect 7606 59814 7658 59866
rect 7670 59814 7722 59866
rect 7734 59814 7786 59866
rect 388 59576 440 59628
rect 8300 59576 8352 59628
rect 9312 59551 9364 59560
rect 9312 59517 9321 59551
rect 9321 59517 9355 59551
rect 9355 59517 9364 59551
rect 9312 59508 9364 59517
rect 1400 59372 1452 59424
rect 2582 59270 2634 59322
rect 2646 59270 2698 59322
rect 2710 59270 2762 59322
rect 2774 59270 2826 59322
rect 2838 59270 2890 59322
rect 5846 59270 5898 59322
rect 5910 59270 5962 59322
rect 5974 59270 6026 59322
rect 6038 59270 6090 59322
rect 6102 59270 6154 59322
rect 9110 59270 9162 59322
rect 9174 59270 9226 59322
rect 9238 59270 9290 59322
rect 9302 59270 9354 59322
rect 9366 59270 9418 59322
rect 480 58964 532 59016
rect 2780 58964 2832 59016
rect 5080 58964 5132 59016
rect 10140 59007 10192 59016
rect 10140 58973 10149 59007
rect 10149 58973 10183 59007
rect 10183 58973 10192 59007
rect 10140 58964 10192 58973
rect 1584 58871 1636 58880
rect 1584 58837 1593 58871
rect 1593 58837 1627 58871
rect 1627 58837 1636 58871
rect 1584 58828 1636 58837
rect 2320 58871 2372 58880
rect 2320 58837 2329 58871
rect 2329 58837 2363 58871
rect 2363 58837 2372 58871
rect 2320 58828 2372 58837
rect 3056 58871 3108 58880
rect 3056 58837 3065 58871
rect 3065 58837 3099 58871
rect 3099 58837 3108 58871
rect 3056 58828 3108 58837
rect 9956 58871 10008 58880
rect 9956 58837 9965 58871
rect 9965 58837 9999 58871
rect 9999 58837 10008 58871
rect 9956 58828 10008 58837
rect 4214 58726 4266 58778
rect 4278 58726 4330 58778
rect 4342 58726 4394 58778
rect 4406 58726 4458 58778
rect 4470 58726 4522 58778
rect 7478 58726 7530 58778
rect 7542 58726 7594 58778
rect 7606 58726 7658 58778
rect 7670 58726 7722 58778
rect 7734 58726 7786 58778
rect 1492 58556 1544 58608
rect 2688 58624 2740 58676
rect 2780 58624 2832 58676
rect 3056 58624 3108 58676
rect 2688 58488 2740 58540
rect 10140 58531 10192 58540
rect 10140 58497 10149 58531
rect 10149 58497 10183 58531
rect 10183 58497 10192 58531
rect 10140 58488 10192 58497
rect 9588 58352 9640 58404
rect 1124 58284 1176 58336
rect 9680 58284 9732 58336
rect 2582 58182 2634 58234
rect 2646 58182 2698 58234
rect 2710 58182 2762 58234
rect 2774 58182 2826 58234
rect 2838 58182 2890 58234
rect 5846 58182 5898 58234
rect 5910 58182 5962 58234
rect 5974 58182 6026 58234
rect 6038 58182 6090 58234
rect 6102 58182 6154 58234
rect 9110 58182 9162 58234
rect 9174 58182 9226 58234
rect 9238 58182 9290 58234
rect 9302 58182 9354 58234
rect 9366 58182 9418 58234
rect 1492 57944 1544 57996
rect 1676 57919 1728 57928
rect 1676 57885 1685 57919
rect 1685 57885 1719 57919
rect 1719 57885 1728 57919
rect 1676 57876 1728 57885
rect 2320 58012 2372 58064
rect 2688 58012 2740 58064
rect 2596 57876 2648 57928
rect 2780 57876 2832 57928
rect 1492 57740 1544 57792
rect 1676 57740 1728 57792
rect 1860 57740 1912 57792
rect 2596 57740 2648 57792
rect 4214 57638 4266 57690
rect 4278 57638 4330 57690
rect 4342 57638 4394 57690
rect 4406 57638 4458 57690
rect 4470 57638 4522 57690
rect 7478 57638 7530 57690
rect 7542 57638 7594 57690
rect 7606 57638 7658 57690
rect 7670 57638 7722 57690
rect 7734 57638 7786 57690
rect 2412 57536 2464 57588
rect 3332 57536 3384 57588
rect 296 57400 348 57452
rect 1308 57332 1360 57384
rect 3056 57400 3108 57452
rect 3148 57400 3200 57452
rect 9496 57332 9548 57384
rect 2504 57264 2556 57316
rect 2780 57264 2832 57316
rect 3332 57264 3384 57316
rect 6276 57264 6328 57316
rect 1492 57196 1544 57248
rect 2412 57196 2464 57248
rect 3056 57239 3108 57248
rect 3056 57205 3065 57239
rect 3065 57205 3099 57239
rect 3099 57205 3108 57239
rect 3056 57196 3108 57205
rect 2582 57094 2634 57146
rect 2646 57094 2698 57146
rect 2710 57094 2762 57146
rect 2774 57094 2826 57146
rect 2838 57094 2890 57146
rect 5846 57094 5898 57146
rect 5910 57094 5962 57146
rect 5974 57094 6026 57146
rect 6038 57094 6090 57146
rect 6102 57094 6154 57146
rect 9110 57094 9162 57146
rect 9174 57094 9226 57146
rect 9238 57094 9290 57146
rect 9302 57094 9354 57146
rect 9366 57094 9418 57146
rect 2964 57035 3016 57044
rect 1492 56924 1544 56976
rect 2964 57001 2973 57035
rect 2973 57001 3007 57035
rect 3007 57001 3016 57035
rect 2964 56992 3016 57001
rect 4068 56992 4120 57044
rect 9956 56924 10008 56976
rect 2596 56856 2648 56908
rect 6460 56856 6512 56908
rect 2688 56831 2740 56840
rect 2688 56797 2697 56831
rect 2697 56797 2731 56831
rect 2731 56797 2740 56831
rect 2688 56788 2740 56797
rect 3976 56831 4028 56840
rect 2504 56720 2556 56772
rect 1768 56652 1820 56704
rect 2320 56652 2372 56704
rect 3976 56797 3985 56831
rect 3985 56797 4019 56831
rect 4019 56797 4028 56831
rect 3976 56788 4028 56797
rect 9312 56831 9364 56840
rect 9312 56797 9321 56831
rect 9321 56797 9355 56831
rect 9355 56797 9364 56831
rect 9312 56788 9364 56797
rect 4214 56550 4266 56602
rect 4278 56550 4330 56602
rect 4342 56550 4394 56602
rect 4406 56550 4458 56602
rect 4470 56550 4522 56602
rect 7478 56550 7530 56602
rect 7542 56550 7594 56602
rect 7606 56550 7658 56602
rect 7670 56550 7722 56602
rect 7734 56550 7786 56602
rect 3976 56448 4028 56500
rect 2780 56380 2832 56432
rect 3332 56380 3384 56432
rect 848 56312 900 56364
rect 1216 56312 1268 56364
rect 2964 56312 3016 56364
rect 4160 56380 4212 56432
rect 4712 56380 4764 56432
rect 4988 56380 5040 56432
rect 2872 56244 2924 56296
rect 8576 56244 8628 56296
rect 3332 56176 3384 56228
rect 9956 56151 10008 56160
rect 9956 56117 9965 56151
rect 9965 56117 9999 56151
rect 9999 56117 10008 56151
rect 9956 56108 10008 56117
rect 848 56040 900 56092
rect 572 55904 624 55956
rect 848 55904 900 55956
rect 2582 56006 2634 56058
rect 2646 56006 2698 56058
rect 2710 56006 2762 56058
rect 2774 56006 2826 56058
rect 2838 56006 2890 56058
rect 5846 56006 5898 56058
rect 5910 56006 5962 56058
rect 5974 56006 6026 56058
rect 6038 56006 6090 56058
rect 6102 56006 6154 56058
rect 9110 56006 9162 56058
rect 9174 56006 9226 56058
rect 9238 56006 9290 56058
rect 9302 56006 9354 56058
rect 9366 56006 9418 56058
rect 3148 55904 3200 55956
rect 3332 55836 3384 55888
rect 664 55700 716 55752
rect 2320 55700 2372 55752
rect 3332 55700 3384 55752
rect 3976 55836 4028 55888
rect 5448 55768 5500 55820
rect 4160 55700 4212 55752
rect 4620 55743 4672 55752
rect 4620 55709 4629 55743
rect 4629 55709 4663 55743
rect 4663 55709 4672 55743
rect 4620 55700 4672 55709
rect 9312 55743 9364 55752
rect 9312 55709 9321 55743
rect 9321 55709 9355 55743
rect 9355 55709 9364 55743
rect 9312 55700 9364 55709
rect 6368 55632 6420 55684
rect 3148 55564 3200 55616
rect 3424 55564 3476 55616
rect 10140 55564 10192 55616
rect 4214 55462 4266 55514
rect 4278 55462 4330 55514
rect 4342 55462 4394 55514
rect 4406 55462 4458 55514
rect 4470 55462 4522 55514
rect 7478 55462 7530 55514
rect 7542 55462 7594 55514
rect 7606 55462 7658 55514
rect 7670 55462 7722 55514
rect 7734 55462 7786 55514
rect 1676 55360 1728 55412
rect 1768 55360 1820 55412
rect 1952 55360 2004 55412
rect 3424 55403 3476 55412
rect 3424 55369 3433 55403
rect 3433 55369 3467 55403
rect 3467 55369 3476 55403
rect 3424 55360 3476 55369
rect 5540 55360 5592 55412
rect 9680 55360 9732 55412
rect 2504 55267 2556 55276
rect 2504 55233 2513 55267
rect 2513 55233 2547 55267
rect 2547 55233 2556 55267
rect 2504 55224 2556 55233
rect 4160 55224 4212 55276
rect 9496 55224 9548 55276
rect 1584 55156 1636 55208
rect 2320 55156 2372 55208
rect 2596 55156 2648 55208
rect 2964 55156 3016 55208
rect 2872 55088 2924 55140
rect 1952 55063 2004 55072
rect 1952 55029 1961 55063
rect 1961 55029 1995 55063
rect 1995 55029 2004 55063
rect 1952 55020 2004 55029
rect 2504 55020 2556 55072
rect 3424 55020 3476 55072
rect 6552 55020 6604 55072
rect 2582 54918 2634 54970
rect 2646 54918 2698 54970
rect 2710 54918 2762 54970
rect 2774 54918 2826 54970
rect 2838 54918 2890 54970
rect 5846 54918 5898 54970
rect 5910 54918 5962 54970
rect 5974 54918 6026 54970
rect 6038 54918 6090 54970
rect 6102 54918 6154 54970
rect 9110 54918 9162 54970
rect 9174 54918 9226 54970
rect 9238 54918 9290 54970
rect 9302 54918 9354 54970
rect 9366 54918 9418 54970
rect 5540 54816 5592 54868
rect 8300 54680 8352 54732
rect 1492 54612 1544 54664
rect 2320 54612 2372 54664
rect 6644 54612 6696 54664
rect 10140 54655 10192 54664
rect 10140 54621 10149 54655
rect 10149 54621 10183 54655
rect 10183 54621 10192 54655
rect 10140 54612 10192 54621
rect 1584 54587 1636 54596
rect 1584 54553 1593 54587
rect 1593 54553 1627 54587
rect 1627 54553 1636 54587
rect 1584 54544 1636 54553
rect 2320 54476 2372 54528
rect 2780 54476 2832 54528
rect 9864 54476 9916 54528
rect 4214 54374 4266 54426
rect 4278 54374 4330 54426
rect 4342 54374 4394 54426
rect 4406 54374 4458 54426
rect 4470 54374 4522 54426
rect 7478 54374 7530 54426
rect 7542 54374 7594 54426
rect 7606 54374 7658 54426
rect 7670 54374 7722 54426
rect 7734 54374 7786 54426
rect 3056 54272 3108 54324
rect 2320 54204 2372 54256
rect 10232 54204 10284 54256
rect 3056 54179 3108 54188
rect 3056 54145 3065 54179
rect 3065 54145 3099 54179
rect 3099 54145 3108 54179
rect 3056 54136 3108 54145
rect 9864 54179 9916 54188
rect 9864 54145 9873 54179
rect 9873 54145 9907 54179
rect 9907 54145 9916 54179
rect 9864 54136 9916 54145
rect 4436 54068 4488 54120
rect 4528 54000 4580 54052
rect 10048 54043 10100 54052
rect 10048 54009 10057 54043
rect 10057 54009 10091 54043
rect 10091 54009 10100 54043
rect 10048 54000 10100 54009
rect 1400 53932 1452 53984
rect 2320 53975 2372 53984
rect 2320 53941 2329 53975
rect 2329 53941 2363 53975
rect 2363 53941 2372 53975
rect 2320 53932 2372 53941
rect 2582 53830 2634 53882
rect 2646 53830 2698 53882
rect 2710 53830 2762 53882
rect 2774 53830 2826 53882
rect 2838 53830 2890 53882
rect 5846 53830 5898 53882
rect 5910 53830 5962 53882
rect 5974 53830 6026 53882
rect 6038 53830 6090 53882
rect 6102 53830 6154 53882
rect 9110 53830 9162 53882
rect 9174 53830 9226 53882
rect 9238 53830 9290 53882
rect 9302 53830 9354 53882
rect 9366 53830 9418 53882
rect 1492 53524 1544 53576
rect 9956 53524 10008 53576
rect 1584 53431 1636 53440
rect 1584 53397 1593 53431
rect 1593 53397 1627 53431
rect 1627 53397 1636 53431
rect 1584 53388 1636 53397
rect 10048 53431 10100 53440
rect 10048 53397 10057 53431
rect 10057 53397 10091 53431
rect 10091 53397 10100 53431
rect 10048 53388 10100 53397
rect 4214 53286 4266 53338
rect 4278 53286 4330 53338
rect 4342 53286 4394 53338
rect 4406 53286 4458 53338
rect 4470 53286 4522 53338
rect 7478 53286 7530 53338
rect 7542 53286 7594 53338
rect 7606 53286 7658 53338
rect 7670 53286 7722 53338
rect 7734 53286 7786 53338
rect 3056 53184 3108 53236
rect 3516 53116 3568 53168
rect 3976 53116 4028 53168
rect 5356 53116 5408 53168
rect 6184 53116 6236 53168
rect 2320 53091 2372 53100
rect 2320 53057 2329 53091
rect 2329 53057 2363 53091
rect 2363 53057 2372 53091
rect 2320 53048 2372 53057
rect 2964 53048 3016 53100
rect 2504 52980 2556 53032
rect 3056 53023 3108 53032
rect 3056 52989 3065 53023
rect 3065 52989 3099 53023
rect 3099 52989 3108 53023
rect 3056 52980 3108 52989
rect 3332 52980 3384 53032
rect 5080 52912 5132 52964
rect 1400 52844 1452 52896
rect 10048 52887 10100 52896
rect 10048 52853 10057 52887
rect 10057 52853 10091 52887
rect 10091 52853 10100 52887
rect 10048 52844 10100 52853
rect 2582 52742 2634 52794
rect 2646 52742 2698 52794
rect 2710 52742 2762 52794
rect 2774 52742 2826 52794
rect 2838 52742 2890 52794
rect 5846 52742 5898 52794
rect 5910 52742 5962 52794
rect 5974 52742 6026 52794
rect 6038 52742 6090 52794
rect 6102 52742 6154 52794
rect 9110 52742 9162 52794
rect 9174 52742 9226 52794
rect 9238 52742 9290 52794
rect 9302 52742 9354 52794
rect 9366 52742 9418 52794
rect 2320 52615 2372 52624
rect 2320 52581 2329 52615
rect 2329 52581 2363 52615
rect 2363 52581 2372 52615
rect 2320 52572 2372 52581
rect 5632 52436 5684 52488
rect 10140 52479 10192 52488
rect 10140 52445 10149 52479
rect 10149 52445 10183 52479
rect 10183 52445 10192 52479
rect 10140 52436 10192 52445
rect 2596 52368 2648 52420
rect 1492 52300 1544 52352
rect 9864 52300 9916 52352
rect 4214 52198 4266 52250
rect 4278 52198 4330 52250
rect 4342 52198 4394 52250
rect 4406 52198 4458 52250
rect 4470 52198 4522 52250
rect 7478 52198 7530 52250
rect 7542 52198 7594 52250
rect 7606 52198 7658 52250
rect 7670 52198 7722 52250
rect 7734 52198 7786 52250
rect 2228 52139 2280 52148
rect 2228 52105 2237 52139
rect 2237 52105 2271 52139
rect 2271 52105 2280 52139
rect 2228 52096 2280 52105
rect 10140 52096 10192 52148
rect 2228 51960 2280 52012
rect 2412 52003 2464 52012
rect 2412 51969 2421 52003
rect 2421 51969 2455 52003
rect 2455 51969 2464 52003
rect 2412 51960 2464 51969
rect 2964 51960 3016 52012
rect 3332 51960 3384 52012
rect 9864 52003 9916 52012
rect 9864 51969 9873 52003
rect 9873 51969 9907 52003
rect 9907 51969 9916 52003
rect 9864 51960 9916 51969
rect 2504 51892 2556 51944
rect 2964 51824 3016 51876
rect 10140 51824 10192 51876
rect 1584 51799 1636 51808
rect 1584 51765 1593 51799
rect 1593 51765 1627 51799
rect 1627 51765 1636 51799
rect 1584 51756 1636 51765
rect 10048 51799 10100 51808
rect 10048 51765 10057 51799
rect 10057 51765 10091 51799
rect 10091 51765 10100 51799
rect 10048 51756 10100 51765
rect 2582 51654 2634 51706
rect 2646 51654 2698 51706
rect 2710 51654 2762 51706
rect 2774 51654 2826 51706
rect 2838 51654 2890 51706
rect 5846 51654 5898 51706
rect 5910 51654 5962 51706
rect 5974 51654 6026 51706
rect 6038 51654 6090 51706
rect 6102 51654 6154 51706
rect 9110 51654 9162 51706
rect 9174 51654 9226 51706
rect 9238 51654 9290 51706
rect 9302 51654 9354 51706
rect 9366 51654 9418 51706
rect 2412 51552 2464 51604
rect 1124 51484 1176 51536
rect 572 51416 624 51468
rect 1768 51416 1820 51468
rect 2320 51416 2372 51468
rect 1124 51348 1176 51400
rect 2412 51348 2464 51400
rect 3056 51348 3108 51400
rect 9864 51391 9916 51400
rect 9864 51357 9873 51391
rect 9873 51357 9907 51391
rect 9907 51357 9916 51391
rect 9864 51348 9916 51357
rect 2964 51280 3016 51332
rect 1584 51255 1636 51264
rect 1584 51221 1593 51255
rect 1593 51221 1627 51255
rect 1627 51221 1636 51255
rect 1584 51212 1636 51221
rect 10048 51255 10100 51264
rect 10048 51221 10057 51255
rect 10057 51221 10091 51255
rect 10091 51221 10100 51255
rect 10048 51212 10100 51221
rect 4214 51110 4266 51162
rect 4278 51110 4330 51162
rect 4342 51110 4394 51162
rect 4406 51110 4458 51162
rect 4470 51110 4522 51162
rect 7478 51110 7530 51162
rect 7542 51110 7594 51162
rect 7606 51110 7658 51162
rect 7670 51110 7722 51162
rect 7734 51110 7786 51162
rect 1308 51008 1360 51060
rect 3424 51008 3476 51060
rect 3976 51008 4028 51060
rect 5172 51008 5224 51060
rect 6736 51008 6788 51060
rect 9864 51008 9916 51060
rect 1216 50940 1268 50992
rect 5264 50940 5316 50992
rect 1216 50804 1268 50856
rect 1308 50804 1360 50856
rect 3792 50872 3844 50924
rect 4068 50872 4120 50924
rect 10140 50915 10192 50924
rect 10140 50881 10149 50915
rect 10149 50881 10183 50915
rect 10183 50881 10192 50915
rect 10140 50872 10192 50881
rect 5632 50804 5684 50856
rect 1952 50736 2004 50788
rect 1308 50668 1360 50720
rect 2582 50566 2634 50618
rect 2646 50566 2698 50618
rect 2710 50566 2762 50618
rect 2774 50566 2826 50618
rect 2838 50566 2890 50618
rect 5846 50566 5898 50618
rect 5910 50566 5962 50618
rect 5974 50566 6026 50618
rect 6038 50566 6090 50618
rect 6102 50566 6154 50618
rect 9110 50566 9162 50618
rect 9174 50566 9226 50618
rect 9238 50566 9290 50618
rect 9302 50566 9354 50618
rect 9366 50566 9418 50618
rect 1308 50464 1360 50516
rect 204 50396 256 50448
rect 756 50328 808 50380
rect 204 50260 256 50312
rect 4712 50464 4764 50516
rect 6828 50464 6880 50516
rect 6552 50396 6604 50448
rect 1492 50260 1544 50312
rect 1952 50328 2004 50380
rect 4712 50328 4764 50380
rect 4988 50328 5040 50380
rect 1768 50303 1820 50312
rect 1768 50269 1777 50303
rect 1777 50269 1811 50303
rect 1811 50269 1820 50303
rect 1768 50260 1820 50269
rect 5540 50260 5592 50312
rect 9864 50303 9916 50312
rect 9864 50269 9873 50303
rect 9873 50269 9907 50303
rect 9907 50269 9916 50303
rect 9864 50260 9916 50269
rect 1952 50167 2004 50176
rect 1952 50133 1961 50167
rect 1961 50133 1995 50167
rect 1995 50133 2004 50167
rect 1952 50124 2004 50133
rect 2780 50124 2832 50176
rect 10048 50167 10100 50176
rect 10048 50133 10057 50167
rect 10057 50133 10091 50167
rect 10091 50133 10100 50167
rect 10048 50124 10100 50133
rect 940 49988 992 50040
rect 4214 50022 4266 50074
rect 4278 50022 4330 50074
rect 4342 50022 4394 50074
rect 4406 50022 4458 50074
rect 4470 50022 4522 50074
rect 7478 50022 7530 50074
rect 7542 50022 7594 50074
rect 7606 50022 7658 50074
rect 7670 50022 7722 50074
rect 7734 50022 7786 50074
rect 3240 49920 3292 49972
rect 9588 49920 9640 49972
rect 1676 49895 1728 49904
rect 1676 49861 1685 49895
rect 1685 49861 1719 49895
rect 1719 49861 1728 49895
rect 1676 49852 1728 49861
rect 1492 49784 1544 49836
rect 1768 49827 1820 49836
rect 1768 49793 1777 49827
rect 1777 49793 1811 49827
rect 1811 49793 1820 49827
rect 1768 49784 1820 49793
rect 4528 49852 4580 49904
rect 1952 49623 2004 49632
rect 1952 49589 1961 49623
rect 1961 49589 1995 49623
rect 1995 49589 2004 49623
rect 1952 49580 2004 49589
rect 2228 49580 2280 49632
rect 9680 49784 9732 49836
rect 3332 49648 3384 49700
rect 6276 49580 6328 49632
rect 2582 49478 2634 49530
rect 2646 49478 2698 49530
rect 2710 49478 2762 49530
rect 2774 49478 2826 49530
rect 2838 49478 2890 49530
rect 5846 49478 5898 49530
rect 5910 49478 5962 49530
rect 5974 49478 6026 49530
rect 6038 49478 6090 49530
rect 6102 49478 6154 49530
rect 9110 49478 9162 49530
rect 9174 49478 9226 49530
rect 9238 49478 9290 49530
rect 9302 49478 9354 49530
rect 9366 49478 9418 49530
rect 3332 49376 3384 49428
rect 3516 49376 3568 49428
rect 2504 49308 2556 49360
rect 3240 49308 3292 49360
rect 3884 49308 3936 49360
rect 5264 49240 5316 49292
rect 1492 49172 1544 49224
rect 1768 49215 1820 49224
rect 1768 49181 1777 49215
rect 1777 49181 1811 49215
rect 1811 49181 1820 49215
rect 1768 49172 1820 49181
rect 1676 49147 1728 49156
rect 1676 49113 1685 49147
rect 1685 49113 1719 49147
rect 1719 49113 1728 49147
rect 2780 49172 2832 49224
rect 3056 49172 3108 49224
rect 3976 49172 4028 49224
rect 9956 49172 10008 49224
rect 1676 49104 1728 49113
rect 2688 49104 2740 49156
rect 2872 49104 2924 49156
rect 6460 49104 6512 49156
rect 1400 49036 1452 49088
rect 3976 49079 4028 49088
rect 3976 49045 3985 49079
rect 3985 49045 4019 49079
rect 4019 49045 4028 49079
rect 3976 49036 4028 49045
rect 10048 49079 10100 49088
rect 10048 49045 10057 49079
rect 10057 49045 10091 49079
rect 10091 49045 10100 49079
rect 10048 49036 10100 49045
rect 4214 48934 4266 48986
rect 4278 48934 4330 48986
rect 4342 48934 4394 48986
rect 4406 48934 4458 48986
rect 4470 48934 4522 48986
rect 7478 48934 7530 48986
rect 7542 48934 7594 48986
rect 7606 48934 7658 48986
rect 7670 48934 7722 48986
rect 7734 48934 7786 48986
rect 3056 48832 3108 48884
rect 2872 48764 2924 48816
rect 3332 48764 3384 48816
rect 3608 48832 3660 48884
rect 1492 48696 1544 48748
rect 1308 48628 1360 48680
rect 1768 48739 1820 48748
rect 1768 48705 1777 48739
rect 1777 48705 1811 48739
rect 1811 48705 1820 48739
rect 1768 48696 1820 48705
rect 1676 48560 1728 48612
rect 3148 48696 3200 48748
rect 3424 48696 3476 48748
rect 3332 48628 3384 48680
rect 2320 48560 2372 48612
rect 3056 48560 3108 48612
rect 1308 48492 1360 48544
rect 1492 48492 1544 48544
rect 3332 48492 3384 48544
rect 3424 48492 3476 48544
rect 3792 48535 3844 48544
rect 3792 48501 3801 48535
rect 3801 48501 3835 48535
rect 3835 48501 3844 48535
rect 3792 48492 3844 48501
rect 9864 48832 9916 48884
rect 4068 48696 4120 48748
rect 4528 48560 4580 48612
rect 5540 48560 5592 48612
rect 8484 48492 8536 48544
rect 2582 48390 2634 48442
rect 2646 48390 2698 48442
rect 2710 48390 2762 48442
rect 2774 48390 2826 48442
rect 2838 48390 2890 48442
rect 5846 48390 5898 48442
rect 5910 48390 5962 48442
rect 5974 48390 6026 48442
rect 6038 48390 6090 48442
rect 6102 48390 6154 48442
rect 9110 48390 9162 48442
rect 9174 48390 9226 48442
rect 9238 48390 9290 48442
rect 9302 48390 9354 48442
rect 9366 48390 9418 48442
rect 2228 48288 2280 48340
rect 848 48220 900 48272
rect 2504 48220 2556 48272
rect 3700 48220 3752 48272
rect 4344 48220 4396 48272
rect 9680 48220 9732 48272
rect 756 48152 808 48204
rect 4528 48152 4580 48204
rect 7104 48152 7156 48204
rect 940 48084 992 48136
rect 2412 48127 2464 48136
rect 756 48016 808 48068
rect 2412 48093 2421 48127
rect 2421 48093 2455 48127
rect 2455 48093 2464 48127
rect 2412 48084 2464 48093
rect 5264 48084 5316 48136
rect 9496 48084 9548 48136
rect 7012 48016 7064 48068
rect 848 47948 900 48000
rect 1584 47991 1636 48000
rect 1584 47957 1593 47991
rect 1593 47957 1627 47991
rect 1627 47957 1636 47991
rect 1584 47948 1636 47957
rect 10048 47991 10100 48000
rect 10048 47957 10057 47991
rect 10057 47957 10091 47991
rect 10091 47957 10100 47991
rect 10048 47948 10100 47957
rect 4214 47846 4266 47898
rect 4278 47846 4330 47898
rect 4342 47846 4394 47898
rect 4406 47846 4458 47898
rect 4470 47846 4522 47898
rect 7478 47846 7530 47898
rect 7542 47846 7594 47898
rect 7606 47846 7658 47898
rect 7670 47846 7722 47898
rect 7734 47846 7786 47898
rect 1952 47676 2004 47728
rect 2320 47676 2372 47728
rect 1400 47651 1452 47660
rect 1400 47617 1409 47651
rect 1409 47617 1443 47651
rect 1443 47617 1452 47651
rect 1400 47608 1452 47617
rect 3792 47608 3844 47660
rect 8300 47608 8352 47660
rect 1952 47540 2004 47592
rect 1584 47447 1636 47456
rect 1584 47413 1593 47447
rect 1593 47413 1627 47447
rect 1627 47413 1636 47447
rect 1584 47404 1636 47413
rect 3792 47404 3844 47456
rect 3976 47404 4028 47456
rect 10048 47447 10100 47456
rect 10048 47413 10057 47447
rect 10057 47413 10091 47447
rect 10091 47413 10100 47447
rect 10048 47404 10100 47413
rect 2582 47302 2634 47354
rect 2646 47302 2698 47354
rect 2710 47302 2762 47354
rect 2774 47302 2826 47354
rect 2838 47302 2890 47354
rect 5846 47302 5898 47354
rect 5910 47302 5962 47354
rect 5974 47302 6026 47354
rect 6038 47302 6090 47354
rect 6102 47302 6154 47354
rect 9110 47302 9162 47354
rect 9174 47302 9226 47354
rect 9238 47302 9290 47354
rect 9302 47302 9354 47354
rect 9366 47302 9418 47354
rect 1584 47200 1636 47252
rect 1768 47200 1820 47252
rect 1952 47243 2004 47252
rect 1952 47209 1961 47243
rect 1961 47209 1995 47243
rect 1995 47209 2004 47243
rect 1952 47200 2004 47209
rect 2412 47200 2464 47252
rect 9496 47200 9548 47252
rect 9956 47243 10008 47252
rect 9956 47209 9965 47243
rect 9965 47209 9999 47243
rect 9999 47209 10008 47243
rect 9956 47200 10008 47209
rect 3976 47175 4028 47184
rect 3976 47141 3985 47175
rect 3985 47141 4019 47175
rect 4019 47141 4028 47175
rect 3976 47132 4028 47141
rect 4436 47132 4488 47184
rect 6460 47132 6512 47184
rect 2504 47039 2556 47048
rect 2504 47005 2513 47039
rect 2513 47005 2547 47039
rect 2547 47005 2556 47039
rect 2504 46996 2556 47005
rect 2688 47064 2740 47116
rect 2964 46996 3016 47048
rect 4436 46996 4488 47048
rect 6552 47064 6604 47116
rect 4252 46928 4304 46980
rect 20 46724 72 46776
rect 4214 46758 4266 46810
rect 4278 46758 4330 46810
rect 4342 46758 4394 46810
rect 4406 46758 4458 46810
rect 4470 46758 4522 46810
rect 7478 46758 7530 46810
rect 7542 46758 7594 46810
rect 7606 46758 7658 46810
rect 7670 46758 7722 46810
rect 7734 46758 7786 46810
rect 756 46656 808 46708
rect 3056 46656 3108 46708
rect 3424 46656 3476 46708
rect 8300 46656 8352 46708
rect 3424 46520 3476 46572
rect 6552 46563 6604 46572
rect 6552 46529 6561 46563
rect 6561 46529 6595 46563
rect 6595 46529 6604 46563
rect 6552 46520 6604 46529
rect 8116 46520 8168 46572
rect 664 46452 716 46504
rect 1952 46495 2004 46504
rect 1952 46461 1961 46495
rect 1961 46461 1995 46495
rect 1995 46461 2004 46495
rect 1952 46452 2004 46461
rect 4068 46452 4120 46504
rect 10048 46427 10100 46436
rect 10048 46393 10057 46427
rect 10057 46393 10091 46427
rect 10091 46393 10100 46427
rect 10048 46384 10100 46393
rect 20 46316 72 46368
rect 1032 46316 1084 46368
rect 2504 46316 2556 46368
rect 4528 46316 4580 46368
rect 4712 46316 4764 46368
rect 2582 46214 2634 46266
rect 2646 46214 2698 46266
rect 2710 46214 2762 46266
rect 2774 46214 2826 46266
rect 2838 46214 2890 46266
rect 5846 46214 5898 46266
rect 5910 46214 5962 46266
rect 5974 46214 6026 46266
rect 6038 46214 6090 46266
rect 6102 46214 6154 46266
rect 9110 46214 9162 46266
rect 9174 46214 9226 46266
rect 9238 46214 9290 46266
rect 9302 46214 9354 46266
rect 9366 46214 9418 46266
rect 112 46112 164 46164
rect 1032 46112 1084 46164
rect 1952 46112 2004 46164
rect 4712 46112 4764 46164
rect 4896 46112 4948 46164
rect 3332 46044 3384 46096
rect 3516 46044 3568 46096
rect 1492 45976 1544 46028
rect 1952 45976 2004 46028
rect 2964 45976 3016 46028
rect 2872 45951 2924 45960
rect 2872 45917 2881 45951
rect 2881 45917 2915 45951
rect 2915 45917 2924 45951
rect 2872 45908 2924 45917
rect 3056 45908 3108 45960
rect 3332 45908 3384 45960
rect 6920 45908 6972 45960
rect 4068 45840 4120 45892
rect 4528 45840 4580 45892
rect 4988 45840 5040 45892
rect 1584 45772 1636 45824
rect 3056 45815 3108 45824
rect 3056 45781 3065 45815
rect 3065 45781 3099 45815
rect 3099 45781 3108 45815
rect 3056 45772 3108 45781
rect 10048 45815 10100 45824
rect 10048 45781 10057 45815
rect 10057 45781 10091 45815
rect 10091 45781 10100 45815
rect 10048 45772 10100 45781
rect 4214 45670 4266 45722
rect 4278 45670 4330 45722
rect 4342 45670 4394 45722
rect 4406 45670 4458 45722
rect 4470 45670 4522 45722
rect 7478 45670 7530 45722
rect 7542 45670 7594 45722
rect 7606 45670 7658 45722
rect 7670 45670 7722 45722
rect 7734 45670 7786 45722
rect 2320 45611 2372 45620
rect 2320 45577 2329 45611
rect 2329 45577 2363 45611
rect 2363 45577 2372 45611
rect 2320 45568 2372 45577
rect 3792 45500 3844 45552
rect 5540 45500 5592 45552
rect 1308 45432 1360 45484
rect 2872 45475 2924 45484
rect 2872 45441 2881 45475
rect 2881 45441 2915 45475
rect 2915 45441 2924 45475
rect 2872 45432 2924 45441
rect 5356 45432 5408 45484
rect 4160 45364 4212 45416
rect 2596 45296 2648 45348
rect 6920 45296 6972 45348
rect 1584 45271 1636 45280
rect 1584 45237 1593 45271
rect 1593 45237 1627 45271
rect 1627 45237 1636 45271
rect 1584 45228 1636 45237
rect 2582 45126 2634 45178
rect 2646 45126 2698 45178
rect 2710 45126 2762 45178
rect 2774 45126 2826 45178
rect 2838 45126 2890 45178
rect 5846 45126 5898 45178
rect 5910 45126 5962 45178
rect 5974 45126 6026 45178
rect 6038 45126 6090 45178
rect 6102 45126 6154 45178
rect 9110 45126 9162 45178
rect 9174 45126 9226 45178
rect 9238 45126 9290 45178
rect 9302 45126 9354 45178
rect 9366 45126 9418 45178
rect 5356 45067 5408 45076
rect 5356 45033 5365 45067
rect 5365 45033 5399 45067
rect 5399 45033 5408 45067
rect 5356 45024 5408 45033
rect 8116 45024 8168 45076
rect 1492 44956 1544 45008
rect 1492 44863 1544 44872
rect 1492 44829 1501 44863
rect 1501 44829 1535 44863
rect 1535 44829 1544 44863
rect 1492 44820 1544 44829
rect 2320 44888 2372 44940
rect 8576 44888 8628 44940
rect 1584 44684 1636 44736
rect 2964 44727 3016 44736
rect 2964 44693 2973 44727
rect 2973 44693 3007 44727
rect 3007 44693 3016 44727
rect 2964 44684 3016 44693
rect 5540 44820 5592 44872
rect 9864 44863 9916 44872
rect 9864 44829 9873 44863
rect 9873 44829 9907 44863
rect 9907 44829 9916 44863
rect 9864 44820 9916 44829
rect 6552 44752 6604 44804
rect 5632 44684 5684 44736
rect 6184 44684 6236 44736
rect 6644 44684 6696 44736
rect 10048 44727 10100 44736
rect 10048 44693 10057 44727
rect 10057 44693 10091 44727
rect 10091 44693 10100 44727
rect 10048 44684 10100 44693
rect 4214 44582 4266 44634
rect 4278 44582 4330 44634
rect 4342 44582 4394 44634
rect 4406 44582 4458 44634
rect 4470 44582 4522 44634
rect 7478 44582 7530 44634
rect 7542 44582 7594 44634
rect 7606 44582 7658 44634
rect 7670 44582 7722 44634
rect 7734 44582 7786 44634
rect 2964 44480 3016 44532
rect 3332 44480 3384 44532
rect 9864 44480 9916 44532
rect 848 44344 900 44396
rect 3792 44344 3844 44396
rect 6552 44387 6604 44396
rect 6552 44353 6561 44387
rect 6561 44353 6595 44387
rect 6595 44353 6604 44387
rect 6552 44344 6604 44353
rect 9864 44387 9916 44396
rect 9864 44353 9873 44387
rect 9873 44353 9907 44387
rect 9907 44353 9916 44387
rect 9864 44344 9916 44353
rect 3332 44276 3384 44328
rect 3148 44183 3200 44192
rect 3148 44149 3157 44183
rect 3157 44149 3191 44183
rect 3191 44149 3200 44183
rect 3148 44140 3200 44149
rect 10048 44183 10100 44192
rect 10048 44149 10057 44183
rect 10057 44149 10091 44183
rect 10091 44149 10100 44183
rect 10048 44140 10100 44149
rect 2582 44038 2634 44090
rect 2646 44038 2698 44090
rect 2710 44038 2762 44090
rect 2774 44038 2826 44090
rect 2838 44038 2890 44090
rect 5846 44038 5898 44090
rect 5910 44038 5962 44090
rect 5974 44038 6026 44090
rect 6038 44038 6090 44090
rect 6102 44038 6154 44090
rect 9110 44038 9162 44090
rect 9174 44038 9226 44090
rect 9238 44038 9290 44090
rect 9302 44038 9354 44090
rect 9366 44038 9418 44090
rect 1492 43936 1544 43988
rect 3332 43936 3384 43988
rect 3792 43936 3844 43988
rect 3976 43936 4028 43988
rect 6552 43936 6604 43988
rect 5632 43868 5684 43920
rect 848 43664 900 43716
rect 2596 43732 2648 43784
rect 3056 43732 3108 43784
rect 3148 43732 3200 43784
rect 3332 43732 3384 43784
rect 6644 43732 6696 43784
rect 9956 43732 10008 43784
rect 5540 43664 5592 43716
rect 3976 43639 4028 43648
rect 3976 43605 3985 43639
rect 3985 43605 4019 43639
rect 4019 43605 4028 43639
rect 3976 43596 4028 43605
rect 10048 43639 10100 43648
rect 10048 43605 10057 43639
rect 10057 43605 10091 43639
rect 10091 43605 10100 43639
rect 10048 43596 10100 43605
rect 4214 43494 4266 43546
rect 4278 43494 4330 43546
rect 4342 43494 4394 43546
rect 4406 43494 4458 43546
rect 4470 43494 4522 43546
rect 7478 43494 7530 43546
rect 7542 43494 7594 43546
rect 7606 43494 7658 43546
rect 7670 43494 7722 43546
rect 7734 43494 7786 43546
rect 940 43392 992 43444
rect 3148 43392 3200 43444
rect 3332 43435 3384 43444
rect 3332 43401 3341 43435
rect 3341 43401 3375 43435
rect 3375 43401 3384 43435
rect 3332 43392 3384 43401
rect 6368 43392 6420 43444
rect 6920 43392 6972 43444
rect 9956 43435 10008 43444
rect 9956 43401 9965 43435
rect 9965 43401 9999 43435
rect 9999 43401 10008 43435
rect 9956 43392 10008 43401
rect 1768 43324 1820 43376
rect 1492 43231 1544 43240
rect 1492 43197 1501 43231
rect 1501 43197 1535 43231
rect 1535 43197 1544 43231
rect 1492 43188 1544 43197
rect 2964 43299 3016 43308
rect 2964 43265 2973 43299
rect 2973 43265 3007 43299
rect 3007 43265 3016 43299
rect 2964 43256 3016 43265
rect 3148 43299 3200 43308
rect 3148 43265 3157 43299
rect 3157 43265 3191 43299
rect 3191 43265 3200 43299
rect 3148 43256 3200 43265
rect 3332 43256 3384 43308
rect 3700 43256 3752 43308
rect 9680 43256 9732 43308
rect 9772 43188 9824 43240
rect 848 43120 900 43172
rect 2596 43120 2648 43172
rect 3608 43120 3660 43172
rect 3976 43163 4028 43172
rect 3976 43129 3985 43163
rect 3985 43129 4019 43163
rect 4019 43129 4028 43163
rect 3976 43120 4028 43129
rect 3792 43052 3844 43104
rect 2582 42950 2634 43002
rect 2646 42950 2698 43002
rect 2710 42950 2762 43002
rect 2774 42950 2826 43002
rect 2838 42950 2890 43002
rect 5846 42950 5898 43002
rect 5910 42950 5962 43002
rect 5974 42950 6026 43002
rect 6038 42950 6090 43002
rect 6102 42950 6154 43002
rect 9110 42950 9162 43002
rect 9174 42950 9226 43002
rect 9238 42950 9290 43002
rect 9302 42950 9354 43002
rect 9366 42950 9418 43002
rect 1492 42848 1544 42900
rect 3332 42848 3384 42900
rect 6276 42712 6328 42764
rect 8392 42712 8444 42764
rect 848 42644 900 42696
rect 1676 42576 1728 42628
rect 3148 42644 3200 42696
rect 3516 42644 3568 42696
rect 4160 42644 4212 42696
rect 6460 42687 6512 42696
rect 6460 42653 6469 42687
rect 6469 42653 6503 42687
rect 6503 42653 6512 42687
rect 6460 42644 6512 42653
rect 9956 42644 10008 42696
rect 2780 42551 2832 42560
rect 2780 42517 2789 42551
rect 2789 42517 2823 42551
rect 2823 42517 2832 42551
rect 3976 42551 4028 42560
rect 2780 42508 2832 42517
rect 3976 42517 3985 42551
rect 3985 42517 4019 42551
rect 4019 42517 4028 42551
rect 3976 42508 4028 42517
rect 9864 42508 9916 42560
rect 10048 42551 10100 42560
rect 10048 42517 10057 42551
rect 10057 42517 10091 42551
rect 10091 42517 10100 42551
rect 10048 42508 10100 42517
rect 4214 42406 4266 42458
rect 4278 42406 4330 42458
rect 4342 42406 4394 42458
rect 4406 42406 4458 42458
rect 4470 42406 4522 42458
rect 7478 42406 7530 42458
rect 7542 42406 7594 42458
rect 7606 42406 7658 42458
rect 7670 42406 7722 42458
rect 7734 42406 7786 42458
rect 3332 42304 3384 42356
rect 3976 42304 4028 42356
rect 4436 42236 4488 42288
rect 4804 42236 4856 42288
rect 1768 42168 1820 42220
rect 2136 42211 2188 42220
rect 2136 42177 2145 42211
rect 2145 42177 2179 42211
rect 2179 42177 2188 42211
rect 2136 42168 2188 42177
rect 2872 42211 2924 42220
rect 2872 42177 2881 42211
rect 2881 42177 2915 42211
rect 2915 42177 2924 42211
rect 2872 42168 2924 42177
rect 9496 42168 9548 42220
rect 2320 42100 2372 42152
rect 2136 42032 2188 42084
rect 1584 42007 1636 42016
rect 1584 41973 1593 42007
rect 1593 41973 1627 42007
rect 1627 41973 1636 42007
rect 1584 41964 1636 41973
rect 2320 42007 2372 42016
rect 2320 41973 2329 42007
rect 2329 41973 2363 42007
rect 2363 41973 2372 42007
rect 2320 41964 2372 41973
rect 3056 42007 3108 42016
rect 3056 41973 3065 42007
rect 3065 41973 3099 42007
rect 3099 41973 3108 42007
rect 3056 41964 3108 41973
rect 10048 42007 10100 42016
rect 10048 41973 10057 42007
rect 10057 41973 10091 42007
rect 10091 41973 10100 42007
rect 10048 41964 10100 41973
rect 2582 41862 2634 41914
rect 2646 41862 2698 41914
rect 2710 41862 2762 41914
rect 2774 41862 2826 41914
rect 2838 41862 2890 41914
rect 5846 41862 5898 41914
rect 5910 41862 5962 41914
rect 5974 41862 6026 41914
rect 6038 41862 6090 41914
rect 6102 41862 6154 41914
rect 9110 41862 9162 41914
rect 9174 41862 9226 41914
rect 9238 41862 9290 41914
rect 9302 41862 9354 41914
rect 9366 41862 9418 41914
rect 664 41760 716 41812
rect 9680 41760 9732 41812
rect 9956 41803 10008 41812
rect 9956 41769 9965 41803
rect 9965 41769 9999 41803
rect 9999 41769 10008 41803
rect 9956 41760 10008 41769
rect 6368 41692 6420 41744
rect 664 41624 716 41676
rect 1400 41624 1452 41676
rect 2320 41624 2372 41676
rect 2872 41624 2924 41676
rect 848 41488 900 41540
rect 1400 41488 1452 41540
rect 1768 41531 1820 41540
rect 1768 41497 1777 41531
rect 1777 41497 1811 41531
rect 1811 41497 1820 41531
rect 1768 41488 1820 41497
rect 2688 41556 2740 41608
rect 3700 41624 3752 41676
rect 5264 41624 5316 41676
rect 3056 41556 3108 41608
rect 5448 41556 5500 41608
rect 5908 41556 5960 41608
rect 6368 41556 6420 41608
rect 9772 41556 9824 41608
rect 5816 41488 5868 41540
rect 6644 41488 6696 41540
rect 2320 41420 2372 41472
rect 5080 41420 5132 41472
rect 7012 41420 7064 41472
rect 4214 41318 4266 41370
rect 4278 41318 4330 41370
rect 4342 41318 4394 41370
rect 4406 41318 4458 41370
rect 4470 41318 4522 41370
rect 7478 41318 7530 41370
rect 7542 41318 7594 41370
rect 7606 41318 7658 41370
rect 7670 41318 7722 41370
rect 7734 41318 7786 41370
rect 756 41216 808 41268
rect 1492 41216 1544 41268
rect 1768 41216 1820 41268
rect 2688 41216 2740 41268
rect 2872 41259 2924 41268
rect 2872 41225 2881 41259
rect 2881 41225 2915 41259
rect 2915 41225 2924 41259
rect 2872 41216 2924 41225
rect 6460 41216 6512 41268
rect 3516 41148 3568 41200
rect 5540 41148 5592 41200
rect 6920 41148 6972 41200
rect 1400 41080 1452 41132
rect 2780 41080 2832 41132
rect 3056 41012 3108 41064
rect 4436 41012 4488 41064
rect 5632 41080 5684 41132
rect 5908 41080 5960 41132
rect 7012 41080 7064 41132
rect 5816 41012 5868 41064
rect 6460 41012 6512 41064
rect 2780 40944 2832 40996
rect 10048 40987 10100 40996
rect 10048 40953 10057 40987
rect 10057 40953 10091 40987
rect 10091 40953 10100 40987
rect 10048 40944 10100 40953
rect 3056 40876 3108 40928
rect 4988 40876 5040 40928
rect 5448 40876 5500 40928
rect 2582 40774 2634 40826
rect 2646 40774 2698 40826
rect 2710 40774 2762 40826
rect 2774 40774 2826 40826
rect 2838 40774 2890 40826
rect 5846 40774 5898 40826
rect 5910 40774 5962 40826
rect 5974 40774 6026 40826
rect 6038 40774 6090 40826
rect 6102 40774 6154 40826
rect 9110 40774 9162 40826
rect 9174 40774 9226 40826
rect 9238 40774 9290 40826
rect 9302 40774 9354 40826
rect 9366 40774 9418 40826
rect 1032 40672 1084 40724
rect 2136 40604 2188 40656
rect 9496 40672 9548 40724
rect 2872 40604 2924 40656
rect 4436 40604 4488 40656
rect 4988 40604 5040 40656
rect 5356 40604 5408 40656
rect 3884 40536 3936 40588
rect 2136 40511 2188 40520
rect 2136 40477 2145 40511
rect 2145 40477 2179 40511
rect 2179 40477 2188 40511
rect 2136 40468 2188 40477
rect 5356 40468 5408 40520
rect 9864 40511 9916 40520
rect 9864 40477 9873 40511
rect 9873 40477 9907 40511
rect 9907 40477 9916 40511
rect 9864 40468 9916 40477
rect 112 40400 164 40452
rect 1768 40400 1820 40452
rect 1584 40375 1636 40384
rect 1584 40341 1593 40375
rect 1593 40341 1627 40375
rect 1627 40341 1636 40375
rect 1584 40332 1636 40341
rect 3976 40375 4028 40384
rect 3976 40341 3985 40375
rect 3985 40341 4019 40375
rect 4019 40341 4028 40375
rect 3976 40332 4028 40341
rect 10048 40375 10100 40384
rect 10048 40341 10057 40375
rect 10057 40341 10091 40375
rect 10091 40341 10100 40375
rect 10048 40332 10100 40341
rect 4214 40230 4266 40282
rect 4278 40230 4330 40282
rect 4342 40230 4394 40282
rect 4406 40230 4458 40282
rect 4470 40230 4522 40282
rect 7478 40230 7530 40282
rect 7542 40230 7594 40282
rect 7606 40230 7658 40282
rect 7670 40230 7722 40282
rect 7734 40230 7786 40282
rect 2136 40128 2188 40180
rect 9864 40128 9916 40180
rect 664 40060 716 40112
rect 2964 40060 3016 40112
rect 5448 40060 5500 40112
rect 6920 40060 6972 40112
rect 1032 39992 1084 40044
rect 1400 39992 1452 40044
rect 2412 39992 2464 40044
rect 2504 39992 2556 40044
rect 2780 39992 2832 40044
rect 9864 40035 9916 40044
rect 9864 40001 9873 40035
rect 9873 40001 9907 40035
rect 9907 40001 9916 40035
rect 9864 39992 9916 40001
rect 5448 39924 5500 39976
rect 5632 39924 5684 39976
rect 2872 39856 2924 39908
rect 3976 39831 4028 39840
rect 3976 39797 3985 39831
rect 3985 39797 4019 39831
rect 4019 39797 4028 39831
rect 3976 39788 4028 39797
rect 10048 39831 10100 39840
rect 10048 39797 10057 39831
rect 10057 39797 10091 39831
rect 10091 39797 10100 39831
rect 10048 39788 10100 39797
rect 2582 39686 2634 39738
rect 2646 39686 2698 39738
rect 2710 39686 2762 39738
rect 2774 39686 2826 39738
rect 2838 39686 2890 39738
rect 5846 39686 5898 39738
rect 5910 39686 5962 39738
rect 5974 39686 6026 39738
rect 6038 39686 6090 39738
rect 6102 39686 6154 39738
rect 9110 39686 9162 39738
rect 9174 39686 9226 39738
rect 9238 39686 9290 39738
rect 9302 39686 9354 39738
rect 9366 39686 9418 39738
rect 6920 39584 6972 39636
rect 9864 39627 9916 39636
rect 9864 39593 9873 39627
rect 9873 39593 9907 39627
rect 9907 39593 9916 39627
rect 9864 39584 9916 39593
rect 6368 39516 6420 39568
rect 7012 39516 7064 39568
rect 3056 39448 3108 39500
rect 112 39380 164 39432
rect 2504 39380 2556 39432
rect 2872 39423 2924 39432
rect 2872 39389 2881 39423
rect 2881 39389 2915 39423
rect 2915 39389 2924 39423
rect 2872 39380 2924 39389
rect 2780 39312 2832 39364
rect 4068 39380 4120 39432
rect 3056 39312 3108 39364
rect 5632 39380 5684 39432
rect 6736 39380 6788 39432
rect 8760 39380 8812 39432
rect 1400 39244 1452 39296
rect 3976 39287 4028 39296
rect 3976 39253 3985 39287
rect 3985 39253 4019 39287
rect 4019 39253 4028 39287
rect 3976 39244 4028 39253
rect 4214 39142 4266 39194
rect 4278 39142 4330 39194
rect 4342 39142 4394 39194
rect 4406 39142 4458 39194
rect 4470 39142 4522 39194
rect 7478 39142 7530 39194
rect 7542 39142 7594 39194
rect 7606 39142 7658 39194
rect 7670 39142 7722 39194
rect 7734 39142 7786 39194
rect 1032 39040 1084 39092
rect 2412 39040 2464 39092
rect 6736 39083 6788 39092
rect 6736 39049 6745 39083
rect 6745 39049 6779 39083
rect 6779 39049 6788 39083
rect 6736 39040 6788 39049
rect 480 38904 532 38956
rect 3700 38972 3752 39024
rect 4436 38972 4488 39024
rect 5632 38972 5684 39024
rect 4712 38904 4764 38956
rect 6460 38904 6512 38956
rect 8208 38904 8260 38956
rect 4344 38836 4396 38888
rect 2780 38768 2832 38820
rect 4252 38768 4304 38820
rect 4528 38768 4580 38820
rect 4712 38768 4764 38820
rect 2964 38743 3016 38752
rect 2964 38709 2973 38743
rect 2973 38709 3007 38743
rect 3007 38709 3016 38743
rect 2964 38700 3016 38709
rect 3700 38743 3752 38752
rect 3700 38709 3709 38743
rect 3709 38709 3743 38743
rect 3743 38709 3752 38743
rect 3700 38700 3752 38709
rect 4620 38700 4672 38752
rect 7104 38700 7156 38752
rect 10048 38743 10100 38752
rect 10048 38709 10057 38743
rect 10057 38709 10091 38743
rect 10091 38709 10100 38743
rect 10048 38700 10100 38709
rect 2582 38598 2634 38650
rect 2646 38598 2698 38650
rect 2710 38598 2762 38650
rect 2774 38598 2826 38650
rect 2838 38598 2890 38650
rect 5846 38598 5898 38650
rect 5910 38598 5962 38650
rect 5974 38598 6026 38650
rect 6038 38598 6090 38650
rect 6102 38598 6154 38650
rect 9110 38598 9162 38650
rect 9174 38598 9226 38650
rect 9238 38598 9290 38650
rect 9302 38598 9354 38650
rect 9366 38598 9418 38650
rect 1492 38496 1544 38548
rect 2412 38496 2464 38548
rect 5356 38496 5408 38548
rect 388 38360 440 38412
rect 4436 38360 4488 38412
rect 3700 38292 3752 38344
rect 4252 38292 4304 38344
rect 2688 38224 2740 38276
rect 3516 38224 3568 38276
rect 5356 38292 5408 38344
rect 8484 38292 8536 38344
rect 5724 38224 5776 38276
rect 10048 38199 10100 38208
rect 10048 38165 10057 38199
rect 10057 38165 10091 38199
rect 10091 38165 10100 38199
rect 10048 38156 10100 38165
rect 4214 38054 4266 38106
rect 4278 38054 4330 38106
rect 4342 38054 4394 38106
rect 4406 38054 4458 38106
rect 4470 38054 4522 38106
rect 7478 38054 7530 38106
rect 7542 38054 7594 38106
rect 7606 38054 7658 38106
rect 7670 38054 7722 38106
rect 7734 38054 7786 38106
rect 1492 37952 1544 38004
rect 2688 37995 2740 38004
rect 2688 37961 2697 37995
rect 2697 37961 2731 37995
rect 2731 37961 2740 37995
rect 2688 37952 2740 37961
rect 9772 37952 9824 38004
rect 1032 37884 1084 37936
rect 2780 37884 2832 37936
rect 3424 37927 3476 37936
rect 3424 37893 3433 37927
rect 3433 37893 3467 37927
rect 3467 37893 3476 37927
rect 3424 37884 3476 37893
rect 1032 37748 1084 37800
rect 2596 37816 2648 37868
rect 2964 37816 3016 37868
rect 5356 37816 5408 37868
rect 1584 37612 1636 37664
rect 2582 37510 2634 37562
rect 2646 37510 2698 37562
rect 2710 37510 2762 37562
rect 2774 37510 2826 37562
rect 2838 37510 2890 37562
rect 5846 37510 5898 37562
rect 5910 37510 5962 37562
rect 5974 37510 6026 37562
rect 6038 37510 6090 37562
rect 6102 37510 6154 37562
rect 9110 37510 9162 37562
rect 9174 37510 9226 37562
rect 9238 37510 9290 37562
rect 9302 37510 9354 37562
rect 9366 37510 9418 37562
rect 2412 37340 2464 37392
rect 5724 37272 5776 37324
rect 2596 37204 2648 37256
rect 2964 37204 3016 37256
rect 3792 37247 3844 37256
rect 3792 37213 3801 37247
rect 3801 37213 3835 37247
rect 3835 37213 3844 37247
rect 3792 37204 3844 37213
rect 8576 37204 8628 37256
rect 2412 37136 2464 37188
rect 6368 37136 6420 37188
rect 2688 37068 2740 37120
rect 3976 37111 4028 37120
rect 3976 37077 3985 37111
rect 3985 37077 4019 37111
rect 4019 37077 4028 37111
rect 3976 37068 4028 37077
rect 8208 37111 8260 37120
rect 8208 37077 8217 37111
rect 8217 37077 8251 37111
rect 8251 37077 8260 37111
rect 8208 37068 8260 37077
rect 10048 37111 10100 37120
rect 10048 37077 10057 37111
rect 10057 37077 10091 37111
rect 10091 37077 10100 37111
rect 10048 37068 10100 37077
rect 4214 36966 4266 37018
rect 4278 36966 4330 37018
rect 4342 36966 4394 37018
rect 4406 36966 4458 37018
rect 4470 36966 4522 37018
rect 7478 36966 7530 37018
rect 7542 36966 7594 37018
rect 7606 36966 7658 37018
rect 7670 36966 7722 37018
rect 7734 36966 7786 37018
rect 2412 36907 2464 36916
rect 2412 36873 2421 36907
rect 2421 36873 2455 36907
rect 2455 36873 2464 36907
rect 2412 36864 2464 36873
rect 3792 36864 3844 36916
rect 6368 36907 6420 36916
rect 6368 36873 6377 36907
rect 6377 36873 6411 36907
rect 6411 36873 6420 36907
rect 6368 36864 6420 36873
rect 8484 36864 8536 36916
rect 2596 36728 2648 36780
rect 6828 36796 6880 36848
rect 3148 36728 3200 36780
rect 3516 36728 3568 36780
rect 6552 36771 6604 36780
rect 6552 36737 6561 36771
rect 6561 36737 6595 36771
rect 6595 36737 6604 36771
rect 6552 36728 6604 36737
rect 7196 36771 7248 36780
rect 7196 36737 7205 36771
rect 7205 36737 7239 36771
rect 7239 36737 7248 36771
rect 7196 36728 7248 36737
rect 9864 36771 9916 36780
rect 9864 36737 9873 36771
rect 9873 36737 9907 36771
rect 9907 36737 9916 36771
rect 9864 36728 9916 36737
rect 1584 36660 1636 36712
rect 2412 36660 2464 36712
rect 940 36592 992 36644
rect 4068 36592 4120 36644
rect 4620 36592 4672 36644
rect 5448 36592 5500 36644
rect 5080 36524 5132 36576
rect 5356 36524 5408 36576
rect 5540 36524 5592 36576
rect 6460 36524 6512 36576
rect 10048 36567 10100 36576
rect 10048 36533 10057 36567
rect 10057 36533 10091 36567
rect 10091 36533 10100 36567
rect 10048 36524 10100 36533
rect 2582 36422 2634 36474
rect 2646 36422 2698 36474
rect 2710 36422 2762 36474
rect 2774 36422 2826 36474
rect 2838 36422 2890 36474
rect 5846 36422 5898 36474
rect 5910 36422 5962 36474
rect 5974 36422 6026 36474
rect 6038 36422 6090 36474
rect 6102 36422 6154 36474
rect 9110 36422 9162 36474
rect 9174 36422 9226 36474
rect 9238 36422 9290 36474
rect 9302 36422 9354 36474
rect 9366 36422 9418 36474
rect 1952 36363 2004 36372
rect 1952 36329 1961 36363
rect 1961 36329 1995 36363
rect 1995 36329 2004 36363
rect 1952 36320 2004 36329
rect 3976 36363 4028 36372
rect 3976 36329 3985 36363
rect 3985 36329 4019 36363
rect 4019 36329 4028 36363
rect 3976 36320 4028 36329
rect 9864 36320 9916 36372
rect 6644 36252 6696 36304
rect 6276 36184 6328 36236
rect 4712 36159 4764 36168
rect 4712 36125 4721 36159
rect 4721 36125 4755 36159
rect 4755 36125 4764 36159
rect 4712 36116 4764 36125
rect 9864 36159 9916 36168
rect 9864 36125 9873 36159
rect 9873 36125 9907 36159
rect 9907 36125 9916 36159
rect 9864 36116 9916 36125
rect 1952 36048 2004 36100
rect 2780 35980 2832 36032
rect 10048 36023 10100 36032
rect 10048 35989 10057 36023
rect 10057 35989 10091 36023
rect 10091 35989 10100 36023
rect 10048 35980 10100 35989
rect 4214 35878 4266 35930
rect 4278 35878 4330 35930
rect 4342 35878 4394 35930
rect 4406 35878 4458 35930
rect 4470 35878 4522 35930
rect 7478 35878 7530 35930
rect 7542 35878 7594 35930
rect 7606 35878 7658 35930
rect 7670 35878 7722 35930
rect 7734 35878 7786 35930
rect 4712 35776 4764 35828
rect 6552 35776 6604 35828
rect 7196 35776 7248 35828
rect 2136 35640 2188 35692
rect 2964 35640 3016 35692
rect 3976 35683 4028 35692
rect 3976 35649 3985 35683
rect 3985 35649 4019 35683
rect 4019 35649 4028 35683
rect 3976 35640 4028 35649
rect 5540 35640 5592 35692
rect 6276 35640 6328 35692
rect 4620 35572 4672 35624
rect 6368 35615 6420 35624
rect 6368 35581 6377 35615
rect 6377 35581 6411 35615
rect 6411 35581 6420 35615
rect 6368 35572 6420 35581
rect 1400 35504 1452 35556
rect 2136 35504 2188 35556
rect 2412 35504 2464 35556
rect 1584 35479 1636 35488
rect 1584 35445 1593 35479
rect 1593 35445 1627 35479
rect 1627 35445 1636 35479
rect 1584 35436 1636 35445
rect 2582 35334 2634 35386
rect 2646 35334 2698 35386
rect 2710 35334 2762 35386
rect 2774 35334 2826 35386
rect 2838 35334 2890 35386
rect 5846 35334 5898 35386
rect 5910 35334 5962 35386
rect 5974 35334 6026 35386
rect 6038 35334 6090 35386
rect 6102 35334 6154 35386
rect 9110 35334 9162 35386
rect 9174 35334 9226 35386
rect 9238 35334 9290 35386
rect 9302 35334 9354 35386
rect 9366 35334 9418 35386
rect 9864 35232 9916 35284
rect 1492 35164 1544 35216
rect 2596 35164 2648 35216
rect 1676 35028 1728 35080
rect 2044 35028 2096 35080
rect 3148 35028 3200 35080
rect 4068 35028 4120 35080
rect 1584 34935 1636 34944
rect 1584 34901 1593 34935
rect 1593 34901 1627 34935
rect 1627 34901 1636 34935
rect 1584 34892 1636 34901
rect 2320 34935 2372 34944
rect 2320 34901 2329 34935
rect 2329 34901 2363 34935
rect 2363 34901 2372 34935
rect 2320 34892 2372 34901
rect 10048 34935 10100 34944
rect 10048 34901 10057 34935
rect 10057 34901 10091 34935
rect 10091 34901 10100 34935
rect 10048 34892 10100 34901
rect 4214 34790 4266 34842
rect 4278 34790 4330 34842
rect 4342 34790 4394 34842
rect 4406 34790 4458 34842
rect 4470 34790 4522 34842
rect 7478 34790 7530 34842
rect 7542 34790 7594 34842
rect 7606 34790 7658 34842
rect 7670 34790 7722 34842
rect 7734 34790 7786 34842
rect 1492 34688 1544 34740
rect 4068 34688 4120 34740
rect 9588 34688 9640 34740
rect 572 34552 624 34604
rect 1860 34552 1912 34604
rect 2596 34552 2648 34604
rect 2228 34484 2280 34536
rect 5540 34552 5592 34604
rect 572 34416 624 34468
rect 1860 34416 1912 34468
rect 2136 34416 2188 34468
rect 3976 34416 4028 34468
rect 2228 34348 2280 34400
rect 3056 34391 3108 34400
rect 3056 34357 3065 34391
rect 3065 34357 3099 34391
rect 3099 34357 3108 34391
rect 3056 34348 3108 34357
rect 2582 34246 2634 34298
rect 2646 34246 2698 34298
rect 2710 34246 2762 34298
rect 2774 34246 2826 34298
rect 2838 34246 2890 34298
rect 5846 34246 5898 34298
rect 5910 34246 5962 34298
rect 5974 34246 6026 34298
rect 6038 34246 6090 34298
rect 6102 34246 6154 34298
rect 9110 34246 9162 34298
rect 9174 34246 9226 34298
rect 9238 34246 9290 34298
rect 9302 34246 9354 34298
rect 9366 34246 9418 34298
rect 848 34144 900 34196
rect 8576 34144 8628 34196
rect 204 34076 256 34128
rect 5632 34076 5684 34128
rect 5816 34076 5868 34128
rect 848 33940 900 33992
rect 5632 33940 5684 33992
rect 6276 33940 6328 33992
rect 2136 33872 2188 33924
rect 2964 33872 3016 33924
rect 2412 33804 2464 33856
rect 6368 33804 6420 33856
rect 4214 33702 4266 33754
rect 4278 33702 4330 33754
rect 4342 33702 4394 33754
rect 4406 33702 4458 33754
rect 4470 33702 4522 33754
rect 7478 33702 7530 33754
rect 7542 33702 7594 33754
rect 7606 33702 7658 33754
rect 7670 33702 7722 33754
rect 7734 33702 7786 33754
rect 1860 33600 1912 33652
rect 2136 33643 2188 33652
rect 2136 33609 2145 33643
rect 2145 33609 2179 33643
rect 2179 33609 2188 33643
rect 2136 33600 2188 33609
rect 2964 33643 3016 33652
rect 2964 33609 2973 33643
rect 2973 33609 3007 33643
rect 3007 33609 3016 33643
rect 2964 33600 3016 33609
rect 3976 33600 4028 33652
rect 5540 33600 5592 33652
rect 8760 33600 8812 33652
rect 1400 33532 1452 33584
rect 2412 33532 2464 33584
rect 1952 33507 2004 33516
rect 1952 33473 1961 33507
rect 1961 33473 1995 33507
rect 1995 33473 2004 33507
rect 1952 33464 2004 33473
rect 1032 33328 1084 33380
rect 1860 33328 1912 33380
rect 1952 33328 2004 33380
rect 2412 33328 2464 33380
rect 2964 33260 3016 33312
rect 5632 33464 5684 33516
rect 9864 33507 9916 33516
rect 9864 33473 9873 33507
rect 9873 33473 9907 33507
rect 9907 33473 9916 33507
rect 9864 33464 9916 33473
rect 4620 33396 4672 33448
rect 5632 33328 5684 33380
rect 5816 33328 5868 33380
rect 10048 33371 10100 33380
rect 10048 33337 10057 33371
rect 10057 33337 10091 33371
rect 10091 33337 10100 33371
rect 10048 33328 10100 33337
rect 2582 33158 2634 33210
rect 2646 33158 2698 33210
rect 2710 33158 2762 33210
rect 2774 33158 2826 33210
rect 2838 33158 2890 33210
rect 5846 33158 5898 33210
rect 5910 33158 5962 33210
rect 5974 33158 6026 33210
rect 6038 33158 6090 33210
rect 6102 33158 6154 33210
rect 9110 33158 9162 33210
rect 9174 33158 9226 33210
rect 9238 33158 9290 33210
rect 9302 33158 9354 33210
rect 9366 33158 9418 33210
rect 296 33056 348 33108
rect 3148 33099 3200 33108
rect 3148 33065 3157 33099
rect 3157 33065 3191 33099
rect 3191 33065 3200 33099
rect 3148 33056 3200 33065
rect 3700 32988 3752 33040
rect 1676 32920 1728 32972
rect 2320 32852 2372 32904
rect 2596 32784 2648 32836
rect 2964 32895 3016 32904
rect 2964 32861 2973 32895
rect 2973 32861 3007 32895
rect 3007 32861 3016 32895
rect 9680 32920 9732 32972
rect 2964 32852 3016 32861
rect 7840 32852 7892 32904
rect 3976 32759 4028 32768
rect 3976 32725 3985 32759
rect 3985 32725 4019 32759
rect 4019 32725 4028 32759
rect 3976 32716 4028 32725
rect 10048 32759 10100 32768
rect 10048 32725 10057 32759
rect 10057 32725 10091 32759
rect 10091 32725 10100 32759
rect 10048 32716 10100 32725
rect 4214 32614 4266 32666
rect 4278 32614 4330 32666
rect 4342 32614 4394 32666
rect 4406 32614 4458 32666
rect 4470 32614 4522 32666
rect 7478 32614 7530 32666
rect 7542 32614 7594 32666
rect 7606 32614 7658 32666
rect 7670 32614 7722 32666
rect 7734 32614 7786 32666
rect 756 32512 808 32564
rect 2596 32555 2648 32564
rect 2596 32521 2605 32555
rect 2605 32521 2639 32555
rect 2639 32521 2648 32555
rect 2596 32512 2648 32521
rect 3240 32555 3292 32564
rect 3240 32521 3249 32555
rect 3249 32521 3283 32555
rect 3283 32521 3292 32555
rect 3240 32512 3292 32521
rect 1768 32376 1820 32428
rect 1860 32376 1912 32428
rect 3700 32376 3752 32428
rect 4436 32444 4488 32496
rect 4804 32444 4856 32496
rect 848 32308 900 32360
rect 3240 32308 3292 32360
rect 3424 32308 3476 32360
rect 5632 32240 5684 32292
rect 3976 32215 4028 32224
rect 3976 32181 3985 32215
rect 3985 32181 4019 32215
rect 4019 32181 4028 32215
rect 3976 32172 4028 32181
rect 2582 32070 2634 32122
rect 2646 32070 2698 32122
rect 2710 32070 2762 32122
rect 2774 32070 2826 32122
rect 2838 32070 2890 32122
rect 5846 32070 5898 32122
rect 5910 32070 5962 32122
rect 5974 32070 6026 32122
rect 6038 32070 6090 32122
rect 6102 32070 6154 32122
rect 9110 32070 9162 32122
rect 9174 32070 9226 32122
rect 9238 32070 9290 32122
rect 9302 32070 9354 32122
rect 9366 32070 9418 32122
rect 1768 32011 1820 32020
rect 1768 31977 1777 32011
rect 1777 31977 1811 32011
rect 1811 31977 1820 32011
rect 1768 31968 1820 31977
rect 940 31900 992 31952
rect 1676 31900 1728 31952
rect 2412 31968 2464 32020
rect 4620 31968 4672 32020
rect 4896 31968 4948 32020
rect 2044 31900 2096 31952
rect 1492 31764 1544 31816
rect 1860 31764 1912 31816
rect 2688 31900 2740 31952
rect 3424 31900 3476 31952
rect 3884 31900 3936 31952
rect 4436 31832 4488 31884
rect 2412 31764 2464 31816
rect 2780 31807 2832 31816
rect 1676 31696 1728 31748
rect 2136 31696 2188 31748
rect 940 31628 992 31680
rect 1768 31628 1820 31680
rect 1860 31628 1912 31680
rect 2780 31773 2789 31807
rect 2789 31773 2823 31807
rect 2823 31773 2832 31807
rect 2780 31764 2832 31773
rect 3332 31764 3384 31816
rect 4804 31764 4856 31816
rect 3332 31628 3384 31680
rect 4712 31628 4764 31680
rect 10048 31943 10100 31952
rect 10048 31909 10057 31943
rect 10057 31909 10091 31943
rect 10091 31909 10100 31943
rect 10048 31900 10100 31909
rect 7932 31764 7984 31816
rect 4214 31526 4266 31578
rect 4278 31526 4330 31578
rect 4342 31526 4394 31578
rect 4406 31526 4458 31578
rect 4470 31526 4522 31578
rect 7478 31526 7530 31578
rect 7542 31526 7594 31578
rect 7606 31526 7658 31578
rect 7670 31526 7722 31578
rect 7734 31526 7786 31578
rect 572 31424 624 31476
rect 1032 31424 1084 31476
rect 3056 31424 3108 31476
rect 3240 31424 3292 31476
rect 5080 31424 5132 31476
rect 5264 31424 5316 31476
rect 6184 31356 6236 31408
rect 2044 31331 2096 31340
rect 2044 31297 2053 31331
rect 2053 31297 2087 31331
rect 2087 31297 2096 31331
rect 2044 31288 2096 31297
rect 2320 31288 2372 31340
rect 2596 31288 2648 31340
rect 3608 31288 3660 31340
rect 5080 31288 5132 31340
rect 2228 31084 2280 31136
rect 3608 31195 3660 31204
rect 3608 31161 3617 31195
rect 3617 31161 3651 31195
rect 3651 31161 3660 31195
rect 3608 31152 3660 31161
rect 2964 31084 3016 31136
rect 10048 31127 10100 31136
rect 10048 31093 10057 31127
rect 10057 31093 10091 31127
rect 10091 31093 10100 31127
rect 10048 31084 10100 31093
rect 2582 30982 2634 31034
rect 2646 30982 2698 31034
rect 2710 30982 2762 31034
rect 2774 30982 2826 31034
rect 2838 30982 2890 31034
rect 5846 30982 5898 31034
rect 5910 30982 5962 31034
rect 5974 30982 6026 31034
rect 6038 30982 6090 31034
rect 6102 30982 6154 31034
rect 9110 30982 9162 31034
rect 9174 30982 9226 31034
rect 9238 30982 9290 31034
rect 9302 30982 9354 31034
rect 9366 30982 9418 31034
rect 2044 30880 2096 30932
rect 1492 30744 1544 30796
rect 1860 30744 1912 30796
rect 2044 30744 2096 30796
rect 756 30676 808 30728
rect 8392 30676 8444 30728
rect 1492 30651 1544 30660
rect 1492 30617 1501 30651
rect 1501 30617 1535 30651
rect 1535 30617 1544 30651
rect 1492 30608 1544 30617
rect 6460 30608 6512 30660
rect 10048 30583 10100 30592
rect 10048 30549 10057 30583
rect 10057 30549 10091 30583
rect 10091 30549 10100 30583
rect 10048 30540 10100 30549
rect 4214 30438 4266 30490
rect 4278 30438 4330 30490
rect 4342 30438 4394 30490
rect 4406 30438 4458 30490
rect 4470 30438 4522 30490
rect 7478 30438 7530 30490
rect 7542 30438 7594 30490
rect 7606 30438 7658 30490
rect 7670 30438 7722 30490
rect 7734 30438 7786 30490
rect 1860 30243 1912 30252
rect 1860 30209 1869 30243
rect 1869 30209 1903 30243
rect 1903 30209 1912 30243
rect 1860 30200 1912 30209
rect 2596 30200 2648 30252
rect 8668 30132 8720 30184
rect 2780 30064 2832 30116
rect 2582 29894 2634 29946
rect 2646 29894 2698 29946
rect 2710 29894 2762 29946
rect 2774 29894 2826 29946
rect 2838 29894 2890 29946
rect 5846 29894 5898 29946
rect 5910 29894 5962 29946
rect 5974 29894 6026 29946
rect 6038 29894 6090 29946
rect 6102 29894 6154 29946
rect 9110 29894 9162 29946
rect 9174 29894 9226 29946
rect 9238 29894 9290 29946
rect 9302 29894 9354 29946
rect 9366 29894 9418 29946
rect 8392 29792 8444 29844
rect 2044 29767 2096 29776
rect 2044 29733 2053 29767
rect 2053 29733 2087 29767
rect 2087 29733 2096 29767
rect 2044 29724 2096 29733
rect 1400 29588 1452 29640
rect 2044 29588 2096 29640
rect 3240 29588 3292 29640
rect 10140 29631 10192 29640
rect 10140 29597 10149 29631
rect 10149 29597 10183 29631
rect 10183 29597 10192 29631
rect 10140 29588 10192 29597
rect 1492 29520 1544 29572
rect 4214 29350 4266 29402
rect 4278 29350 4330 29402
rect 4342 29350 4394 29402
rect 4406 29350 4458 29402
rect 4470 29350 4522 29402
rect 7478 29350 7530 29402
rect 7542 29350 7594 29402
rect 7606 29350 7658 29402
rect 7670 29350 7722 29402
rect 7734 29350 7786 29402
rect 664 29248 716 29300
rect 3884 29180 3936 29232
rect 1400 29112 1452 29164
rect 2964 29112 3016 29164
rect 1768 29044 1820 29096
rect 4068 29044 4120 29096
rect 2872 28976 2924 29028
rect 3884 28976 3936 29028
rect 10140 29019 10192 29028
rect 10140 28985 10149 29019
rect 10149 28985 10183 29019
rect 10183 28985 10192 29019
rect 10140 28976 10192 28985
rect 2504 28908 2556 28960
rect 2582 28806 2634 28858
rect 2646 28806 2698 28858
rect 2710 28806 2762 28858
rect 2774 28806 2826 28858
rect 2838 28806 2890 28858
rect 5846 28806 5898 28858
rect 5910 28806 5962 28858
rect 5974 28806 6026 28858
rect 6038 28806 6090 28858
rect 6102 28806 6154 28858
rect 9110 28806 9162 28858
rect 9174 28806 9226 28858
rect 9238 28806 9290 28858
rect 9302 28806 9354 28858
rect 9366 28806 9418 28858
rect 2504 28704 2556 28756
rect 9864 28704 9916 28756
rect 1768 28636 1820 28688
rect 2964 28636 3016 28688
rect 2412 28543 2464 28552
rect 2412 28509 2421 28543
rect 2421 28509 2455 28543
rect 2455 28509 2464 28543
rect 2412 28500 2464 28509
rect 2596 28543 2648 28552
rect 2596 28509 2605 28543
rect 2605 28509 2639 28543
rect 2639 28509 2648 28543
rect 2596 28500 2648 28509
rect 1768 28475 1820 28484
rect 1768 28441 1777 28475
rect 1777 28441 1811 28475
rect 1811 28441 1820 28475
rect 1768 28432 1820 28441
rect 1952 28475 2004 28484
rect 1952 28441 1961 28475
rect 1961 28441 1995 28475
rect 1995 28441 2004 28475
rect 1952 28432 2004 28441
rect 2320 28432 2372 28484
rect 4214 28262 4266 28314
rect 4278 28262 4330 28314
rect 4342 28262 4394 28314
rect 4406 28262 4458 28314
rect 4470 28262 4522 28314
rect 7478 28262 7530 28314
rect 7542 28262 7594 28314
rect 7606 28262 7658 28314
rect 7670 28262 7722 28314
rect 7734 28262 7786 28314
rect 1768 28160 1820 28212
rect 3056 28092 3108 28144
rect 756 28024 808 28076
rect 2964 28024 3016 28076
rect 3056 27956 3108 28008
rect 9956 27999 10008 28008
rect 9956 27965 9965 27999
rect 9965 27965 9999 27999
rect 9999 27965 10008 27999
rect 9956 27956 10008 27965
rect 2582 27718 2634 27770
rect 2646 27718 2698 27770
rect 2710 27718 2762 27770
rect 2774 27718 2826 27770
rect 2838 27718 2890 27770
rect 5846 27718 5898 27770
rect 5910 27718 5962 27770
rect 5974 27718 6026 27770
rect 6038 27718 6090 27770
rect 6102 27718 6154 27770
rect 9110 27718 9162 27770
rect 9174 27718 9226 27770
rect 9238 27718 9290 27770
rect 9302 27718 9354 27770
rect 9366 27718 9418 27770
rect 1032 27548 1084 27600
rect 3332 27480 3384 27532
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 3056 27344 3108 27396
rect 9956 27319 10008 27328
rect 9956 27285 9965 27319
rect 9965 27285 9999 27319
rect 9999 27285 10008 27319
rect 9956 27276 10008 27285
rect 4214 27174 4266 27226
rect 4278 27174 4330 27226
rect 4342 27174 4394 27226
rect 4406 27174 4458 27226
rect 4470 27174 4522 27226
rect 7478 27174 7530 27226
rect 7542 27174 7594 27226
rect 7606 27174 7658 27226
rect 7670 27174 7722 27226
rect 7734 27174 7786 27226
rect 756 27004 808 27056
rect 2044 26936 2096 26988
rect 4528 27004 4580 27056
rect 2136 26911 2188 26920
rect 2136 26877 2145 26911
rect 2145 26877 2179 26911
rect 2179 26877 2188 26911
rect 2136 26868 2188 26877
rect 1676 26843 1728 26852
rect 1676 26809 1685 26843
rect 1685 26809 1719 26843
rect 1719 26809 1728 26843
rect 1676 26800 1728 26809
rect 10140 26775 10192 26784
rect 10140 26741 10149 26775
rect 10149 26741 10183 26775
rect 10183 26741 10192 26775
rect 10140 26732 10192 26741
rect 2582 26630 2634 26682
rect 2646 26630 2698 26682
rect 2710 26630 2762 26682
rect 2774 26630 2826 26682
rect 2838 26630 2890 26682
rect 5846 26630 5898 26682
rect 5910 26630 5962 26682
rect 5974 26630 6026 26682
rect 6038 26630 6090 26682
rect 6102 26630 6154 26682
rect 9110 26630 9162 26682
rect 9174 26630 9226 26682
rect 9238 26630 9290 26682
rect 9302 26630 9354 26682
rect 9366 26630 9418 26682
rect 2044 26571 2096 26580
rect 2044 26537 2053 26571
rect 2053 26537 2087 26571
rect 2087 26537 2096 26571
rect 2044 26528 2096 26537
rect 1676 26460 1728 26512
rect 2136 26460 2188 26512
rect 3148 26460 3200 26512
rect 756 26392 808 26444
rect 940 26324 992 26376
rect 1492 26324 1544 26376
rect 2596 26299 2648 26308
rect 2596 26265 2605 26299
rect 2605 26265 2639 26299
rect 2639 26265 2648 26299
rect 2596 26256 2648 26265
rect 3056 26188 3108 26240
rect 3332 26188 3384 26240
rect 4214 26086 4266 26138
rect 4278 26086 4330 26138
rect 4342 26086 4394 26138
rect 4406 26086 4458 26138
rect 4470 26086 4522 26138
rect 7478 26086 7530 26138
rect 7542 26086 7594 26138
rect 7606 26086 7658 26138
rect 7670 26086 7722 26138
rect 7734 26086 7786 26138
rect 20 25984 72 26036
rect 3424 26027 3476 26036
rect 3424 25993 3433 26027
rect 3433 25993 3467 26027
rect 3467 25993 3476 26027
rect 3424 25984 3476 25993
rect 3608 25916 3660 25968
rect 2044 25848 2096 25900
rect 2964 25848 3016 25900
rect 3332 25891 3384 25900
rect 3332 25857 3341 25891
rect 3341 25857 3375 25891
rect 3375 25857 3384 25891
rect 3332 25848 3384 25857
rect 10140 25687 10192 25696
rect 10140 25653 10149 25687
rect 10149 25653 10183 25687
rect 10183 25653 10192 25687
rect 10140 25644 10192 25653
rect 2582 25542 2634 25594
rect 2646 25542 2698 25594
rect 2710 25542 2762 25594
rect 2774 25542 2826 25594
rect 2838 25542 2890 25594
rect 5846 25542 5898 25594
rect 5910 25542 5962 25594
rect 5974 25542 6026 25594
rect 6038 25542 6090 25594
rect 6102 25542 6154 25594
rect 9110 25542 9162 25594
rect 9174 25542 9226 25594
rect 9238 25542 9290 25594
rect 9302 25542 9354 25594
rect 9366 25542 9418 25594
rect 1860 25440 1912 25492
rect 3792 25440 3844 25492
rect 3056 25372 3108 25424
rect 10140 25279 10192 25288
rect 10140 25245 10149 25279
rect 10149 25245 10183 25279
rect 10183 25245 10192 25279
rect 10140 25236 10192 25245
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 3884 25211 3936 25220
rect 3884 25177 3893 25211
rect 3893 25177 3927 25211
rect 3927 25177 3936 25211
rect 3884 25168 3936 25177
rect 2872 25100 2924 25152
rect 4214 24998 4266 25050
rect 4278 24998 4330 25050
rect 4342 24998 4394 25050
rect 4406 24998 4458 25050
rect 4470 24998 4522 25050
rect 7478 24998 7530 25050
rect 7542 24998 7594 25050
rect 7606 24998 7658 25050
rect 7670 24998 7722 25050
rect 7734 24998 7786 25050
rect 2320 24828 2372 24880
rect 1124 24692 1176 24744
rect 2136 24692 2188 24744
rect 2964 24760 3016 24812
rect 3240 24692 3292 24744
rect 3792 24556 3844 24608
rect 2582 24454 2634 24506
rect 2646 24454 2698 24506
rect 2710 24454 2762 24506
rect 2774 24454 2826 24506
rect 2838 24454 2890 24506
rect 5846 24454 5898 24506
rect 5910 24454 5962 24506
rect 5974 24454 6026 24506
rect 6038 24454 6090 24506
rect 6102 24454 6154 24506
rect 9110 24454 9162 24506
rect 9174 24454 9226 24506
rect 9238 24454 9290 24506
rect 9302 24454 9354 24506
rect 9366 24454 9418 24506
rect 2228 24284 2280 24336
rect 3792 24259 3844 24268
rect 3792 24225 3801 24259
rect 3801 24225 3835 24259
rect 3835 24225 3844 24259
rect 3792 24216 3844 24225
rect 7840 24216 7892 24268
rect 2688 24191 2740 24200
rect 2688 24157 2697 24191
rect 2697 24157 2731 24191
rect 2731 24157 2740 24191
rect 2688 24148 2740 24157
rect 2964 24148 3016 24200
rect 10140 24191 10192 24200
rect 10140 24157 10149 24191
rect 10149 24157 10183 24191
rect 10183 24157 10192 24191
rect 10140 24148 10192 24157
rect 3056 24080 3108 24132
rect 3792 24012 3844 24064
rect 4214 23910 4266 23962
rect 4278 23910 4330 23962
rect 4342 23910 4394 23962
rect 4406 23910 4458 23962
rect 4470 23910 4522 23962
rect 7478 23910 7530 23962
rect 7542 23910 7594 23962
rect 7606 23910 7658 23962
rect 7670 23910 7722 23962
rect 7734 23910 7786 23962
rect 3056 23851 3108 23860
rect 3056 23817 3065 23851
rect 3065 23817 3099 23851
rect 3099 23817 3108 23851
rect 3056 23808 3108 23817
rect 3976 23808 4028 23860
rect 5080 23851 5132 23860
rect 5080 23817 5089 23851
rect 5089 23817 5123 23851
rect 5123 23817 5132 23851
rect 5080 23808 5132 23817
rect 5264 23808 5316 23860
rect 756 23740 808 23792
rect 1584 23672 1636 23724
rect 3056 23672 3108 23724
rect 3792 23715 3844 23724
rect 3792 23681 3801 23715
rect 3801 23681 3835 23715
rect 3835 23681 3844 23715
rect 3792 23672 3844 23681
rect 1124 23604 1176 23656
rect 2780 23604 2832 23656
rect 3332 23604 3384 23656
rect 3792 23536 3844 23588
rect 4528 23740 4580 23792
rect 4896 23672 4948 23724
rect 5080 23672 5132 23724
rect 5264 23715 5316 23724
rect 5264 23681 5273 23715
rect 5273 23681 5307 23715
rect 5307 23681 5316 23715
rect 5264 23672 5316 23681
rect 7932 23604 7984 23656
rect 3240 23468 3292 23520
rect 4068 23468 4120 23520
rect 10140 23511 10192 23520
rect 10140 23477 10149 23511
rect 10149 23477 10183 23511
rect 10183 23477 10192 23511
rect 10140 23468 10192 23477
rect 2582 23366 2634 23418
rect 2646 23366 2698 23418
rect 2710 23366 2762 23418
rect 2774 23366 2826 23418
rect 2838 23366 2890 23418
rect 5846 23366 5898 23418
rect 5910 23366 5962 23418
rect 5974 23366 6026 23418
rect 6038 23366 6090 23418
rect 6102 23366 6154 23418
rect 9110 23366 9162 23418
rect 9174 23366 9226 23418
rect 9238 23366 9290 23418
rect 9302 23366 9354 23418
rect 9366 23366 9418 23418
rect 4160 23264 4212 23316
rect 4988 23264 5040 23316
rect 5724 23196 5776 23248
rect 3056 23128 3108 23180
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2136 23060 2188 23112
rect 3884 23060 3936 23112
rect 4528 22992 4580 23044
rect 1768 22924 1820 22976
rect 2320 22924 2372 22976
rect 4712 22924 4764 22976
rect 4214 22822 4266 22874
rect 4278 22822 4330 22874
rect 4342 22822 4394 22874
rect 4406 22822 4458 22874
rect 4470 22822 4522 22874
rect 7478 22822 7530 22874
rect 7542 22822 7594 22874
rect 7606 22822 7658 22874
rect 7670 22822 7722 22874
rect 7734 22822 7786 22874
rect 3056 22720 3108 22772
rect 3240 22720 3292 22772
rect 3516 22720 3568 22772
rect 5264 22652 5316 22704
rect 3516 22627 3568 22636
rect 2320 22516 2372 22568
rect 3516 22593 3525 22627
rect 3525 22593 3559 22627
rect 3559 22593 3568 22627
rect 3516 22584 3568 22593
rect 2964 22516 3016 22568
rect 3056 22448 3108 22500
rect 10140 22491 10192 22500
rect 10140 22457 10149 22491
rect 10149 22457 10183 22491
rect 10183 22457 10192 22491
rect 10140 22448 10192 22457
rect 3148 22380 3200 22432
rect 3976 22380 4028 22432
rect 2582 22278 2634 22330
rect 2646 22278 2698 22330
rect 2710 22278 2762 22330
rect 2774 22278 2826 22330
rect 2838 22278 2890 22330
rect 5846 22278 5898 22330
rect 5910 22278 5962 22330
rect 5974 22278 6026 22330
rect 6038 22278 6090 22330
rect 6102 22278 6154 22330
rect 9110 22278 9162 22330
rect 9174 22278 9226 22330
rect 9238 22278 9290 22330
rect 9302 22278 9354 22330
rect 9366 22278 9418 22330
rect 2320 22176 2372 22228
rect 3148 22176 3200 22228
rect 3608 22176 3660 22228
rect 2228 22108 2280 22160
rect 10140 22151 10192 22160
rect 10140 22117 10149 22151
rect 10149 22117 10183 22151
rect 10183 22117 10192 22151
rect 10140 22108 10192 22117
rect 1952 22040 2004 22092
rect 2136 22040 2188 22092
rect 2320 22040 2372 22092
rect 5080 22040 5132 22092
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 3056 21972 3108 22024
rect 4214 21734 4266 21786
rect 4278 21734 4330 21786
rect 4342 21734 4394 21786
rect 4406 21734 4458 21786
rect 4470 21734 4522 21786
rect 7478 21734 7530 21786
rect 7542 21734 7594 21786
rect 7606 21734 7658 21786
rect 7670 21734 7722 21786
rect 7734 21734 7786 21786
rect 4804 21632 4856 21684
rect 5448 21564 5500 21616
rect 3056 21496 3108 21548
rect 4804 21496 4856 21548
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 3976 21428 4028 21480
rect 10140 21335 10192 21344
rect 10140 21301 10149 21335
rect 10149 21301 10183 21335
rect 10183 21301 10192 21335
rect 10140 21292 10192 21301
rect 2582 21190 2634 21242
rect 2646 21190 2698 21242
rect 2710 21190 2762 21242
rect 2774 21190 2826 21242
rect 2838 21190 2890 21242
rect 5846 21190 5898 21242
rect 5910 21190 5962 21242
rect 5974 21190 6026 21242
rect 6038 21190 6090 21242
rect 6102 21190 6154 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 9238 21190 9290 21242
rect 9302 21190 9354 21242
rect 9366 21190 9418 21242
rect 3424 21088 3476 21140
rect 1032 21020 1084 21072
rect 1216 20952 1268 21004
rect 1952 20884 2004 20936
rect 2964 20884 3016 20936
rect 3424 20884 3476 20936
rect 4214 20646 4266 20698
rect 4278 20646 4330 20698
rect 4342 20646 4394 20698
rect 4406 20646 4458 20698
rect 4470 20646 4522 20698
rect 7478 20646 7530 20698
rect 7542 20646 7594 20698
rect 7606 20646 7658 20698
rect 7670 20646 7722 20698
rect 7734 20646 7786 20698
rect 1676 20451 1728 20460
rect 1676 20417 1685 20451
rect 1685 20417 1719 20451
rect 1719 20417 1728 20451
rect 1676 20408 1728 20417
rect 2780 20408 2832 20460
rect 3148 20408 3200 20460
rect 10140 20408 10192 20460
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 10048 20315 10100 20324
rect 10048 20281 10057 20315
rect 10057 20281 10091 20315
rect 10091 20281 10100 20315
rect 10048 20272 10100 20281
rect 2582 20102 2634 20154
rect 2646 20102 2698 20154
rect 2710 20102 2762 20154
rect 2774 20102 2826 20154
rect 2838 20102 2890 20154
rect 5846 20102 5898 20154
rect 5910 20102 5962 20154
rect 5974 20102 6026 20154
rect 6038 20102 6090 20154
rect 6102 20102 6154 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 9238 20102 9290 20154
rect 9302 20102 9354 20154
rect 9366 20102 9418 20154
rect 3056 20043 3108 20052
rect 3056 20009 3065 20043
rect 3065 20009 3099 20043
rect 3099 20009 3108 20043
rect 3056 20000 3108 20009
rect 1584 19864 1636 19916
rect 1768 19864 1820 19916
rect 2136 19864 2188 19916
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 3240 19796 3292 19848
rect 9220 19796 9272 19848
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 4214 19558 4266 19610
rect 4278 19558 4330 19610
rect 4342 19558 4394 19610
rect 4406 19558 4458 19610
rect 4470 19558 4522 19610
rect 7478 19558 7530 19610
rect 7542 19558 7594 19610
rect 7606 19558 7658 19610
rect 7670 19558 7722 19610
rect 7734 19558 7786 19610
rect 9220 19499 9272 19508
rect 9220 19465 9229 19499
rect 9229 19465 9263 19499
rect 9263 19465 9272 19499
rect 9220 19456 9272 19465
rect 3608 19388 3660 19440
rect 1492 19320 1544 19372
rect 2964 19320 3016 19372
rect 3516 19320 3568 19372
rect 1400 19295 1452 19304
rect 1400 19261 1409 19295
rect 1409 19261 1443 19295
rect 1443 19261 1452 19295
rect 1400 19252 1452 19261
rect 5172 19184 5224 19236
rect 9864 19159 9916 19168
rect 9864 19125 9873 19159
rect 9873 19125 9907 19159
rect 9907 19125 9916 19159
rect 9864 19116 9916 19125
rect 2582 19014 2634 19066
rect 2646 19014 2698 19066
rect 2710 19014 2762 19066
rect 2774 19014 2826 19066
rect 2838 19014 2890 19066
rect 5846 19014 5898 19066
rect 5910 19014 5962 19066
rect 5974 19014 6026 19066
rect 6038 19014 6090 19066
rect 6102 19014 6154 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 9238 19014 9290 19066
rect 9302 19014 9354 19066
rect 9366 19014 9418 19066
rect 2136 18912 2188 18964
rect 1216 18776 1268 18828
rect 2504 18776 2556 18828
rect 2780 18776 2832 18828
rect 3240 18776 3292 18828
rect 3976 18751 4028 18760
rect 3976 18717 3985 18751
rect 3985 18717 4019 18751
rect 4019 18717 4028 18751
rect 3976 18708 4028 18717
rect 9864 18751 9916 18760
rect 9864 18717 9873 18751
rect 9873 18717 9907 18751
rect 9907 18717 9916 18751
rect 9864 18708 9916 18717
rect 3240 18640 3292 18692
rect 3884 18640 3936 18692
rect 10048 18615 10100 18624
rect 10048 18581 10057 18615
rect 10057 18581 10091 18615
rect 10091 18581 10100 18615
rect 10048 18572 10100 18581
rect 4214 18470 4266 18522
rect 4278 18470 4330 18522
rect 4342 18470 4394 18522
rect 4406 18470 4458 18522
rect 4470 18470 4522 18522
rect 7478 18470 7530 18522
rect 7542 18470 7594 18522
rect 7606 18470 7658 18522
rect 7670 18470 7722 18522
rect 7734 18470 7786 18522
rect 2964 18368 3016 18420
rect 1952 18300 2004 18352
rect 3148 18300 3200 18352
rect 2688 18232 2740 18284
rect 3700 18275 3752 18284
rect 2320 18164 2372 18216
rect 3700 18241 3709 18275
rect 3709 18241 3743 18275
rect 3743 18241 3752 18275
rect 3700 18232 3752 18241
rect 9864 18275 9916 18284
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 2504 18139 2556 18148
rect 2504 18105 2513 18139
rect 2513 18105 2547 18139
rect 2547 18105 2556 18139
rect 2504 18096 2556 18105
rect 3056 18164 3108 18216
rect 2964 18028 3016 18080
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 2582 17926 2634 17978
rect 2646 17926 2698 17978
rect 2710 17926 2762 17978
rect 2774 17926 2826 17978
rect 2838 17926 2890 17978
rect 5846 17926 5898 17978
rect 5910 17926 5962 17978
rect 5974 17926 6026 17978
rect 6038 17926 6090 17978
rect 6102 17926 6154 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 9238 17926 9290 17978
rect 9302 17926 9354 17978
rect 9366 17926 9418 17978
rect 1952 17824 2004 17876
rect 3608 17824 3660 17876
rect 3884 17756 3936 17808
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 2504 17620 2556 17672
rect 3056 17688 3108 17740
rect 3148 17663 3200 17672
rect 3148 17629 3157 17663
rect 3157 17629 3191 17663
rect 3191 17629 3200 17663
rect 3148 17620 3200 17629
rect 9036 17620 9088 17672
rect 1676 17552 1728 17604
rect 3516 17552 3568 17604
rect 3976 17527 4028 17536
rect 3976 17493 4001 17527
rect 4001 17493 4028 17527
rect 10048 17527 10100 17536
rect 3976 17484 4028 17493
rect 10048 17493 10057 17527
rect 10057 17493 10091 17527
rect 10091 17493 10100 17527
rect 10048 17484 10100 17493
rect 4214 17382 4266 17434
rect 4278 17382 4330 17434
rect 4342 17382 4394 17434
rect 4406 17382 4458 17434
rect 4470 17382 4522 17434
rect 7478 17382 7530 17434
rect 7542 17382 7594 17434
rect 7606 17382 7658 17434
rect 7670 17382 7722 17434
rect 7734 17382 7786 17434
rect 1124 17280 1176 17332
rect 4712 17280 4764 17332
rect 4988 17280 5040 17332
rect 9864 17280 9916 17332
rect 3884 17212 3936 17264
rect 2964 17187 3016 17196
rect 2964 17153 2973 17187
rect 2973 17153 3007 17187
rect 3007 17153 3016 17187
rect 2964 17144 3016 17153
rect 3976 17144 4028 17196
rect 3240 17119 3292 17128
rect 3240 17085 3249 17119
rect 3249 17085 3283 17119
rect 3283 17085 3292 17119
rect 3240 17076 3292 17085
rect 4620 16940 4672 16992
rect 4804 16940 4856 16992
rect 2582 16838 2634 16890
rect 2646 16838 2698 16890
rect 2710 16838 2762 16890
rect 2774 16838 2826 16890
rect 2838 16838 2890 16890
rect 5846 16838 5898 16890
rect 5910 16838 5962 16890
rect 5974 16838 6026 16890
rect 6038 16838 6090 16890
rect 6102 16838 6154 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 9238 16838 9290 16890
rect 9302 16838 9354 16890
rect 9366 16838 9418 16890
rect 1216 16532 1268 16584
rect 2412 16575 2464 16584
rect 2412 16541 2421 16575
rect 2421 16541 2455 16575
rect 2455 16541 2464 16575
rect 2412 16532 2464 16541
rect 3056 16575 3108 16584
rect 3056 16541 3065 16575
rect 3065 16541 3099 16575
rect 3099 16541 3108 16575
rect 3056 16532 3108 16541
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 9220 16532 9272 16584
rect 1584 16396 1636 16448
rect 2228 16439 2280 16448
rect 2228 16405 2237 16439
rect 2237 16405 2271 16439
rect 2271 16405 2280 16439
rect 2228 16396 2280 16405
rect 3332 16464 3384 16516
rect 3240 16396 3292 16448
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 4214 16294 4266 16346
rect 4278 16294 4330 16346
rect 4342 16294 4394 16346
rect 4406 16294 4458 16346
rect 4470 16294 4522 16346
rect 7478 16294 7530 16346
rect 7542 16294 7594 16346
rect 7606 16294 7658 16346
rect 7670 16294 7722 16346
rect 7734 16294 7786 16346
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 1400 16056 1452 16108
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 2872 16099 2924 16108
rect 2872 16065 2881 16099
rect 2881 16065 2915 16099
rect 2915 16065 2924 16099
rect 2872 16056 2924 16065
rect 3700 16056 3752 16108
rect 9956 16056 10008 16108
rect 1492 15852 1544 15904
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 2136 15852 2188 15904
rect 10048 15895 10100 15904
rect 10048 15861 10057 15895
rect 10057 15861 10091 15895
rect 10091 15861 10100 15895
rect 10048 15852 10100 15861
rect 2582 15750 2634 15802
rect 2646 15750 2698 15802
rect 2710 15750 2762 15802
rect 2774 15750 2826 15802
rect 2838 15750 2890 15802
rect 5846 15750 5898 15802
rect 5910 15750 5962 15802
rect 5974 15750 6026 15802
rect 6038 15750 6090 15802
rect 6102 15750 6154 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 9238 15750 9290 15802
rect 9302 15750 9354 15802
rect 9366 15750 9418 15802
rect 2136 15648 2188 15700
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 4988 15580 5040 15632
rect 2044 15512 2096 15564
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 3240 15444 3292 15496
rect 3516 15376 3568 15428
rect 2136 15351 2188 15360
rect 2136 15317 2145 15351
rect 2145 15317 2179 15351
rect 2179 15317 2188 15351
rect 2136 15308 2188 15317
rect 2412 15308 2464 15360
rect 4214 15206 4266 15258
rect 4278 15206 4330 15258
rect 4342 15206 4394 15258
rect 4406 15206 4458 15258
rect 4470 15206 4522 15258
rect 7478 15206 7530 15258
rect 7542 15206 7594 15258
rect 7606 15206 7658 15258
rect 7670 15206 7722 15258
rect 7734 15206 7786 15258
rect 8576 15104 8628 15156
rect 3056 15036 3108 15088
rect 2964 14968 3016 15020
rect 9496 14968 9548 15020
rect 10048 14875 10100 14884
rect 10048 14841 10057 14875
rect 10057 14841 10091 14875
rect 10091 14841 10100 14875
rect 10048 14832 10100 14841
rect 1676 14764 1728 14816
rect 2582 14662 2634 14714
rect 2646 14662 2698 14714
rect 2710 14662 2762 14714
rect 2774 14662 2826 14714
rect 2838 14662 2890 14714
rect 5846 14662 5898 14714
rect 5910 14662 5962 14714
rect 5974 14662 6026 14714
rect 6038 14662 6090 14714
rect 6102 14662 6154 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 9238 14662 9290 14714
rect 9302 14662 9354 14714
rect 9366 14662 9418 14714
rect 1768 14560 1820 14612
rect 2504 14560 2556 14612
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2136 14424 2188 14476
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 2320 14399 2372 14408
rect 2320 14365 2329 14399
rect 2329 14365 2363 14399
rect 2363 14365 2372 14399
rect 2320 14356 2372 14365
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 1584 14220 1636 14272
rect 1952 14220 2004 14272
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 4214 14118 4266 14170
rect 4278 14118 4330 14170
rect 4342 14118 4394 14170
rect 4406 14118 4458 14170
rect 4470 14118 4522 14170
rect 7478 14118 7530 14170
rect 7542 14118 7594 14170
rect 7606 14118 7658 14170
rect 7670 14118 7722 14170
rect 7734 14118 7786 14170
rect 2228 13948 2280 14000
rect 1492 13880 1544 13932
rect 3608 13948 3660 14000
rect 9496 14016 9548 14068
rect 9588 14016 9640 14068
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 1768 13812 1820 13864
rect 1400 13719 1452 13728
rect 1400 13685 1409 13719
rect 1409 13685 1443 13719
rect 1443 13685 1452 13719
rect 1400 13676 1452 13685
rect 2412 13676 2464 13728
rect 2582 13574 2634 13626
rect 2646 13574 2698 13626
rect 2710 13574 2762 13626
rect 2774 13574 2826 13626
rect 2838 13574 2890 13626
rect 5846 13574 5898 13626
rect 5910 13574 5962 13626
rect 5974 13574 6026 13626
rect 6038 13574 6090 13626
rect 6102 13574 6154 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 9238 13574 9290 13626
rect 9302 13574 9354 13626
rect 9366 13574 9418 13626
rect 3056 13515 3108 13524
rect 2044 13404 2096 13456
rect 2504 13447 2556 13456
rect 2504 13413 2513 13447
rect 2513 13413 2547 13447
rect 2547 13413 2556 13447
rect 2504 13404 2556 13413
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 2228 13268 2280 13320
rect 3056 13481 3065 13515
rect 3065 13481 3099 13515
rect 3099 13481 3108 13515
rect 3056 13472 3108 13481
rect 9036 13472 9088 13524
rect 9864 13472 9916 13524
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 3884 13200 3936 13252
rect 1676 13132 1728 13184
rect 2412 13132 2464 13184
rect 3240 13132 3292 13184
rect 4214 13030 4266 13082
rect 4278 13030 4330 13082
rect 4342 13030 4394 13082
rect 4406 13030 4458 13082
rect 4470 13030 4522 13082
rect 7478 13030 7530 13082
rect 7542 13030 7594 13082
rect 7606 13030 7658 13082
rect 7670 13030 7722 13082
rect 7734 13030 7786 13082
rect 2320 12928 2372 12980
rect 3056 12928 3108 12980
rect 1400 12903 1452 12912
rect 1400 12869 1409 12903
rect 1409 12869 1443 12903
rect 1443 12869 1452 12903
rect 1400 12860 1452 12869
rect 1768 12860 1820 12912
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 3240 12792 3292 12844
rect 3792 12792 3844 12844
rect 9496 12724 9548 12776
rect 2964 12656 3016 12708
rect 3148 12656 3200 12708
rect 3700 12656 3752 12708
rect 3976 12656 4028 12708
rect 10048 12631 10100 12640
rect 10048 12597 10057 12631
rect 10057 12597 10091 12631
rect 10091 12597 10100 12631
rect 10048 12588 10100 12597
rect 2582 12486 2634 12538
rect 2646 12486 2698 12538
rect 2710 12486 2762 12538
rect 2774 12486 2826 12538
rect 2838 12486 2890 12538
rect 5846 12486 5898 12538
rect 5910 12486 5962 12538
rect 5974 12486 6026 12538
rect 6038 12486 6090 12538
rect 6102 12486 6154 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 9238 12486 9290 12538
rect 9302 12486 9354 12538
rect 9366 12486 9418 12538
rect 4712 12384 4764 12436
rect 3884 12248 3936 12300
rect 1216 12180 1268 12232
rect 2136 12180 2188 12232
rect 4620 12180 4672 12232
rect 4712 12180 4764 12232
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 4214 11942 4266 11994
rect 4278 11942 4330 11994
rect 4342 11942 4394 11994
rect 4406 11942 4458 11994
rect 4470 11942 4522 11994
rect 7478 11942 7530 11994
rect 7542 11942 7594 11994
rect 7606 11942 7658 11994
rect 7670 11942 7722 11994
rect 7734 11942 7786 11994
rect 3056 11883 3108 11892
rect 3056 11849 3065 11883
rect 3065 11849 3099 11883
rect 3099 11849 3108 11883
rect 3056 11840 3108 11849
rect 10140 11840 10192 11892
rect 3240 11772 3292 11824
rect 3056 11704 3108 11756
rect 3700 11747 3752 11756
rect 3700 11713 3709 11747
rect 3709 11713 3743 11747
rect 3743 11713 3752 11747
rect 3700 11704 3752 11713
rect 3884 11704 3936 11756
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 2964 11568 3016 11620
rect 3700 11500 3752 11552
rect 2582 11398 2634 11450
rect 2646 11398 2698 11450
rect 2710 11398 2762 11450
rect 2774 11398 2826 11450
rect 2838 11398 2890 11450
rect 5846 11398 5898 11450
rect 5910 11398 5962 11450
rect 5974 11398 6026 11450
rect 6038 11398 6090 11450
rect 6102 11398 6154 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 9238 11398 9290 11450
rect 9302 11398 9354 11450
rect 9366 11398 9418 11450
rect 3332 11296 3384 11348
rect 3424 11228 3476 11280
rect 10048 11271 10100 11280
rect 10048 11237 10057 11271
rect 10057 11237 10091 11271
rect 10091 11237 10100 11271
rect 10048 11228 10100 11237
rect 2136 11160 2188 11212
rect 1492 11092 1544 11144
rect 3056 11160 3108 11212
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 3332 11024 3384 11076
rect 4214 10854 4266 10906
rect 4278 10854 4330 10906
rect 4342 10854 4394 10906
rect 4406 10854 4458 10906
rect 4470 10854 4522 10906
rect 7478 10854 7530 10906
rect 7542 10854 7594 10906
rect 7606 10854 7658 10906
rect 7670 10854 7722 10906
rect 7734 10854 7786 10906
rect 9864 10752 9916 10804
rect 1952 10616 2004 10668
rect 3240 10616 3292 10668
rect 3516 10616 3568 10668
rect 4068 10616 4120 10668
rect 9864 10659 9916 10668
rect 9864 10625 9873 10659
rect 9873 10625 9907 10659
rect 9907 10625 9916 10659
rect 9864 10616 9916 10625
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 4896 10480 4948 10532
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 2582 10310 2634 10362
rect 2646 10310 2698 10362
rect 2710 10310 2762 10362
rect 2774 10310 2826 10362
rect 2838 10310 2890 10362
rect 5846 10310 5898 10362
rect 5910 10310 5962 10362
rect 5974 10310 6026 10362
rect 6038 10310 6090 10362
rect 6102 10310 6154 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 9238 10310 9290 10362
rect 9302 10310 9354 10362
rect 9366 10310 9418 10362
rect 3976 10251 4028 10260
rect 3976 10217 3985 10251
rect 3985 10217 4019 10251
rect 4019 10217 4028 10251
rect 3976 10208 4028 10217
rect 4712 10140 4764 10192
rect 1768 10072 1820 10124
rect 1492 10004 1544 10056
rect 3148 10004 3200 10056
rect 3976 10004 4028 10056
rect 4214 9766 4266 9818
rect 4278 9766 4330 9818
rect 4342 9766 4394 9818
rect 4406 9766 4458 9818
rect 4470 9766 4522 9818
rect 7478 9766 7530 9818
rect 7542 9766 7594 9818
rect 7606 9766 7658 9818
rect 7670 9766 7722 9818
rect 7734 9766 7786 9818
rect 3884 9596 3936 9648
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 3424 9528 3476 9580
rect 4712 9528 4764 9580
rect 3056 9392 3108 9444
rect 9864 9392 9916 9444
rect 10048 9435 10100 9444
rect 10048 9401 10057 9435
rect 10057 9401 10091 9435
rect 10091 9401 10100 9435
rect 10048 9392 10100 9401
rect 8300 9324 8352 9376
rect 2582 9222 2634 9274
rect 2646 9222 2698 9274
rect 2710 9222 2762 9274
rect 2774 9222 2826 9274
rect 2838 9222 2890 9274
rect 5846 9222 5898 9274
rect 5910 9222 5962 9274
rect 5974 9222 6026 9274
rect 6038 9222 6090 9274
rect 6102 9222 6154 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 9238 9222 9290 9274
rect 9302 9222 9354 9274
rect 9366 9222 9418 9274
rect 3056 9120 3108 9172
rect 3884 9120 3936 9172
rect 2044 8984 2096 9036
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 3056 8823 3108 8832
rect 3056 8789 3065 8823
rect 3065 8789 3099 8823
rect 3099 8789 3108 8823
rect 3056 8780 3108 8789
rect 10048 8823 10100 8832
rect 10048 8789 10057 8823
rect 10057 8789 10091 8823
rect 10091 8789 10100 8823
rect 10048 8780 10100 8789
rect 4214 8678 4266 8730
rect 4278 8678 4330 8730
rect 4342 8678 4394 8730
rect 4406 8678 4458 8730
rect 4470 8678 4522 8730
rect 7478 8678 7530 8730
rect 7542 8678 7594 8730
rect 7606 8678 7658 8730
rect 7670 8678 7722 8730
rect 7734 8678 7786 8730
rect 3608 8576 3660 8628
rect 2412 8440 2464 8492
rect 2964 8440 3016 8492
rect 3056 8440 3108 8492
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 2872 8304 2924 8356
rect 3056 8304 3108 8356
rect 10048 8347 10100 8356
rect 10048 8313 10057 8347
rect 10057 8313 10091 8347
rect 10091 8313 10100 8347
rect 10048 8304 10100 8313
rect 2582 8134 2634 8186
rect 2646 8134 2698 8186
rect 2710 8134 2762 8186
rect 2774 8134 2826 8186
rect 2838 8134 2890 8186
rect 5846 8134 5898 8186
rect 5910 8134 5962 8186
rect 5974 8134 6026 8186
rect 6038 8134 6090 8186
rect 6102 8134 6154 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 9238 8134 9290 8186
rect 9302 8134 9354 8186
rect 9366 8134 9418 8186
rect 5356 8032 5408 8084
rect 2228 7896 2280 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 1584 7828 1636 7880
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 3884 7828 3936 7880
rect 9864 7692 9916 7744
rect 4214 7590 4266 7642
rect 4278 7590 4330 7642
rect 4342 7590 4394 7642
rect 4406 7590 4458 7642
rect 4470 7590 4522 7642
rect 7478 7590 7530 7642
rect 7542 7590 7594 7642
rect 7606 7590 7658 7642
rect 7670 7590 7722 7642
rect 7734 7590 7786 7642
rect 3516 7488 3568 7540
rect 3792 7488 3844 7540
rect 2688 7420 2740 7472
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 2964 7284 3016 7336
rect 2412 7148 2464 7200
rect 9864 7148 9916 7200
rect 10048 7191 10100 7200
rect 10048 7157 10057 7191
rect 10057 7157 10091 7191
rect 10091 7157 10100 7191
rect 10048 7148 10100 7157
rect 2582 7046 2634 7098
rect 2646 7046 2698 7098
rect 2710 7046 2762 7098
rect 2774 7046 2826 7098
rect 2838 7046 2890 7098
rect 5846 7046 5898 7098
rect 5910 7046 5962 7098
rect 5974 7046 6026 7098
rect 6038 7046 6090 7098
rect 6102 7046 6154 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 9238 7046 9290 7098
rect 9302 7046 9354 7098
rect 9366 7046 9418 7098
rect 3148 6808 3200 6860
rect 4620 6808 4672 6860
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 2136 6740 2188 6792
rect 2504 6740 2556 6792
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 3148 6672 3200 6724
rect 1676 6604 1728 6656
rect 10048 6647 10100 6656
rect 10048 6613 10057 6647
rect 10057 6613 10091 6647
rect 10091 6613 10100 6647
rect 10048 6604 10100 6613
rect 4214 6502 4266 6554
rect 4278 6502 4330 6554
rect 4342 6502 4394 6554
rect 4406 6502 4458 6554
rect 4470 6502 4522 6554
rect 7478 6502 7530 6554
rect 7542 6502 7594 6554
rect 7606 6502 7658 6554
rect 7670 6502 7722 6554
rect 7734 6502 7786 6554
rect 1860 6443 1912 6452
rect 1860 6409 1869 6443
rect 1869 6409 1903 6443
rect 1903 6409 1912 6443
rect 1860 6400 1912 6409
rect 2596 6443 2648 6452
rect 2596 6409 2605 6443
rect 2605 6409 2639 6443
rect 2639 6409 2648 6443
rect 2596 6400 2648 6409
rect 3056 6332 3108 6384
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 9036 6060 9088 6112
rect 2582 5958 2634 6010
rect 2646 5958 2698 6010
rect 2710 5958 2762 6010
rect 2774 5958 2826 6010
rect 2838 5958 2890 6010
rect 5846 5958 5898 6010
rect 5910 5958 5962 6010
rect 5974 5958 6026 6010
rect 6038 5958 6090 6010
rect 6102 5958 6154 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 9238 5958 9290 6010
rect 9302 5958 9354 6010
rect 9366 5958 9418 6010
rect 2964 5856 3016 5908
rect 3976 5856 4028 5908
rect 3424 5720 3476 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 2228 5652 2280 5704
rect 4160 5652 4212 5704
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 4214 5414 4266 5466
rect 4278 5414 4330 5466
rect 4342 5414 4394 5466
rect 4406 5414 4458 5466
rect 4470 5414 4522 5466
rect 7478 5414 7530 5466
rect 7542 5414 7594 5466
rect 7606 5414 7658 5466
rect 7670 5414 7722 5466
rect 7734 5414 7786 5466
rect 2872 5355 2924 5364
rect 2872 5321 2881 5355
rect 2881 5321 2915 5355
rect 2915 5321 2924 5355
rect 2872 5312 2924 5321
rect 3240 5312 3292 5364
rect 1308 5176 1360 5228
rect 1952 5176 2004 5228
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 4528 5219 4580 5228
rect 4528 5185 4537 5219
rect 4537 5185 4571 5219
rect 4571 5185 4580 5219
rect 4528 5176 4580 5185
rect 9036 5176 9088 5228
rect 4712 5108 4764 5160
rect 9864 4972 9916 5024
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 2582 4870 2634 4922
rect 2646 4870 2698 4922
rect 2710 4870 2762 4922
rect 2774 4870 2826 4922
rect 2838 4870 2890 4922
rect 5846 4870 5898 4922
rect 5910 4870 5962 4922
rect 5974 4870 6026 4922
rect 6038 4870 6090 4922
rect 6102 4870 6154 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 9238 4870 9290 4922
rect 9302 4870 9354 4922
rect 9366 4870 9418 4922
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 4528 4768 4580 4820
rect 3700 4632 3752 4684
rect 3884 4632 3936 4684
rect 1860 4564 1912 4616
rect 2504 4607 2556 4616
rect 2504 4573 2513 4607
rect 2513 4573 2547 4607
rect 2547 4573 2556 4607
rect 2504 4564 2556 4573
rect 2780 4564 2832 4616
rect 3056 4564 3108 4616
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 9864 4607 9916 4616
rect 9864 4573 9873 4607
rect 9873 4573 9907 4607
rect 9907 4573 9916 4607
rect 9864 4564 9916 4573
rect 2320 4496 2372 4548
rect 2688 4496 2740 4548
rect 4160 4539 4212 4548
rect 4160 4505 4169 4539
rect 4169 4505 4203 4539
rect 4203 4505 4212 4539
rect 4160 4496 4212 4505
rect 9864 4428 9916 4480
rect 10048 4471 10100 4480
rect 10048 4437 10057 4471
rect 10057 4437 10091 4471
rect 10091 4437 10100 4471
rect 10048 4428 10100 4437
rect 4214 4326 4266 4378
rect 4278 4326 4330 4378
rect 4342 4326 4394 4378
rect 4406 4326 4458 4378
rect 4470 4326 4522 4378
rect 7478 4326 7530 4378
rect 7542 4326 7594 4378
rect 7606 4326 7658 4378
rect 7670 4326 7722 4378
rect 7734 4326 7786 4378
rect 4804 4224 4856 4276
rect 2412 4088 2464 4140
rect 2780 4131 2832 4140
rect 2780 4097 2789 4131
rect 2789 4097 2823 4131
rect 2823 4097 2832 4131
rect 2780 4088 2832 4097
rect 1768 4020 1820 4072
rect 2688 4020 2740 4072
rect 1216 3952 1268 4004
rect 2044 3884 2096 3936
rect 4620 3884 4672 3936
rect 5080 3927 5132 3936
rect 5080 3893 5089 3927
rect 5089 3893 5123 3927
rect 5123 3893 5132 3927
rect 5080 3884 5132 3893
rect 2582 3782 2634 3834
rect 2646 3782 2698 3834
rect 2710 3782 2762 3834
rect 2774 3782 2826 3834
rect 2838 3782 2890 3834
rect 5846 3782 5898 3834
rect 5910 3782 5962 3834
rect 5974 3782 6026 3834
rect 6038 3782 6090 3834
rect 6102 3782 6154 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 9238 3782 9290 3834
rect 9302 3782 9354 3834
rect 9366 3782 9418 3834
rect 2228 3680 2280 3732
rect 5540 3612 5592 3664
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 2412 3476 2464 3528
rect 4160 3476 4212 3528
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 9680 3408 9732 3460
rect 9864 3340 9916 3392
rect 10048 3383 10100 3392
rect 10048 3349 10057 3383
rect 10057 3349 10091 3383
rect 10091 3349 10100 3383
rect 10048 3340 10100 3349
rect 4214 3238 4266 3290
rect 4278 3238 4330 3290
rect 4342 3238 4394 3290
rect 4406 3238 4458 3290
rect 4470 3238 4522 3290
rect 7478 3238 7530 3290
rect 7542 3238 7594 3290
rect 7606 3238 7658 3290
rect 7670 3238 7722 3290
rect 7734 3238 7786 3290
rect 1676 3136 1728 3188
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 2504 3136 2556 3188
rect 3332 3179 3384 3188
rect 3332 3145 3341 3179
rect 3341 3145 3375 3179
rect 3375 3145 3384 3179
rect 3332 3136 3384 3145
rect 1400 3000 1452 3052
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 2964 3000 3016 3052
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 5080 3000 5132 3052
rect 9864 3043 9916 3052
rect 9864 3009 9873 3043
rect 9873 3009 9907 3043
rect 9907 3009 9916 3043
rect 9864 3000 9916 3009
rect 9496 2796 9548 2848
rect 10048 2839 10100 2848
rect 10048 2805 10057 2839
rect 10057 2805 10091 2839
rect 10091 2805 10100 2839
rect 10048 2796 10100 2805
rect 2582 2694 2634 2746
rect 2646 2694 2698 2746
rect 2710 2694 2762 2746
rect 2774 2694 2826 2746
rect 2838 2694 2890 2746
rect 5846 2694 5898 2746
rect 5910 2694 5962 2746
rect 5974 2694 6026 2746
rect 6038 2694 6090 2746
rect 6102 2694 6154 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 9238 2694 9290 2746
rect 9302 2694 9354 2746
rect 9366 2694 9418 2746
rect 2412 2592 2464 2644
rect 3884 2592 3936 2644
rect 2320 2524 2372 2576
rect 3976 2524 4028 2576
rect 1492 2388 1544 2440
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5540 2388 5592 2440
rect 9680 2388 9732 2440
rect 2780 2320 2832 2372
rect 1768 2252 1820 2304
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 9588 2252 9640 2304
rect 4214 2150 4266 2202
rect 4278 2150 4330 2202
rect 4342 2150 4394 2202
rect 4406 2150 4458 2202
rect 4470 2150 4522 2202
rect 7478 2150 7530 2202
rect 7542 2150 7594 2202
rect 7606 2150 7658 2202
rect 7670 2150 7722 2202
rect 7734 2150 7786 2202
rect 2872 1028 2924 1080
rect 4620 1028 4672 1080
<< metal2 >>
rect 1398 79248 1454 79257
rect 5998 79200 6054 80000
rect 9954 79520 10010 79529
rect 9954 79455 10010 79464
rect 1398 79183 1454 79192
rect 1306 78840 1362 78849
rect 1306 78775 1362 78784
rect 1320 77042 1348 78775
rect 1412 77586 1440 79183
rect 9586 78704 9642 78713
rect 9586 78639 9642 78648
rect 3882 78432 3938 78441
rect 3882 78367 3938 78376
rect 2582 77820 2890 77840
rect 2582 77818 2588 77820
rect 2644 77818 2668 77820
rect 2724 77818 2748 77820
rect 2804 77818 2828 77820
rect 2884 77818 2890 77820
rect 2644 77766 2646 77818
rect 2826 77766 2828 77818
rect 2582 77764 2588 77766
rect 2644 77764 2668 77766
rect 2724 77764 2748 77766
rect 2804 77764 2828 77766
rect 2884 77764 2890 77766
rect 2582 77744 2890 77764
rect 3606 77616 3662 77625
rect 1400 77580 1452 77586
rect 3606 77551 3662 77560
rect 3792 77580 3844 77586
rect 1400 77522 1452 77528
rect 1768 77512 1820 77518
rect 1768 77454 1820 77460
rect 2872 77512 2924 77518
rect 2872 77454 2924 77460
rect 1308 77036 1360 77042
rect 1308 76978 1360 76984
rect 1492 77036 1544 77042
rect 1492 76978 1544 76984
rect 1400 76832 1452 76838
rect 1400 76774 1452 76780
rect 1216 73704 1268 73710
rect 1216 73646 1268 73652
rect 664 72208 716 72214
rect 664 72150 716 72156
rect 572 69488 624 69494
rect 572 69430 624 69436
rect 204 66156 256 66162
rect 204 66098 256 66104
rect 20 62280 72 62286
rect 20 62222 72 62228
rect 32 46782 60 62222
rect 112 60036 164 60042
rect 112 59978 164 59984
rect 20 46776 72 46782
rect 20 46718 72 46724
rect 20 46368 72 46374
rect 20 46310 72 46316
rect 32 45914 60 46310
rect 124 46170 152 59978
rect 216 50454 244 66098
rect 480 65544 532 65550
rect 480 65486 532 65492
rect 492 59945 520 65486
rect 584 62336 612 69430
rect 676 65618 704 72150
rect 1228 72146 1256 73646
rect 1412 72842 1440 76774
rect 1504 75857 1532 76978
rect 1676 76084 1728 76090
rect 1676 76026 1728 76032
rect 1584 75948 1636 75954
rect 1584 75890 1636 75896
rect 1490 75848 1546 75857
rect 1490 75783 1546 75792
rect 1492 74724 1544 74730
rect 1492 74666 1544 74672
rect 1320 72814 1440 72842
rect 1216 72140 1268 72146
rect 1216 72082 1268 72088
rect 1320 71482 1348 72814
rect 1400 72684 1452 72690
rect 1400 72626 1452 72632
rect 1412 71641 1440 72626
rect 1504 72570 1532 74666
rect 1596 74633 1624 75890
rect 1582 74624 1638 74633
rect 1582 74559 1638 74568
rect 1584 73772 1636 73778
rect 1584 73714 1636 73720
rect 1596 72865 1624 73714
rect 1582 72856 1638 72865
rect 1582 72791 1638 72800
rect 1504 72542 1624 72570
rect 1492 72480 1544 72486
rect 1492 72422 1544 72428
rect 1398 71632 1454 71641
rect 1398 71567 1454 71576
rect 1320 71454 1440 71482
rect 940 70984 992 70990
rect 940 70926 992 70932
rect 952 70417 980 70926
rect 1124 70848 1176 70854
rect 1124 70790 1176 70796
rect 938 70408 994 70417
rect 938 70343 994 70352
rect 1136 69986 1164 70790
rect 1412 70666 1440 71454
rect 1504 70854 1532 72422
rect 1596 72185 1624 72542
rect 1582 72176 1638 72185
rect 1582 72111 1638 72120
rect 1584 72072 1636 72078
rect 1584 72014 1636 72020
rect 1596 71233 1624 72014
rect 1688 71670 1716 76026
rect 1676 71664 1728 71670
rect 1676 71606 1728 71612
rect 1676 71528 1728 71534
rect 1676 71470 1728 71476
rect 1582 71224 1638 71233
rect 1582 71159 1638 71168
rect 1688 71108 1716 71470
rect 1596 71080 1716 71108
rect 1492 70848 1544 70854
rect 1492 70790 1544 70796
rect 1320 70638 1440 70666
rect 1216 70440 1268 70446
rect 1216 70382 1268 70388
rect 1320 70394 1348 70638
rect 1596 70514 1624 71080
rect 1584 70508 1636 70514
rect 1584 70450 1636 70456
rect 1490 70408 1546 70417
rect 1044 69958 1164 69986
rect 940 67652 992 67658
rect 940 67594 992 67600
rect 848 66700 900 66706
rect 848 66642 900 66648
rect 664 65612 716 65618
rect 664 65554 716 65560
rect 584 62308 704 62336
rect 572 62212 624 62218
rect 572 62154 624 62160
rect 478 59936 534 59945
rect 478 59871 534 59880
rect 388 59628 440 59634
rect 388 59570 440 59576
rect 296 57452 348 57458
rect 296 57394 348 57400
rect 204 50448 256 50454
rect 204 50390 256 50396
rect 204 50312 256 50318
rect 204 50254 256 50260
rect 112 46164 164 46170
rect 112 46106 164 46112
rect 32 45886 152 45914
rect 18 45826 74 45835
rect 18 45761 74 45770
rect 32 26042 60 45761
rect 124 40458 152 45886
rect 112 40452 164 40458
rect 112 40394 164 40400
rect 110 39944 166 39953
rect 110 39879 166 39888
rect 124 39438 152 39879
rect 112 39432 164 39438
rect 112 39374 164 39380
rect 216 34134 244 50254
rect 204 34128 256 34134
rect 204 34070 256 34076
rect 308 33114 336 57394
rect 400 38418 428 59570
rect 480 59016 532 59022
rect 480 58958 532 58964
rect 492 38962 520 58958
rect 584 55962 612 62154
rect 676 56953 704 62308
rect 756 60104 808 60110
rect 756 60046 808 60052
rect 662 56944 718 56953
rect 662 56879 718 56888
rect 572 55956 624 55962
rect 572 55898 624 55904
rect 664 55752 716 55758
rect 664 55694 716 55700
rect 572 51468 624 51474
rect 572 51410 624 51416
rect 480 38956 532 38962
rect 480 38898 532 38904
rect 388 38412 440 38418
rect 388 38354 440 38360
rect 584 34610 612 51410
rect 676 46594 704 55694
rect 768 50386 796 60046
rect 860 56370 888 66642
rect 952 61606 980 67594
rect 1044 64394 1072 69958
rect 1124 65612 1176 65618
rect 1124 65554 1176 65560
rect 1032 64388 1084 64394
rect 1032 64330 1084 64336
rect 940 61600 992 61606
rect 940 61542 992 61548
rect 1032 61192 1084 61198
rect 1032 61134 1084 61140
rect 940 61124 992 61130
rect 940 61066 992 61072
rect 848 56364 900 56370
rect 848 56306 900 56312
rect 846 56094 902 56103
rect 846 56029 902 56038
rect 848 55956 900 55962
rect 848 55898 900 55904
rect 756 50380 808 50386
rect 756 50322 808 50328
rect 860 50266 888 55898
rect 768 50238 888 50266
rect 768 48210 796 50238
rect 952 50130 980 61066
rect 860 50102 980 50130
rect 860 48278 888 50102
rect 940 50040 992 50046
rect 940 49982 992 49988
rect 848 48272 900 48278
rect 848 48214 900 48220
rect 756 48204 808 48210
rect 756 48146 808 48152
rect 952 48142 980 49982
rect 940 48136 992 48142
rect 940 48078 992 48084
rect 756 48068 808 48074
rect 756 48010 808 48016
rect 768 46714 796 48010
rect 848 48000 900 48006
rect 848 47942 900 47948
rect 756 46708 808 46714
rect 756 46650 808 46656
rect 676 46566 796 46594
rect 664 46504 716 46510
rect 664 46446 716 46452
rect 676 41818 704 46446
rect 664 41812 716 41818
rect 664 41754 716 41760
rect 664 41676 716 41682
rect 664 41618 716 41624
rect 676 40118 704 41618
rect 768 41414 796 46566
rect 860 44402 888 47942
rect 1044 47138 1072 61134
rect 1136 60734 1164 65554
rect 1228 65550 1256 70382
rect 1320 70366 1440 70394
rect 1308 70100 1360 70106
rect 1308 70042 1360 70048
rect 1320 68746 1348 70042
rect 1412 70009 1440 70366
rect 1490 70343 1546 70352
rect 1398 70000 1454 70009
rect 1398 69935 1454 69944
rect 1400 69760 1452 69766
rect 1400 69702 1452 69708
rect 1412 69358 1440 69702
rect 1400 69352 1452 69358
rect 1400 69294 1452 69300
rect 1400 69216 1452 69222
rect 1400 69158 1452 69164
rect 1308 68740 1360 68746
rect 1308 68682 1360 68688
rect 1320 68406 1348 68682
rect 1308 68400 1360 68406
rect 1308 68342 1360 68348
rect 1320 67794 1348 68342
rect 1308 67788 1360 67794
rect 1308 67730 1360 67736
rect 1412 67266 1440 69158
rect 1504 68814 1532 70343
rect 1596 70106 1624 70450
rect 1780 70145 1808 77454
rect 2228 77376 2280 77382
rect 2228 77318 2280 77324
rect 1952 76560 2004 76566
rect 1952 76502 2004 76508
rect 1860 75540 1912 75546
rect 1860 75482 1912 75488
rect 1872 73030 1900 75482
rect 1964 74769 1992 76502
rect 2136 76492 2188 76498
rect 2136 76434 2188 76440
rect 2044 76424 2096 76430
rect 2044 76366 2096 76372
rect 2056 75886 2084 76366
rect 2148 76362 2176 76434
rect 2136 76356 2188 76362
rect 2136 76298 2188 76304
rect 2044 75880 2096 75886
rect 2044 75822 2096 75828
rect 2056 75206 2084 75822
rect 2148 75818 2176 76298
rect 2136 75812 2188 75818
rect 2136 75754 2188 75760
rect 2148 75274 2176 75754
rect 2240 75342 2268 77318
rect 2884 76945 2912 77454
rect 3056 77376 3108 77382
rect 3056 77318 3108 77324
rect 2964 77036 3016 77042
rect 2964 76978 3016 76984
rect 2870 76936 2926 76945
rect 2504 76900 2556 76906
rect 2870 76871 2926 76880
rect 2504 76842 2556 76848
rect 2320 76832 2372 76838
rect 2320 76774 2372 76780
rect 2228 75336 2280 75342
rect 2228 75278 2280 75284
rect 2136 75268 2188 75274
rect 2136 75210 2188 75216
rect 2044 75200 2096 75206
rect 2044 75142 2096 75148
rect 2056 74866 2084 75142
rect 2148 75002 2176 75210
rect 2136 74996 2188 75002
rect 2136 74938 2188 74944
rect 2044 74860 2096 74866
rect 2044 74802 2096 74808
rect 1950 74760 2006 74769
rect 1950 74695 2006 74704
rect 1952 74656 2004 74662
rect 1952 74598 2004 74604
rect 1860 73024 1912 73030
rect 1860 72966 1912 72972
rect 1860 71936 1912 71942
rect 1860 71878 1912 71884
rect 1872 70689 1900 71878
rect 1858 70680 1914 70689
rect 1858 70615 1914 70624
rect 1964 70394 1992 74598
rect 2056 74254 2084 74802
rect 2044 74248 2096 74254
rect 2044 74190 2096 74196
rect 2148 74186 2176 74938
rect 2136 74180 2188 74186
rect 2136 74122 2188 74128
rect 2044 73568 2096 73574
rect 2044 73510 2096 73516
rect 1872 70366 1992 70394
rect 1766 70136 1822 70145
rect 1584 70100 1636 70106
rect 1766 70071 1822 70080
rect 1584 70042 1636 70048
rect 1584 69896 1636 69902
rect 1582 69864 1584 69873
rect 1676 69896 1728 69902
rect 1636 69864 1638 69873
rect 1676 69838 1728 69844
rect 1582 69799 1638 69808
rect 1688 69465 1716 69838
rect 1768 69760 1820 69766
rect 1768 69702 1820 69708
rect 1674 69456 1730 69465
rect 1584 69420 1636 69426
rect 1674 69391 1730 69400
rect 1584 69362 1636 69368
rect 1492 68808 1544 68814
rect 1492 68750 1544 68756
rect 1492 68672 1544 68678
rect 1492 68614 1544 68620
rect 1504 67658 1532 68614
rect 1596 68241 1624 69362
rect 1676 69352 1728 69358
rect 1676 69294 1728 69300
rect 1582 68232 1638 68241
rect 1582 68167 1638 68176
rect 1584 67720 1636 67726
rect 1584 67662 1636 67668
rect 1492 67652 1544 67658
rect 1492 67594 1544 67600
rect 1596 67425 1624 67662
rect 1582 67416 1638 67425
rect 1582 67351 1638 67360
rect 1688 67266 1716 69294
rect 1412 67238 1532 67266
rect 1400 67176 1452 67182
rect 1400 67118 1452 67124
rect 1412 67017 1440 67118
rect 1398 67008 1454 67017
rect 1398 66943 1454 66952
rect 1400 66632 1452 66638
rect 1400 66574 1452 66580
rect 1412 66473 1440 66574
rect 1398 66464 1454 66473
rect 1398 66399 1454 66408
rect 1400 66088 1452 66094
rect 1306 66056 1362 66065
rect 1400 66030 1452 66036
rect 1306 65991 1362 66000
rect 1320 65618 1348 65991
rect 1412 65657 1440 66030
rect 1398 65648 1454 65657
rect 1308 65612 1360 65618
rect 1398 65583 1454 65592
rect 1308 65554 1360 65560
rect 1216 65544 1268 65550
rect 1216 65486 1268 65492
rect 1216 65204 1268 65210
rect 1216 65146 1268 65152
rect 1228 61402 1256 65146
rect 1398 65104 1454 65113
rect 1398 65039 1454 65048
rect 1412 63034 1440 65039
rect 1400 63028 1452 63034
rect 1400 62970 1452 62976
rect 1504 62880 1532 67238
rect 1596 67238 1716 67266
rect 1596 65113 1624 67238
rect 1676 67176 1728 67182
rect 1676 67118 1728 67124
rect 1688 66337 1716 67118
rect 1674 66328 1730 66337
rect 1674 66263 1730 66272
rect 1676 65544 1728 65550
rect 1676 65486 1728 65492
rect 1582 65104 1638 65113
rect 1582 65039 1638 65048
rect 1688 64977 1716 65486
rect 1674 64968 1730 64977
rect 1584 64932 1636 64938
rect 1674 64903 1730 64912
rect 1584 64874 1636 64880
rect 1596 63617 1624 64874
rect 1676 64864 1728 64870
rect 1676 64806 1728 64812
rect 1582 63608 1638 63617
rect 1582 63543 1638 63552
rect 1584 63300 1636 63306
rect 1584 63242 1636 63248
rect 1596 62898 1624 63242
rect 1320 62852 1532 62880
rect 1584 62892 1636 62898
rect 1216 61396 1268 61402
rect 1216 61338 1268 61344
rect 1136 60706 1256 60734
rect 1124 58336 1176 58342
rect 1124 58278 1176 58284
rect 1136 51542 1164 58278
rect 1228 56817 1256 60706
rect 1320 57916 1348 62852
rect 1584 62834 1636 62840
rect 1596 62762 1624 62834
rect 1400 62756 1452 62762
rect 1400 62698 1452 62704
rect 1584 62756 1636 62762
rect 1584 62698 1636 62704
rect 1412 61674 1440 62698
rect 1688 62665 1716 64806
rect 1674 62656 1730 62665
rect 1674 62591 1730 62600
rect 1584 62144 1636 62150
rect 1584 62086 1636 62092
rect 1400 61668 1452 61674
rect 1400 61610 1452 61616
rect 1412 60586 1440 61610
rect 1596 61441 1624 62086
rect 1780 61826 1808 69702
rect 1872 69494 1900 70366
rect 1950 70272 2006 70281
rect 1950 70207 2006 70216
rect 1860 69488 1912 69494
rect 1860 69430 1912 69436
rect 1860 69216 1912 69222
rect 1860 69158 1912 69164
rect 1688 61810 1808 61826
rect 1676 61804 1808 61810
rect 1728 61798 1808 61804
rect 1676 61746 1728 61752
rect 1676 61600 1728 61606
rect 1676 61542 1728 61548
rect 1582 61432 1638 61441
rect 1582 61367 1638 61376
rect 1584 61056 1636 61062
rect 1584 60998 1636 61004
rect 1400 60580 1452 60586
rect 1400 60522 1452 60528
rect 1412 60466 1440 60522
rect 1412 60438 1532 60466
rect 1400 59424 1452 59430
rect 1400 59366 1452 59372
rect 1412 58041 1440 59366
rect 1504 58614 1532 60438
rect 1596 60217 1624 60998
rect 1582 60208 1638 60217
rect 1582 60143 1638 60152
rect 1584 59968 1636 59974
rect 1584 59910 1636 59916
rect 1596 59265 1624 59910
rect 1582 59256 1638 59265
rect 1582 59191 1638 59200
rect 1584 58880 1636 58886
rect 1584 58822 1636 58828
rect 1492 58608 1544 58614
rect 1492 58550 1544 58556
rect 1398 58032 1454 58041
rect 1504 58002 1532 58550
rect 1398 57967 1454 57976
rect 1492 57996 1544 58002
rect 1492 57938 1544 57944
rect 1320 57888 1440 57916
rect 1308 57384 1360 57390
rect 1308 57326 1360 57332
rect 1214 56808 1270 56817
rect 1214 56743 1270 56752
rect 1216 56364 1268 56370
rect 1216 56306 1268 56312
rect 1124 51536 1176 51542
rect 1124 51478 1176 51484
rect 1124 51400 1176 51406
rect 1124 51342 1176 51348
rect 952 47110 1072 47138
rect 848 44396 900 44402
rect 848 44338 900 44344
rect 848 43716 900 43722
rect 848 43658 900 43664
rect 860 43330 888 43658
rect 952 43450 980 47110
rect 1030 46880 1086 46889
rect 1030 46815 1086 46824
rect 1044 46374 1072 46815
rect 1032 46368 1084 46374
rect 1032 46310 1084 46316
rect 1032 46164 1084 46170
rect 1032 46106 1084 46112
rect 940 43444 992 43450
rect 940 43386 992 43392
rect 860 43302 980 43330
rect 848 43172 900 43178
rect 848 43114 900 43120
rect 860 42702 888 43114
rect 848 42696 900 42702
rect 848 42638 900 42644
rect 860 41546 888 42638
rect 848 41540 900 41546
rect 848 41482 900 41488
rect 768 41386 888 41414
rect 756 41268 808 41274
rect 756 41210 808 41216
rect 664 40112 716 40118
rect 664 40054 716 40060
rect 662 39944 718 39953
rect 662 39879 718 39888
rect 572 34604 624 34610
rect 572 34546 624 34552
rect 572 34468 624 34474
rect 572 34410 624 34416
rect 296 33108 348 33114
rect 296 33050 348 33056
rect 584 31482 612 34410
rect 572 31476 624 31482
rect 572 31418 624 31424
rect 676 29306 704 39879
rect 768 32570 796 41210
rect 860 34202 888 41386
rect 952 36650 980 43302
rect 1044 40730 1072 46106
rect 1032 40724 1084 40730
rect 1032 40666 1084 40672
rect 1032 40044 1084 40050
rect 1032 39986 1084 39992
rect 1044 39098 1072 39986
rect 1032 39092 1084 39098
rect 1032 39034 1084 39040
rect 1032 37936 1084 37942
rect 1030 37904 1032 37913
rect 1084 37904 1086 37913
rect 1030 37839 1086 37848
rect 1032 37800 1084 37806
rect 1032 37742 1084 37748
rect 940 36644 992 36650
rect 940 36586 992 36592
rect 848 34196 900 34202
rect 848 34138 900 34144
rect 848 33992 900 33998
rect 848 33934 900 33940
rect 756 32564 808 32570
rect 756 32506 808 32512
rect 860 32366 888 33934
rect 1044 33386 1072 37742
rect 1032 33380 1084 33386
rect 1032 33322 1084 33328
rect 848 32360 900 32366
rect 848 32302 900 32308
rect 756 30728 808 30734
rect 756 30670 808 30676
rect 664 29300 716 29306
rect 664 29242 716 29248
rect 768 28082 796 30670
rect 756 28076 808 28082
rect 756 28018 808 28024
rect 768 27062 796 28018
rect 756 27056 808 27062
rect 756 26998 808 27004
rect 768 26450 796 26998
rect 756 26444 808 26450
rect 756 26386 808 26392
rect 20 26036 72 26042
rect 20 25978 72 25984
rect 768 23798 796 26386
rect 756 23792 808 23798
rect 756 23734 808 23740
rect 860 22094 888 32302
rect 940 31952 992 31958
rect 940 31894 992 31900
rect 952 31686 980 31894
rect 940 31680 992 31686
rect 940 31622 992 31628
rect 1032 31476 1084 31482
rect 1032 31418 1084 31424
rect 938 28792 994 28801
rect 938 28727 994 28736
rect 952 26382 980 28727
rect 1044 27606 1072 31418
rect 1032 27600 1084 27606
rect 1032 27542 1084 27548
rect 940 26376 992 26382
rect 940 26318 992 26324
rect 1136 24750 1164 51342
rect 1228 50998 1256 56306
rect 1320 51066 1348 57326
rect 1412 54754 1440 57888
rect 1492 57792 1544 57798
rect 1492 57734 1544 57740
rect 1504 57361 1532 57734
rect 1596 57633 1624 58822
rect 1688 57934 1716 61542
rect 1768 61396 1820 61402
rect 1768 61338 1820 61344
rect 1676 57928 1728 57934
rect 1676 57870 1728 57876
rect 1676 57792 1728 57798
rect 1676 57734 1728 57740
rect 1680 57718 1716 57734
rect 1582 57624 1638 57633
rect 1582 57559 1638 57568
rect 1680 57508 1708 57718
rect 1596 57497 1708 57508
rect 1582 57488 1708 57497
rect 1638 57480 1708 57488
rect 1780 57440 1808 61338
rect 1872 60654 1900 69158
rect 1964 68814 1992 70207
rect 1952 68808 2004 68814
rect 1952 68750 2004 68756
rect 2056 68474 2084 73510
rect 2148 73234 2176 74122
rect 2228 73772 2280 73778
rect 2228 73714 2280 73720
rect 2240 73273 2268 73714
rect 2226 73264 2282 73273
rect 2136 73228 2188 73234
rect 2226 73199 2282 73208
rect 2136 73170 2188 73176
rect 2148 72146 2176 73170
rect 2228 72684 2280 72690
rect 2228 72626 2280 72632
rect 2136 72140 2188 72146
rect 2136 72082 2188 72088
rect 2148 71670 2176 72082
rect 2240 72049 2268 72626
rect 2332 72078 2360 76774
rect 2516 76430 2544 76842
rect 2582 76732 2890 76752
rect 2582 76730 2588 76732
rect 2644 76730 2668 76732
rect 2724 76730 2748 76732
rect 2804 76730 2828 76732
rect 2884 76730 2890 76732
rect 2644 76678 2646 76730
rect 2826 76678 2828 76730
rect 2582 76676 2588 76678
rect 2644 76676 2668 76678
rect 2724 76676 2748 76678
rect 2804 76676 2828 76678
rect 2884 76676 2890 76678
rect 2582 76656 2890 76676
rect 2504 76424 2556 76430
rect 2504 76366 2556 76372
rect 2976 76265 3004 76978
rect 2962 76256 3018 76265
rect 2962 76191 3018 76200
rect 2596 76016 2648 76022
rect 3068 75970 3096 77318
rect 3620 77042 3648 77551
rect 3792 77522 3844 77528
rect 3608 77036 3660 77042
rect 3608 76978 3660 76984
rect 3148 76832 3200 76838
rect 3148 76774 3200 76780
rect 3424 76832 3476 76838
rect 3424 76774 3476 76780
rect 2648 75964 3096 75970
rect 2596 75958 3096 75964
rect 2504 75948 2556 75954
rect 2608 75942 3096 75958
rect 2504 75890 2556 75896
rect 2516 75818 2544 75890
rect 2504 75812 2556 75818
rect 2504 75754 2556 75760
rect 2582 75644 2890 75664
rect 2582 75642 2588 75644
rect 2644 75642 2668 75644
rect 2724 75642 2748 75644
rect 2804 75642 2828 75644
rect 2884 75642 2890 75644
rect 2644 75590 2646 75642
rect 2826 75590 2828 75642
rect 2582 75588 2588 75590
rect 2644 75588 2668 75590
rect 2724 75588 2748 75590
rect 2804 75588 2828 75590
rect 2884 75588 2890 75590
rect 2582 75568 2890 75588
rect 2504 75472 2556 75478
rect 2504 75414 2556 75420
rect 2412 74384 2464 74390
rect 2412 74326 2464 74332
rect 2320 72072 2372 72078
rect 2226 72040 2282 72049
rect 2320 72014 2372 72020
rect 2226 71975 2282 71984
rect 2228 71732 2280 71738
rect 2228 71674 2280 71680
rect 2136 71664 2188 71670
rect 2136 71606 2188 71612
rect 2240 71516 2268 71674
rect 2148 71488 2268 71516
rect 2148 70514 2176 71488
rect 2228 70984 2280 70990
rect 2228 70926 2280 70932
rect 2240 70825 2268 70926
rect 2320 70848 2372 70854
rect 2226 70816 2282 70825
rect 2320 70790 2372 70796
rect 2226 70751 2282 70760
rect 2136 70508 2188 70514
rect 2136 70450 2188 70456
rect 2332 70394 2360 70790
rect 2240 70366 2360 70394
rect 2240 69986 2268 70366
rect 2318 70272 2374 70281
rect 2318 70207 2374 70216
rect 2148 69958 2268 69986
rect 2044 68468 2096 68474
rect 2044 68410 2096 68416
rect 1952 68332 2004 68338
rect 1952 68274 2004 68280
rect 1964 62778 1992 68274
rect 2044 67856 2096 67862
rect 2044 67798 2096 67804
rect 2056 65210 2084 67798
rect 2044 65204 2096 65210
rect 2044 65146 2096 65152
rect 2044 65068 2096 65074
rect 2044 65010 2096 65016
rect 2056 62914 2084 65010
rect 2148 63356 2176 69958
rect 2228 69420 2280 69426
rect 2228 69362 2280 69368
rect 2240 69057 2268 69362
rect 2226 69048 2282 69057
rect 2226 68983 2282 68992
rect 2228 68808 2280 68814
rect 2228 68750 2280 68756
rect 2240 64002 2268 68750
rect 2332 64122 2360 70207
rect 2424 68338 2452 74326
rect 2516 72729 2544 75414
rect 2964 74860 3016 74866
rect 2964 74802 3016 74808
rect 2582 74556 2890 74576
rect 2582 74554 2588 74556
rect 2644 74554 2668 74556
rect 2724 74554 2748 74556
rect 2804 74554 2828 74556
rect 2884 74554 2890 74556
rect 2644 74502 2646 74554
rect 2826 74502 2828 74554
rect 2582 74500 2588 74502
rect 2644 74500 2668 74502
rect 2724 74500 2748 74502
rect 2804 74500 2828 74502
rect 2884 74500 2890 74502
rect 2582 74480 2890 74500
rect 2872 74248 2924 74254
rect 2872 74190 2924 74196
rect 2884 73658 2912 74190
rect 2976 73817 3004 74802
rect 3160 74186 3188 76774
rect 3436 76294 3464 76774
rect 3804 76650 3832 77522
rect 3896 77042 3924 78367
rect 4066 78024 4122 78033
rect 4066 77959 4122 77968
rect 9494 78024 9550 78033
rect 9494 77959 9550 77968
rect 4080 77518 4108 77959
rect 5846 77820 6154 77840
rect 5846 77818 5852 77820
rect 5908 77818 5932 77820
rect 5988 77818 6012 77820
rect 6068 77818 6092 77820
rect 6148 77818 6154 77820
rect 5908 77766 5910 77818
rect 6090 77766 6092 77818
rect 5846 77764 5852 77766
rect 5908 77764 5932 77766
rect 5988 77764 6012 77766
rect 6068 77764 6092 77766
rect 6148 77764 6154 77766
rect 5846 77744 6154 77764
rect 9110 77820 9418 77840
rect 9110 77818 9116 77820
rect 9172 77818 9196 77820
rect 9252 77818 9276 77820
rect 9332 77818 9356 77820
rect 9412 77818 9418 77820
rect 9172 77766 9174 77818
rect 9354 77766 9356 77818
rect 9110 77764 9116 77766
rect 9172 77764 9196 77766
rect 9252 77764 9276 77766
rect 9332 77764 9356 77766
rect 9412 77764 9418 77766
rect 9110 77744 9418 77764
rect 3976 77512 4028 77518
rect 3976 77454 4028 77460
rect 4068 77512 4120 77518
rect 4068 77454 4120 77460
rect 9404 77512 9456 77518
rect 9404 77454 9456 77460
rect 3988 77217 4016 77454
rect 4068 77376 4120 77382
rect 4068 77318 4120 77324
rect 8300 77376 8352 77382
rect 8300 77318 8352 77324
rect 3974 77208 4030 77217
rect 3974 77143 4030 77152
rect 3884 77036 3936 77042
rect 3884 76978 3936 76984
rect 4080 76922 4108 77318
rect 4214 77276 4522 77296
rect 4214 77274 4220 77276
rect 4276 77274 4300 77276
rect 4356 77274 4380 77276
rect 4436 77274 4460 77276
rect 4516 77274 4522 77276
rect 4276 77222 4278 77274
rect 4458 77222 4460 77274
rect 4214 77220 4220 77222
rect 4276 77220 4300 77222
rect 4356 77220 4380 77222
rect 4436 77220 4460 77222
rect 4516 77220 4522 77222
rect 4214 77200 4522 77220
rect 7478 77276 7786 77296
rect 7478 77274 7484 77276
rect 7540 77274 7564 77276
rect 7620 77274 7644 77276
rect 7700 77274 7724 77276
rect 7780 77274 7786 77276
rect 7540 77222 7542 77274
rect 7722 77222 7724 77274
rect 7478 77220 7484 77222
rect 7540 77220 7564 77222
rect 7620 77220 7644 77222
rect 7700 77220 7724 77222
rect 7780 77220 7786 77222
rect 7478 77200 7786 77220
rect 3988 76894 4108 76922
rect 3804 76622 3924 76650
rect 3792 76560 3844 76566
rect 3792 76502 3844 76508
rect 3424 76288 3476 76294
rect 3424 76230 3476 76236
rect 3516 76016 3568 76022
rect 3516 75958 3568 75964
rect 3424 75744 3476 75750
rect 3424 75686 3476 75692
rect 3240 75336 3292 75342
rect 3240 75278 3292 75284
rect 3252 75041 3280 75278
rect 3238 75032 3294 75041
rect 3238 74967 3294 74976
rect 3240 74248 3292 74254
rect 3238 74216 3240 74225
rect 3292 74216 3294 74225
rect 3148 74180 3200 74186
rect 3238 74151 3294 74160
rect 3148 74122 3200 74128
rect 3240 74112 3292 74118
rect 3240 74054 3292 74060
rect 2962 73808 3018 73817
rect 2962 73743 3018 73752
rect 2884 73630 3004 73658
rect 2582 73468 2890 73488
rect 2582 73466 2588 73468
rect 2644 73466 2668 73468
rect 2724 73466 2748 73468
rect 2804 73466 2828 73468
rect 2884 73466 2890 73468
rect 2644 73414 2646 73466
rect 2826 73414 2828 73466
rect 2582 73412 2588 73414
rect 2644 73412 2668 73414
rect 2724 73412 2748 73414
rect 2804 73412 2828 73414
rect 2884 73412 2890 73414
rect 2582 73392 2890 73412
rect 2976 73166 3004 73630
rect 3148 73636 3200 73642
rect 3148 73578 3200 73584
rect 2964 73160 3016 73166
rect 2964 73102 3016 73108
rect 2502 72720 2558 72729
rect 2502 72655 2558 72664
rect 2872 72684 2924 72690
rect 2872 72626 2924 72632
rect 2884 72593 2912 72626
rect 2870 72584 2926 72593
rect 2870 72519 2926 72528
rect 2504 72480 2556 72486
rect 2504 72422 2556 72428
rect 2412 68332 2464 68338
rect 2412 68274 2464 68280
rect 2412 68128 2464 68134
rect 2412 68070 2464 68076
rect 2320 64116 2372 64122
rect 2320 64058 2372 64064
rect 2240 63974 2360 64002
rect 2228 63912 2280 63918
rect 2228 63854 2280 63860
rect 2240 63510 2268 63854
rect 2228 63504 2280 63510
rect 2228 63446 2280 63452
rect 2228 63368 2280 63374
rect 2148 63328 2228 63356
rect 2228 63310 2280 63316
rect 2056 62886 2268 62914
rect 1964 62750 2176 62778
rect 1952 62688 2004 62694
rect 1952 62630 2004 62636
rect 1964 62490 1992 62630
rect 1952 62484 2004 62490
rect 1952 62426 2004 62432
rect 1952 62348 2004 62354
rect 1952 62290 2004 62296
rect 1964 61062 1992 62290
rect 2044 61600 2096 61606
rect 2044 61542 2096 61548
rect 1952 61056 2004 61062
rect 1952 60998 2004 61004
rect 1860 60648 1912 60654
rect 1860 60590 1912 60596
rect 1860 60512 1912 60518
rect 1860 60454 1912 60460
rect 1950 60480 2006 60489
rect 1872 57905 1900 60454
rect 1950 60415 2006 60424
rect 1858 57896 1914 57905
rect 1858 57831 1914 57840
rect 1860 57792 1912 57798
rect 1860 57734 1912 57740
rect 1582 57423 1638 57432
rect 1688 57412 1808 57440
rect 1490 57352 1546 57361
rect 1490 57287 1546 57296
rect 1492 57248 1544 57254
rect 1492 57190 1544 57196
rect 1504 57066 1532 57190
rect 1504 57038 1624 57066
rect 1492 56976 1544 56982
rect 1492 56918 1544 56924
rect 1504 54913 1532 56918
rect 1596 56681 1624 57038
rect 1582 56672 1638 56681
rect 1582 56607 1638 56616
rect 1688 56522 1716 57412
rect 1766 57080 1822 57089
rect 1766 57015 1822 57024
rect 1780 56710 1808 57015
rect 1768 56704 1820 56710
rect 1768 56646 1820 56652
rect 1596 56494 1716 56522
rect 1596 55214 1624 56494
rect 1780 55570 1808 56646
rect 1688 55542 1808 55570
rect 1688 55418 1716 55542
rect 1676 55412 1728 55418
rect 1676 55354 1728 55360
rect 1768 55412 1820 55418
rect 1768 55354 1820 55360
rect 1584 55208 1636 55214
rect 1584 55150 1636 55156
rect 1490 54904 1546 54913
rect 1490 54839 1546 54848
rect 1412 54726 1532 54754
rect 1504 54670 1532 54726
rect 1688 54720 1716 55354
rect 1596 54692 1716 54720
rect 1492 54664 1544 54670
rect 1492 54606 1544 54612
rect 1596 54602 1624 54692
rect 1584 54596 1636 54602
rect 1584 54538 1636 54544
rect 1400 53984 1452 53990
rect 1400 53926 1452 53932
rect 1412 53281 1440 53926
rect 1492 53576 1544 53582
rect 1492 53518 1544 53524
rect 1398 53272 1454 53281
rect 1398 53207 1454 53216
rect 1400 52896 1452 52902
rect 1400 52838 1452 52844
rect 1412 52057 1440 52838
rect 1504 52601 1532 53518
rect 1584 53440 1636 53446
rect 1584 53382 1636 53388
rect 1596 52873 1624 53382
rect 1582 52864 1638 52873
rect 1582 52799 1638 52808
rect 1490 52592 1546 52601
rect 1490 52527 1546 52536
rect 1492 52352 1544 52358
rect 1492 52294 1544 52300
rect 1398 52048 1454 52057
rect 1398 51983 1454 51992
rect 1504 51241 1532 52294
rect 1584 51808 1636 51814
rect 1584 51750 1636 51756
rect 1596 51649 1624 51750
rect 1582 51640 1638 51649
rect 1582 51575 1638 51584
rect 1584 51264 1636 51270
rect 1490 51232 1546 51241
rect 1584 51206 1636 51212
rect 1490 51167 1546 51176
rect 1596 51074 1624 51206
rect 1308 51060 1360 51066
rect 1308 51002 1360 51008
rect 1504 51046 1624 51074
rect 1216 50992 1268 50998
rect 1216 50934 1268 50940
rect 1306 50960 1362 50969
rect 1306 50895 1362 50904
rect 1320 50862 1348 50895
rect 1216 50856 1268 50862
rect 1216 50798 1268 50804
rect 1308 50856 1360 50862
rect 1308 50798 1360 50804
rect 1124 24744 1176 24750
rect 1124 24686 1176 24692
rect 1124 23656 1176 23662
rect 1122 23624 1124 23633
rect 1176 23624 1178 23633
rect 1122 23559 1178 23568
rect 1228 22094 1256 50798
rect 1308 50720 1360 50726
rect 1360 50668 1440 50674
rect 1308 50662 1440 50668
rect 1320 50646 1440 50662
rect 1308 50516 1360 50522
rect 1308 50458 1360 50464
rect 1320 48686 1348 50458
rect 1412 49473 1440 50646
rect 1504 50561 1532 51046
rect 1582 50960 1638 50969
rect 1582 50895 1638 50904
rect 1490 50552 1546 50561
rect 1490 50487 1546 50496
rect 1492 50312 1544 50318
rect 1492 50254 1544 50260
rect 1504 49842 1532 50254
rect 1492 49836 1544 49842
rect 1492 49778 1544 49784
rect 1398 49464 1454 49473
rect 1398 49399 1454 49408
rect 1504 49230 1532 49778
rect 1492 49224 1544 49230
rect 1492 49166 1544 49172
rect 1400 49088 1452 49094
rect 1400 49030 1452 49036
rect 1308 48680 1360 48686
rect 1308 48622 1360 48628
rect 1308 48544 1360 48550
rect 1308 48486 1360 48492
rect 1320 47977 1348 48486
rect 1306 47968 1362 47977
rect 1306 47903 1362 47912
rect 1412 47818 1440 49030
rect 1504 48754 1532 49166
rect 1492 48748 1544 48754
rect 1492 48690 1544 48696
rect 1492 48544 1544 48550
rect 1492 48486 1544 48492
rect 1320 47790 1440 47818
rect 1320 47444 1348 47790
rect 1400 47660 1452 47666
rect 1400 47602 1452 47608
rect 1412 47569 1440 47602
rect 1398 47560 1454 47569
rect 1398 47495 1454 47504
rect 1320 47416 1440 47444
rect 1308 45484 1360 45490
rect 1308 45426 1360 45432
rect 860 22066 1072 22094
rect 1044 21078 1072 22066
rect 1136 22066 1256 22094
rect 1032 21072 1084 21078
rect 1032 21014 1084 21020
rect 1136 17338 1164 22066
rect 1214 21448 1270 21457
rect 1214 21383 1270 21392
rect 1228 21010 1256 21383
rect 1216 21004 1268 21010
rect 1216 20946 1268 20952
rect 1214 19272 1270 19281
rect 1214 19207 1270 19216
rect 1228 18834 1256 19207
rect 1216 18828 1268 18834
rect 1216 18770 1268 18776
rect 1124 17332 1176 17338
rect 1124 17274 1176 17280
rect 1216 16584 1268 16590
rect 1216 16526 1268 16532
rect 1228 15065 1256 16526
rect 1214 15056 1270 15065
rect 1214 14991 1270 15000
rect 1216 12232 1268 12238
rect 1216 12174 1268 12180
rect 1228 11257 1256 12174
rect 1214 11248 1270 11257
rect 1214 11183 1270 11192
rect 1320 6914 1348 45426
rect 1412 41682 1440 47416
rect 1504 46034 1532 48486
rect 1596 48314 1624 50895
rect 1688 50561 1716 54692
rect 1780 51474 1808 55354
rect 1768 51468 1820 51474
rect 1768 51410 1820 51416
rect 1766 51368 1822 51377
rect 1766 51303 1822 51312
rect 1674 50552 1730 50561
rect 1674 50487 1730 50496
rect 1674 50416 1730 50425
rect 1674 50351 1730 50360
rect 1688 49910 1716 50351
rect 1780 50318 1808 51303
rect 1768 50312 1820 50318
rect 1768 50254 1820 50260
rect 1676 49904 1728 49910
rect 1676 49846 1728 49852
rect 1780 49842 1808 50254
rect 1768 49836 1820 49842
rect 1768 49778 1820 49784
rect 1674 49600 1730 49609
rect 1674 49535 1730 49544
rect 1688 49162 1716 49535
rect 1780 49230 1808 49778
rect 1768 49224 1820 49230
rect 1768 49166 1820 49172
rect 1676 49156 1728 49162
rect 1676 49098 1728 49104
rect 1674 48920 1730 48929
rect 1674 48855 1730 48864
rect 1688 48618 1716 48855
rect 1780 48754 1808 49166
rect 1768 48748 1820 48754
rect 1768 48690 1820 48696
rect 1676 48612 1728 48618
rect 1676 48554 1728 48560
rect 1766 48512 1822 48521
rect 1766 48447 1822 48456
rect 1596 48286 1716 48314
rect 1584 48000 1636 48006
rect 1584 47942 1636 47948
rect 1596 47841 1624 47942
rect 1582 47832 1638 47841
rect 1582 47767 1638 47776
rect 1584 47456 1636 47462
rect 1582 47424 1584 47433
rect 1636 47424 1638 47433
rect 1582 47359 1638 47368
rect 1584 47252 1636 47258
rect 1584 47194 1636 47200
rect 1492 46028 1544 46034
rect 1492 45970 1544 45976
rect 1596 45914 1624 47194
rect 1504 45886 1624 45914
rect 1504 45014 1532 45886
rect 1584 45824 1636 45830
rect 1584 45766 1636 45772
rect 1596 45529 1624 45766
rect 1582 45520 1638 45529
rect 1582 45455 1638 45464
rect 1584 45280 1636 45286
rect 1584 45222 1636 45228
rect 1492 45008 1544 45014
rect 1492 44950 1544 44956
rect 1492 44872 1544 44878
rect 1596 44849 1624 45222
rect 1492 44814 1544 44820
rect 1582 44840 1638 44849
rect 1504 43994 1532 44814
rect 1582 44775 1638 44784
rect 1584 44736 1636 44742
rect 1584 44678 1636 44684
rect 1492 43988 1544 43994
rect 1492 43930 1544 43936
rect 1492 43240 1544 43246
rect 1492 43182 1544 43188
rect 1504 42906 1532 43182
rect 1492 42900 1544 42906
rect 1492 42842 1544 42848
rect 1596 42786 1624 44678
rect 1504 42758 1624 42786
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1400 41540 1452 41546
rect 1400 41482 1452 41488
rect 1412 41138 1440 41482
rect 1504 41274 1532 42758
rect 1688 42634 1716 48286
rect 1780 47258 1808 48447
rect 1768 47252 1820 47258
rect 1768 47194 1820 47200
rect 1766 47152 1822 47161
rect 1766 47087 1822 47096
rect 1780 43382 1808 47087
rect 1768 43376 1820 43382
rect 1768 43318 1820 43324
rect 1676 42628 1728 42634
rect 1676 42570 1728 42576
rect 1674 42528 1730 42537
rect 1674 42463 1730 42472
rect 1584 42016 1636 42022
rect 1584 41958 1636 41964
rect 1492 41268 1544 41274
rect 1492 41210 1544 41216
rect 1490 41168 1546 41177
rect 1400 41132 1452 41138
rect 1490 41103 1546 41112
rect 1400 41074 1452 41080
rect 1412 40050 1440 41074
rect 1400 40044 1452 40050
rect 1400 39986 1452 39992
rect 1400 39296 1452 39302
rect 1400 39238 1452 39244
rect 1412 37641 1440 39238
rect 1504 38654 1532 41103
rect 1596 40633 1624 41958
rect 1688 41154 1716 42463
rect 1766 42392 1822 42401
rect 1766 42327 1822 42336
rect 1780 42226 1808 42327
rect 1768 42220 1820 42226
rect 1768 42162 1820 42168
rect 1768 41540 1820 41546
rect 1768 41482 1820 41488
rect 1780 41274 1808 41482
rect 1768 41268 1820 41274
rect 1768 41210 1820 41216
rect 1688 41126 1808 41154
rect 1674 40896 1730 40905
rect 1674 40831 1730 40840
rect 1582 40624 1638 40633
rect 1582 40559 1638 40568
rect 1584 40384 1636 40390
rect 1584 40326 1636 40332
rect 1596 38865 1624 40326
rect 1582 38856 1638 38865
rect 1582 38791 1638 38800
rect 1504 38626 1624 38654
rect 1492 38548 1544 38554
rect 1492 38490 1544 38496
rect 1504 38010 1532 38490
rect 1492 38004 1544 38010
rect 1492 37946 1544 37952
rect 1596 37890 1624 38626
rect 1504 37862 1624 37890
rect 1398 37632 1454 37641
rect 1398 37567 1454 37576
rect 1400 35556 1452 35562
rect 1400 35498 1452 35504
rect 1412 33674 1440 35498
rect 1504 35222 1532 37862
rect 1584 37664 1636 37670
rect 1584 37606 1636 37612
rect 1596 36718 1624 37606
rect 1584 36712 1636 36718
rect 1584 36654 1636 36660
rect 1584 35488 1636 35494
rect 1582 35456 1584 35465
rect 1636 35456 1638 35465
rect 1582 35391 1638 35400
rect 1492 35216 1544 35222
rect 1492 35158 1544 35164
rect 1688 35086 1716 40831
rect 1780 40769 1808 41126
rect 1766 40760 1822 40769
rect 1766 40695 1822 40704
rect 1768 40452 1820 40458
rect 1768 40394 1820 40400
rect 1676 35080 1728 35086
rect 1490 35048 1546 35057
rect 1676 35022 1728 35028
rect 1490 34983 1546 34992
rect 1504 34746 1532 34983
rect 1584 34944 1636 34950
rect 1584 34886 1636 34892
rect 1674 34912 1730 34921
rect 1492 34740 1544 34746
rect 1492 34682 1544 34688
rect 1596 34649 1624 34886
rect 1674 34847 1730 34856
rect 1582 34640 1638 34649
rect 1582 34575 1638 34584
rect 1412 33646 1532 33674
rect 1400 33584 1452 33590
rect 1400 33526 1452 33532
rect 1412 32337 1440 33526
rect 1398 32328 1454 32337
rect 1398 32263 1454 32272
rect 1504 32212 1532 33646
rect 1688 32978 1716 34847
rect 1676 32972 1728 32978
rect 1676 32914 1728 32920
rect 1780 32586 1808 40394
rect 1872 34610 1900 57734
rect 1964 55418 1992 60415
rect 1952 55412 2004 55418
rect 1952 55354 2004 55360
rect 1952 55072 2004 55078
rect 1952 55014 2004 55020
rect 1964 51241 1992 55014
rect 1950 51232 2006 51241
rect 1950 51167 2006 51176
rect 1950 50824 2006 50833
rect 1950 50759 1952 50768
rect 2004 50759 2006 50768
rect 1952 50730 2004 50736
rect 1950 50552 2006 50561
rect 1950 50487 2006 50496
rect 1964 50386 1992 50487
rect 1952 50380 2004 50386
rect 1952 50322 2004 50328
rect 1952 50176 2004 50182
rect 1952 50118 2004 50124
rect 1964 49745 1992 50118
rect 1950 49736 2006 49745
rect 1950 49671 2006 49680
rect 1952 49632 2004 49638
rect 1952 49574 2004 49580
rect 1964 47734 1992 49574
rect 1952 47728 2004 47734
rect 1952 47670 2004 47676
rect 1952 47592 2004 47598
rect 1952 47534 2004 47540
rect 1964 47258 1992 47534
rect 1952 47252 2004 47258
rect 1952 47194 2004 47200
rect 1952 46504 2004 46510
rect 1952 46446 2004 46452
rect 1964 46170 1992 46446
rect 1952 46164 2004 46170
rect 1952 46106 2004 46112
rect 1952 46028 2004 46034
rect 1952 45970 2004 45976
rect 1964 36378 1992 45970
rect 1952 36372 2004 36378
rect 1952 36314 2004 36320
rect 1952 36100 2004 36106
rect 1952 36042 2004 36048
rect 1860 34604 1912 34610
rect 1860 34546 1912 34552
rect 1860 34468 1912 34474
rect 1860 34410 1912 34416
rect 1872 33658 1900 34410
rect 1860 33652 1912 33658
rect 1964 33640 1992 36042
rect 2056 35086 2084 61542
rect 2148 61169 2176 62750
rect 2134 61160 2190 61169
rect 2134 61095 2190 61104
rect 2136 61056 2188 61062
rect 2136 60998 2188 61004
rect 2148 42226 2176 60998
rect 2240 52154 2268 62886
rect 2332 62354 2360 63974
rect 2424 63458 2452 68070
rect 2516 67726 2544 72422
rect 2582 72380 2890 72400
rect 2582 72378 2588 72380
rect 2644 72378 2668 72380
rect 2724 72378 2748 72380
rect 2804 72378 2828 72380
rect 2884 72378 2890 72380
rect 2644 72326 2646 72378
rect 2826 72326 2828 72378
rect 2582 72324 2588 72326
rect 2644 72324 2668 72326
rect 2724 72324 2748 72326
rect 2804 72324 2828 72326
rect 2884 72324 2890 72326
rect 2582 72304 2890 72324
rect 2872 72072 2924 72078
rect 2976 72060 3004 73102
rect 2924 72032 3004 72060
rect 2872 72014 2924 72020
rect 2884 71738 2912 72014
rect 2872 71732 2924 71738
rect 2872 71674 2924 71680
rect 2884 71602 2912 71674
rect 2872 71596 2924 71602
rect 2872 71538 2924 71544
rect 2964 71392 3016 71398
rect 2964 71334 3016 71340
rect 2582 71292 2890 71312
rect 2582 71290 2588 71292
rect 2644 71290 2668 71292
rect 2724 71290 2748 71292
rect 2804 71290 2828 71292
rect 2884 71290 2890 71292
rect 2644 71238 2646 71290
rect 2826 71238 2828 71290
rect 2582 71236 2588 71238
rect 2644 71236 2668 71238
rect 2724 71236 2748 71238
rect 2804 71236 2828 71238
rect 2884 71236 2890 71238
rect 2582 71216 2890 71236
rect 2688 71120 2740 71126
rect 2688 71062 2740 71068
rect 2700 70394 2728 71062
rect 2976 70922 3004 71334
rect 2964 70916 3016 70922
rect 2964 70858 3016 70864
rect 2700 70366 3004 70394
rect 2582 70204 2890 70224
rect 2582 70202 2588 70204
rect 2644 70202 2668 70204
rect 2724 70202 2748 70204
rect 2804 70202 2828 70204
rect 2884 70202 2890 70204
rect 2644 70150 2646 70202
rect 2826 70150 2828 70202
rect 2582 70148 2588 70150
rect 2644 70148 2668 70150
rect 2724 70148 2748 70150
rect 2804 70148 2828 70150
rect 2884 70148 2890 70150
rect 2582 70128 2890 70148
rect 2582 69116 2890 69136
rect 2582 69114 2588 69116
rect 2644 69114 2668 69116
rect 2724 69114 2748 69116
rect 2804 69114 2828 69116
rect 2884 69114 2890 69116
rect 2644 69062 2646 69114
rect 2826 69062 2828 69114
rect 2582 69060 2588 69062
rect 2644 69060 2668 69062
rect 2724 69060 2748 69062
rect 2804 69060 2828 69062
rect 2884 69060 2890 69062
rect 2582 69040 2890 69060
rect 2780 68808 2832 68814
rect 2780 68750 2832 68756
rect 2596 68740 2648 68746
rect 2596 68682 2648 68688
rect 2608 68406 2636 68682
rect 2792 68649 2820 68750
rect 2778 68640 2834 68649
rect 2778 68575 2834 68584
rect 2976 68490 3004 70366
rect 2976 68462 3096 68490
rect 2596 68400 2648 68406
rect 2596 68342 2648 68348
rect 2964 68332 3016 68338
rect 2964 68274 3016 68280
rect 2582 68028 2890 68048
rect 2582 68026 2588 68028
rect 2644 68026 2668 68028
rect 2724 68026 2748 68028
rect 2804 68026 2828 68028
rect 2884 68026 2890 68028
rect 2644 67974 2646 68026
rect 2826 67974 2828 68026
rect 2582 67972 2588 67974
rect 2644 67972 2668 67974
rect 2724 67972 2748 67974
rect 2804 67972 2828 67974
rect 2884 67972 2890 67974
rect 2582 67952 2890 67972
rect 2976 67833 3004 68274
rect 2962 67824 3018 67833
rect 2962 67759 3018 67768
rect 2504 67720 2556 67726
rect 2504 67662 2556 67668
rect 2778 67688 2834 67697
rect 2778 67623 2834 67632
rect 2872 67652 2924 67658
rect 2792 67250 2820 67623
rect 2872 67594 2924 67600
rect 2884 67318 2912 67594
rect 2872 67312 2924 67318
rect 2872 67254 2924 67260
rect 2780 67244 2832 67250
rect 2780 67186 2832 67192
rect 2884 67096 2912 67254
rect 2884 67068 3004 67096
rect 2582 66940 2890 66960
rect 2582 66938 2588 66940
rect 2644 66938 2668 66940
rect 2724 66938 2748 66940
rect 2804 66938 2828 66940
rect 2884 66938 2890 66940
rect 2644 66886 2646 66938
rect 2826 66886 2828 66938
rect 2582 66884 2588 66886
rect 2644 66884 2668 66886
rect 2724 66884 2748 66886
rect 2804 66884 2828 66886
rect 2884 66884 2890 66886
rect 2582 66864 2890 66884
rect 2976 66774 3004 67068
rect 2964 66768 3016 66774
rect 2884 66716 2964 66722
rect 2884 66710 3016 66716
rect 2884 66694 3004 66710
rect 2780 66632 2832 66638
rect 2780 66574 2832 66580
rect 2792 66065 2820 66574
rect 2884 66230 2912 66694
rect 2872 66224 2924 66230
rect 2872 66166 2924 66172
rect 2778 66056 2834 66065
rect 2778 65991 2834 66000
rect 2582 65852 2890 65872
rect 2582 65850 2588 65852
rect 2644 65850 2668 65852
rect 2724 65850 2748 65852
rect 2804 65850 2828 65852
rect 2884 65850 2890 65852
rect 2644 65798 2646 65850
rect 2826 65798 2828 65850
rect 2582 65796 2588 65798
rect 2644 65796 2668 65798
rect 2724 65796 2748 65798
rect 2804 65796 2828 65798
rect 2884 65796 2890 65798
rect 2582 65776 2890 65796
rect 2504 65544 2556 65550
rect 2504 65486 2556 65492
rect 2516 63889 2544 65486
rect 3068 65113 3096 68462
rect 3160 66298 3188 73578
rect 3252 70582 3280 74054
rect 3332 72548 3384 72554
rect 3332 72490 3384 72496
rect 3240 70576 3292 70582
rect 3240 70518 3292 70524
rect 3240 70440 3292 70446
rect 3240 70382 3292 70388
rect 3252 68406 3280 70382
rect 3240 68400 3292 68406
rect 3240 68342 3292 68348
rect 3252 67726 3280 68342
rect 3240 67720 3292 67726
rect 3344 67697 3372 72490
rect 3436 71670 3464 75686
rect 3424 71664 3476 71670
rect 3424 71606 3476 71612
rect 3240 67662 3292 67668
rect 3330 67688 3386 67697
rect 3252 67250 3280 67662
rect 3330 67623 3386 67632
rect 3240 67244 3292 67250
rect 3240 67186 3292 67192
rect 3148 66292 3200 66298
rect 3148 66234 3200 66240
rect 3252 66162 3280 67186
rect 3240 66156 3292 66162
rect 3240 66098 3292 66104
rect 3252 66042 3280 66098
rect 3160 66014 3280 66042
rect 3160 65618 3188 66014
rect 3240 65952 3292 65958
rect 3240 65894 3292 65900
rect 3148 65612 3200 65618
rect 3148 65554 3200 65560
rect 3054 65104 3110 65113
rect 3054 65039 3110 65048
rect 3148 65000 3200 65006
rect 3148 64942 3200 64948
rect 3056 64932 3108 64938
rect 3056 64874 3108 64880
rect 2582 64764 2890 64784
rect 2582 64762 2588 64764
rect 2644 64762 2668 64764
rect 2724 64762 2748 64764
rect 2804 64762 2828 64764
rect 2884 64762 2890 64764
rect 2644 64710 2646 64762
rect 2826 64710 2828 64762
rect 2582 64708 2588 64710
rect 2644 64708 2668 64710
rect 2724 64708 2748 64710
rect 2804 64708 2828 64710
rect 2884 64708 2890 64710
rect 2582 64688 2890 64708
rect 3068 64433 3096 64874
rect 3054 64424 3110 64433
rect 2964 64388 3016 64394
rect 3054 64359 3110 64368
rect 2964 64330 3016 64336
rect 2502 63880 2558 63889
rect 2502 63815 2558 63824
rect 2582 63676 2890 63696
rect 2582 63674 2588 63676
rect 2644 63674 2668 63676
rect 2724 63674 2748 63676
rect 2804 63674 2828 63676
rect 2884 63674 2890 63676
rect 2644 63622 2646 63674
rect 2826 63622 2828 63674
rect 2582 63620 2588 63622
rect 2644 63620 2668 63622
rect 2724 63620 2748 63622
rect 2804 63620 2828 63622
rect 2884 63620 2890 63622
rect 2582 63600 2890 63620
rect 2870 63472 2926 63481
rect 2424 63430 2544 63458
rect 2412 63368 2464 63374
rect 2412 63310 2464 63316
rect 2424 62898 2452 63310
rect 2412 62892 2464 62898
rect 2412 62834 2464 62840
rect 2424 62422 2452 62834
rect 2412 62416 2464 62422
rect 2412 62358 2464 62364
rect 2320 62348 2372 62354
rect 2320 62290 2372 62296
rect 2412 62280 2464 62286
rect 2412 62222 2464 62228
rect 2320 62144 2372 62150
rect 2320 62086 2372 62092
rect 2332 61849 2360 62086
rect 2318 61840 2374 61849
rect 2318 61775 2374 61784
rect 2320 61056 2372 61062
rect 2318 61024 2320 61033
rect 2372 61024 2374 61033
rect 2318 60959 2374 60968
rect 2318 60888 2374 60897
rect 2318 60823 2374 60832
rect 2332 60790 2360 60823
rect 2320 60784 2372 60790
rect 2320 60726 2372 60732
rect 2320 59968 2372 59974
rect 2320 59910 2372 59916
rect 2332 59673 2360 59910
rect 2318 59664 2374 59673
rect 2318 59599 2374 59608
rect 2320 58880 2372 58886
rect 2320 58822 2372 58828
rect 2332 58449 2360 58822
rect 2318 58440 2374 58449
rect 2318 58375 2374 58384
rect 2318 58304 2374 58313
rect 2318 58239 2374 58248
rect 2332 58070 2360 58239
rect 2320 58064 2372 58070
rect 2320 58006 2372 58012
rect 2424 57916 2452 62222
rect 2516 60296 2544 63430
rect 2870 63407 2926 63416
rect 2884 63374 2912 63407
rect 2872 63368 2924 63374
rect 2872 63310 2924 63316
rect 2688 63300 2740 63306
rect 2688 63242 2740 63248
rect 2596 62960 2648 62966
rect 2594 62928 2596 62937
rect 2648 62928 2650 62937
rect 2700 62898 2728 63242
rect 2884 62898 2912 63310
rect 2976 63306 3004 64330
rect 3056 64320 3108 64326
rect 3056 64262 3108 64268
rect 3068 63986 3096 64262
rect 3160 64025 3188 64942
rect 3146 64016 3202 64025
rect 3056 63980 3108 63986
rect 3146 63951 3202 63960
rect 3056 63922 3108 63928
rect 3068 63617 3096 63922
rect 3054 63608 3110 63617
rect 3054 63543 3110 63552
rect 3056 63504 3108 63510
rect 3056 63446 3108 63452
rect 3148 63504 3200 63510
rect 3148 63446 3200 63452
rect 2964 63300 3016 63306
rect 2964 63242 3016 63248
rect 2594 62863 2650 62872
rect 2688 62892 2740 62898
rect 2688 62834 2740 62840
rect 2872 62892 2924 62898
rect 2872 62834 2924 62840
rect 2582 62588 2890 62608
rect 2582 62586 2588 62588
rect 2644 62586 2668 62588
rect 2724 62586 2748 62588
rect 2804 62586 2828 62588
rect 2884 62586 2890 62588
rect 2644 62534 2646 62586
rect 2826 62534 2828 62586
rect 2582 62532 2588 62534
rect 2644 62532 2668 62534
rect 2724 62532 2748 62534
rect 2804 62532 2828 62534
rect 2884 62532 2890 62534
rect 2582 62512 2890 62532
rect 2596 62416 2648 62422
rect 2596 62358 2648 62364
rect 2608 61810 2636 62358
rect 2778 62248 2834 62257
rect 2778 62183 2834 62192
rect 2792 62150 2820 62183
rect 2780 62144 2832 62150
rect 2780 62086 2832 62092
rect 2596 61804 2648 61810
rect 2596 61746 2648 61752
rect 2608 61713 2636 61746
rect 2594 61704 2650 61713
rect 2594 61639 2650 61648
rect 2582 61500 2890 61520
rect 2582 61498 2588 61500
rect 2644 61498 2668 61500
rect 2724 61498 2748 61500
rect 2804 61498 2828 61500
rect 2884 61498 2890 61500
rect 2644 61446 2646 61498
rect 2826 61446 2828 61498
rect 2582 61444 2588 61446
rect 2644 61444 2668 61446
rect 2724 61444 2748 61446
rect 2804 61444 2828 61446
rect 2884 61444 2890 61446
rect 2582 61424 2890 61444
rect 2780 61056 2832 61062
rect 2780 60998 2832 61004
rect 2792 60858 2820 60998
rect 2780 60852 2832 60858
rect 2780 60794 2832 60800
rect 3068 60761 3096 63446
rect 3054 60752 3110 60761
rect 3054 60687 3056 60696
rect 3108 60687 3110 60696
rect 3056 60658 3108 60664
rect 2964 60648 3016 60654
rect 2778 60616 2834 60625
rect 2964 60590 3016 60596
rect 2778 60551 2780 60560
rect 2832 60551 2834 60560
rect 2780 60522 2832 60528
rect 2582 60412 2890 60432
rect 2582 60410 2588 60412
rect 2644 60410 2668 60412
rect 2724 60410 2748 60412
rect 2804 60410 2828 60412
rect 2884 60410 2890 60412
rect 2644 60358 2646 60410
rect 2826 60358 2828 60410
rect 2582 60356 2588 60358
rect 2644 60356 2668 60358
rect 2724 60356 2748 60358
rect 2804 60356 2828 60358
rect 2884 60356 2890 60358
rect 2582 60336 2890 60356
rect 2516 60268 2636 60296
rect 2502 60208 2558 60217
rect 2502 60143 2558 60152
rect 2332 57888 2452 57916
rect 2332 56817 2360 57888
rect 2410 57760 2466 57769
rect 2410 57695 2466 57704
rect 2424 57594 2452 57695
rect 2412 57588 2464 57594
rect 2412 57530 2464 57536
rect 2516 57322 2544 60143
rect 2608 60081 2636 60268
rect 2976 60246 3004 60590
rect 2964 60240 3016 60246
rect 2964 60182 3016 60188
rect 2964 60104 3016 60110
rect 2594 60072 2650 60081
rect 2964 60046 3016 60052
rect 2594 60007 2650 60016
rect 2582 59324 2890 59344
rect 2582 59322 2588 59324
rect 2644 59322 2668 59324
rect 2724 59322 2748 59324
rect 2804 59322 2828 59324
rect 2884 59322 2890 59324
rect 2644 59270 2646 59322
rect 2826 59270 2828 59322
rect 2582 59268 2588 59270
rect 2644 59268 2668 59270
rect 2724 59268 2748 59270
rect 2804 59268 2828 59270
rect 2884 59268 2890 59270
rect 2582 59248 2890 59268
rect 2686 59120 2742 59129
rect 2686 59055 2742 59064
rect 2700 58682 2728 59055
rect 2780 59016 2832 59022
rect 2780 58958 2832 58964
rect 2792 58682 2820 58958
rect 2688 58676 2740 58682
rect 2688 58618 2740 58624
rect 2780 58676 2832 58682
rect 2780 58618 2832 58624
rect 2688 58540 2740 58546
rect 2688 58482 2740 58488
rect 2700 58449 2728 58482
rect 2686 58440 2742 58449
rect 2686 58375 2742 58384
rect 2582 58236 2890 58256
rect 2582 58234 2588 58236
rect 2644 58234 2668 58236
rect 2724 58234 2748 58236
rect 2804 58234 2828 58236
rect 2884 58234 2890 58236
rect 2644 58182 2646 58234
rect 2826 58182 2828 58234
rect 2582 58180 2588 58182
rect 2644 58180 2668 58182
rect 2724 58180 2748 58182
rect 2804 58180 2828 58182
rect 2884 58180 2890 58182
rect 2582 58160 2890 58180
rect 2688 58064 2740 58070
rect 2594 58032 2650 58041
rect 2688 58006 2740 58012
rect 2778 58032 2834 58041
rect 2594 57967 2650 57976
rect 2608 57934 2636 57967
rect 2596 57928 2648 57934
rect 2596 57870 2648 57876
rect 2596 57792 2648 57798
rect 2596 57734 2648 57740
rect 2608 57361 2636 57734
rect 2700 57633 2728 58006
rect 2778 57967 2834 57976
rect 2792 57934 2820 57967
rect 2780 57928 2832 57934
rect 2780 57870 2832 57876
rect 2686 57624 2742 57633
rect 2686 57559 2742 57568
rect 2594 57352 2650 57361
rect 2504 57316 2556 57322
rect 2792 57322 2820 57870
rect 2594 57287 2650 57296
rect 2780 57316 2832 57322
rect 2504 57258 2556 57264
rect 2780 57258 2832 57264
rect 2412 57248 2464 57254
rect 2412 57190 2464 57196
rect 2318 56808 2374 56817
rect 2318 56743 2374 56752
rect 2320 56704 2372 56710
rect 2320 56646 2372 56652
rect 2332 55758 2360 56646
rect 2320 55752 2372 55758
rect 2320 55694 2372 55700
rect 2332 55321 2360 55694
rect 2318 55312 2374 55321
rect 2318 55247 2374 55256
rect 2320 55208 2372 55214
rect 2320 55150 2372 55156
rect 2332 54913 2360 55150
rect 2318 54904 2374 54913
rect 2318 54839 2374 54848
rect 2332 54670 2360 54839
rect 2320 54664 2372 54670
rect 2320 54606 2372 54612
rect 2320 54528 2372 54534
rect 2320 54470 2372 54476
rect 2332 54262 2360 54470
rect 2320 54256 2372 54262
rect 2320 54198 2372 54204
rect 2320 53984 2372 53990
rect 2320 53926 2372 53932
rect 2332 53825 2360 53926
rect 2318 53816 2374 53825
rect 2318 53751 2374 53760
rect 2318 53136 2374 53145
rect 2318 53071 2320 53080
rect 2372 53071 2374 53080
rect 2320 53042 2372 53048
rect 2320 52624 2372 52630
rect 2320 52566 2372 52572
rect 2332 52465 2360 52566
rect 2318 52456 2374 52465
rect 2318 52391 2374 52400
rect 2424 52193 2452 57190
rect 2582 57148 2890 57168
rect 2582 57146 2588 57148
rect 2644 57146 2668 57148
rect 2724 57146 2748 57148
rect 2804 57146 2828 57148
rect 2884 57146 2890 57148
rect 2644 57094 2646 57146
rect 2826 57094 2828 57146
rect 2582 57092 2588 57094
rect 2644 57092 2668 57094
rect 2724 57092 2748 57094
rect 2804 57092 2828 57094
rect 2884 57092 2890 57094
rect 2582 57072 2890 57092
rect 2976 57050 3004 60046
rect 3068 58970 3096 60658
rect 3160 60314 3188 63446
rect 3148 60308 3200 60314
rect 3148 60250 3200 60256
rect 3148 60172 3200 60178
rect 3148 60114 3200 60120
rect 3160 59129 3188 60114
rect 3146 59120 3202 59129
rect 3146 59055 3202 59064
rect 3068 58942 3188 58970
rect 3056 58880 3108 58886
rect 3054 58848 3056 58857
rect 3108 58848 3110 58857
rect 3054 58783 3110 58792
rect 3056 58676 3108 58682
rect 3056 58618 3108 58624
rect 3068 57769 3096 58618
rect 3054 57760 3110 57769
rect 3054 57695 3110 57704
rect 3160 57633 3188 58942
rect 3146 57624 3202 57633
rect 3146 57559 3202 57568
rect 3056 57452 3108 57458
rect 3056 57394 3108 57400
rect 3148 57452 3200 57458
rect 3148 57394 3200 57400
rect 3068 57361 3096 57394
rect 3054 57352 3110 57361
rect 3054 57287 3110 57296
rect 3056 57248 3108 57254
rect 3056 57190 3108 57196
rect 2964 57044 3016 57050
rect 2964 56986 3016 56992
rect 2502 56944 2558 56953
rect 2502 56879 2558 56888
rect 2596 56908 2648 56914
rect 2516 56778 2544 56879
rect 2596 56850 2648 56856
rect 2700 56902 2820 56930
rect 2504 56772 2556 56778
rect 2504 56714 2556 56720
rect 2502 56672 2558 56681
rect 2502 56607 2558 56616
rect 2516 55944 2544 56607
rect 2608 56545 2636 56850
rect 2700 56846 2728 56902
rect 2688 56840 2740 56846
rect 2792 56828 2820 56902
rect 2792 56800 2912 56828
rect 2688 56782 2740 56788
rect 2594 56536 2650 56545
rect 2594 56471 2650 56480
rect 2778 56536 2834 56545
rect 2778 56471 2834 56480
rect 2792 56438 2820 56471
rect 2780 56432 2832 56438
rect 2780 56374 2832 56380
rect 2884 56302 2912 56800
rect 2962 56400 3018 56409
rect 2962 56335 2964 56344
rect 3016 56335 3018 56344
rect 2964 56306 3016 56312
rect 2872 56296 2924 56302
rect 2872 56238 2924 56244
rect 2582 56060 2890 56080
rect 2582 56058 2588 56060
rect 2644 56058 2668 56060
rect 2724 56058 2748 56060
rect 2804 56058 2828 56060
rect 2884 56058 2890 56060
rect 2644 56006 2646 56058
rect 2826 56006 2828 56058
rect 2582 56004 2588 56006
rect 2644 56004 2668 56006
rect 2724 56004 2748 56006
rect 2804 56004 2828 56006
rect 2884 56004 2890 56006
rect 2582 55984 2890 56004
rect 2976 55944 3004 56306
rect 2516 55916 2636 55944
rect 2502 55720 2558 55729
rect 2502 55655 2558 55664
rect 2516 55282 2544 55655
rect 2504 55276 2556 55282
rect 2504 55218 2556 55224
rect 2608 55214 2636 55916
rect 2884 55916 3004 55944
rect 2596 55208 2648 55214
rect 2596 55150 2648 55156
rect 2884 55146 2912 55916
rect 3068 55865 3096 57190
rect 3160 55962 3188 57394
rect 3148 55956 3200 55962
rect 3148 55898 3200 55904
rect 3054 55856 3110 55865
rect 3054 55791 3110 55800
rect 3148 55616 3200 55622
rect 3054 55584 3110 55593
rect 3148 55558 3200 55564
rect 3054 55519 3110 55528
rect 2964 55208 3016 55214
rect 2964 55150 3016 55156
rect 2872 55140 2924 55146
rect 2872 55082 2924 55088
rect 2504 55072 2556 55078
rect 2504 55014 2556 55020
rect 2516 54641 2544 55014
rect 2582 54972 2890 54992
rect 2582 54970 2588 54972
rect 2644 54970 2668 54972
rect 2724 54970 2748 54972
rect 2804 54970 2828 54972
rect 2884 54970 2890 54972
rect 2644 54918 2646 54970
rect 2826 54918 2828 54970
rect 2582 54916 2588 54918
rect 2644 54916 2668 54918
rect 2724 54916 2748 54918
rect 2804 54916 2828 54918
rect 2884 54916 2890 54918
rect 2582 54896 2890 54916
rect 2502 54632 2558 54641
rect 2976 54618 3004 55150
rect 2502 54567 2558 54576
rect 2700 54590 3004 54618
rect 2700 54097 2728 54590
rect 2780 54528 2832 54534
rect 2780 54470 2832 54476
rect 2792 54233 2820 54470
rect 2962 54360 3018 54369
rect 3068 54330 3096 55519
rect 2962 54295 3018 54304
rect 3056 54324 3108 54330
rect 2778 54224 2834 54233
rect 2778 54159 2834 54168
rect 2686 54088 2742 54097
rect 2686 54023 2742 54032
rect 2582 53884 2890 53904
rect 2582 53882 2588 53884
rect 2644 53882 2668 53884
rect 2724 53882 2748 53884
rect 2804 53882 2828 53884
rect 2884 53882 2890 53884
rect 2644 53830 2646 53882
rect 2826 53830 2828 53882
rect 2582 53828 2588 53830
rect 2644 53828 2668 53830
rect 2724 53828 2748 53830
rect 2804 53828 2828 53830
rect 2884 53828 2890 53830
rect 2582 53808 2890 53828
rect 2976 53106 3004 54295
rect 3056 54266 3108 54272
rect 3056 54188 3108 54194
rect 3056 54130 3108 54136
rect 3068 53242 3096 54130
rect 3056 53236 3108 53242
rect 3056 53178 3108 53184
rect 2964 53100 3016 53106
rect 2964 53042 3016 53048
rect 2504 53032 2556 53038
rect 2504 52974 2556 52980
rect 2410 52184 2466 52193
rect 2228 52148 2280 52154
rect 2410 52119 2466 52128
rect 2228 52090 2280 52096
rect 2318 52048 2374 52057
rect 2228 52012 2280 52018
rect 2318 51983 2374 51992
rect 2412 52012 2464 52018
rect 2228 51954 2280 51960
rect 2240 49722 2268 51954
rect 2332 51474 2360 51983
rect 2412 51954 2464 51960
rect 2424 51610 2452 51954
rect 2516 51950 2544 52974
rect 2582 52796 2890 52816
rect 2582 52794 2588 52796
rect 2644 52794 2668 52796
rect 2724 52794 2748 52796
rect 2804 52794 2828 52796
rect 2884 52794 2890 52796
rect 2644 52742 2646 52794
rect 2826 52742 2828 52794
rect 2582 52740 2588 52742
rect 2644 52740 2668 52742
rect 2724 52740 2748 52742
rect 2804 52740 2828 52742
rect 2884 52740 2890 52742
rect 2582 52720 2890 52740
rect 2596 52420 2648 52426
rect 2596 52362 2648 52368
rect 2504 51944 2556 51950
rect 2502 51912 2504 51921
rect 2556 51912 2558 51921
rect 2502 51847 2558 51856
rect 2608 51796 2636 52362
rect 2976 52018 3004 53042
rect 3056 53032 3108 53038
rect 3056 52974 3108 52980
rect 2964 52012 3016 52018
rect 2964 51954 3016 51960
rect 2964 51876 3016 51882
rect 2964 51818 3016 51824
rect 2516 51768 2636 51796
rect 2412 51604 2464 51610
rect 2412 51546 2464 51552
rect 2320 51468 2372 51474
rect 2320 51410 2372 51416
rect 2412 51400 2464 51406
rect 2318 51368 2374 51377
rect 2412 51342 2464 51348
rect 2318 51303 2374 51312
rect 2332 50017 2360 51303
rect 2318 50008 2374 50017
rect 2318 49943 2374 49952
rect 2240 49694 2360 49722
rect 2228 49632 2280 49638
rect 2228 49574 2280 49580
rect 2240 48657 2268 49574
rect 2226 48648 2282 48657
rect 2332 48618 2360 49694
rect 2226 48583 2282 48592
rect 2320 48612 2372 48618
rect 2320 48554 2372 48560
rect 2424 48498 2452 51342
rect 2516 49366 2544 51768
rect 2582 51708 2890 51728
rect 2582 51706 2588 51708
rect 2644 51706 2668 51708
rect 2724 51706 2748 51708
rect 2804 51706 2828 51708
rect 2884 51706 2890 51708
rect 2644 51654 2646 51706
rect 2826 51654 2828 51706
rect 2582 51652 2588 51654
rect 2644 51652 2668 51654
rect 2724 51652 2748 51654
rect 2804 51652 2828 51654
rect 2884 51652 2890 51654
rect 2582 51632 2890 51652
rect 2976 51338 3004 51818
rect 3068 51513 3096 52974
rect 3054 51504 3110 51513
rect 3054 51439 3110 51448
rect 3056 51400 3108 51406
rect 3160 51377 3188 55558
rect 3252 53689 3280 65894
rect 3424 65068 3476 65074
rect 3424 65010 3476 65016
rect 3332 64864 3384 64870
rect 3330 64832 3332 64841
rect 3384 64832 3386 64841
rect 3330 64767 3386 64776
rect 3436 63510 3464 65010
rect 3424 63504 3476 63510
rect 3424 63446 3476 63452
rect 3424 63368 3476 63374
rect 3424 63310 3476 63316
rect 3332 63232 3384 63238
rect 3332 63174 3384 63180
rect 3344 63073 3372 63174
rect 3330 63064 3386 63073
rect 3330 62999 3386 63008
rect 3332 62960 3384 62966
rect 3332 62902 3384 62908
rect 3344 57594 3372 62902
rect 3332 57588 3384 57594
rect 3332 57530 3384 57536
rect 3332 57316 3384 57322
rect 3332 57258 3384 57264
rect 3344 56438 3372 57258
rect 3332 56432 3384 56438
rect 3332 56374 3384 56380
rect 3332 56228 3384 56234
rect 3332 56170 3384 56176
rect 3344 55894 3372 56170
rect 3332 55888 3384 55894
rect 3332 55830 3384 55836
rect 3332 55752 3384 55758
rect 3332 55694 3384 55700
rect 3238 53680 3294 53689
rect 3238 53615 3294 53624
rect 3344 53038 3372 55694
rect 3436 55622 3464 63310
rect 3424 55616 3476 55622
rect 3424 55558 3476 55564
rect 3424 55412 3476 55418
rect 3424 55354 3476 55360
rect 3436 55185 3464 55354
rect 3422 55176 3478 55185
rect 3422 55111 3478 55120
rect 3424 55072 3476 55078
rect 3424 55014 3476 55020
rect 3332 53032 3384 53038
rect 3332 52974 3384 52980
rect 3332 52012 3384 52018
rect 3332 51954 3384 51960
rect 3056 51342 3108 51348
rect 3146 51368 3202 51377
rect 2964 51332 3016 51338
rect 2964 51274 3016 51280
rect 2582 50620 2890 50640
rect 2582 50618 2588 50620
rect 2644 50618 2668 50620
rect 2724 50618 2748 50620
rect 2804 50618 2828 50620
rect 2884 50618 2890 50620
rect 2644 50566 2646 50618
rect 2826 50566 2828 50618
rect 2582 50564 2588 50566
rect 2644 50564 2668 50566
rect 2724 50564 2748 50566
rect 2804 50564 2828 50566
rect 2884 50564 2890 50566
rect 2582 50544 2890 50564
rect 2780 50176 2832 50182
rect 2780 50118 2832 50124
rect 2792 49881 2820 50118
rect 2778 49872 2834 49881
rect 2778 49807 2834 49816
rect 2582 49532 2890 49552
rect 2582 49530 2588 49532
rect 2644 49530 2668 49532
rect 2724 49530 2748 49532
rect 2804 49530 2828 49532
rect 2884 49530 2890 49532
rect 2644 49478 2646 49530
rect 2826 49478 2828 49530
rect 2582 49476 2588 49478
rect 2644 49476 2668 49478
rect 2724 49476 2748 49478
rect 2804 49476 2828 49478
rect 2884 49476 2890 49478
rect 2582 49456 2890 49476
rect 2504 49360 2556 49366
rect 2504 49302 2556 49308
rect 2780 49224 2832 49230
rect 2780 49166 2832 49172
rect 2688 49156 2740 49162
rect 2688 49098 2740 49104
rect 2700 48929 2728 49098
rect 2686 48920 2742 48929
rect 2686 48855 2742 48864
rect 2792 48657 2820 49166
rect 2872 49156 2924 49162
rect 2872 49098 2924 49104
rect 2884 48822 2912 49098
rect 2872 48816 2924 48822
rect 2872 48758 2924 48764
rect 2976 48770 3004 51274
rect 3068 49230 3096 51342
rect 3146 51303 3202 51312
rect 3344 50946 3372 51954
rect 3436 51218 3464 55014
rect 3528 53174 3556 75958
rect 3608 75948 3660 75954
rect 3608 75890 3660 75896
rect 3620 75449 3648 75890
rect 3606 75440 3662 75449
rect 3606 75375 3662 75384
rect 3608 70916 3660 70922
rect 3608 70858 3660 70864
rect 3516 53168 3568 53174
rect 3516 53110 3568 53116
rect 3436 51190 3556 51218
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3160 50918 3372 50946
rect 3056 49224 3108 49230
rect 3056 49166 3108 49172
rect 3054 48920 3110 48929
rect 3054 48855 3056 48864
rect 3108 48855 3110 48864
rect 3056 48826 3108 48832
rect 2976 48742 3096 48770
rect 3160 48754 3188 50918
rect 3238 50824 3294 50833
rect 3238 50759 3294 50768
rect 3252 49978 3280 50759
rect 3240 49972 3292 49978
rect 3240 49914 3292 49920
rect 3332 49700 3384 49706
rect 3332 49642 3384 49648
rect 3344 49434 3372 49642
rect 3332 49428 3384 49434
rect 3332 49370 3384 49376
rect 3240 49360 3292 49366
rect 3240 49302 3292 49308
rect 3330 49328 3386 49337
rect 2778 48648 2834 48657
rect 3068 48618 3096 48742
rect 3148 48748 3200 48754
rect 3148 48690 3200 48696
rect 2778 48583 2834 48592
rect 3056 48612 3108 48618
rect 3056 48554 3108 48560
rect 2240 48470 2452 48498
rect 2240 48346 2268 48470
rect 2582 48444 2890 48464
rect 2582 48442 2588 48444
rect 2644 48442 2668 48444
rect 2724 48442 2748 48444
rect 2804 48442 2828 48444
rect 2884 48442 2890 48444
rect 2644 48390 2646 48442
rect 2826 48390 2828 48442
rect 2582 48388 2588 48390
rect 2644 48388 2668 48390
rect 2724 48388 2748 48390
rect 2804 48388 2828 48390
rect 2884 48388 2890 48390
rect 2318 48376 2374 48385
rect 2228 48340 2280 48346
rect 2582 48368 2890 48388
rect 2962 48376 3018 48385
rect 2318 48311 2374 48320
rect 2962 48311 3018 48320
rect 2228 48282 2280 48288
rect 2332 48226 2360 48311
rect 2240 48198 2360 48226
rect 2504 48272 2556 48278
rect 2504 48214 2556 48220
rect 2136 42220 2188 42226
rect 2136 42162 2188 42168
rect 2136 42084 2188 42090
rect 2136 42026 2188 42032
rect 2148 40662 2176 42026
rect 2240 41313 2268 48198
rect 2412 48136 2464 48142
rect 2412 48078 2464 48084
rect 2320 47728 2372 47734
rect 2320 47670 2372 47676
rect 2332 46617 2360 47670
rect 2424 47258 2452 48078
rect 2412 47252 2464 47258
rect 2412 47194 2464 47200
rect 2516 47138 2544 48214
rect 2582 47356 2890 47376
rect 2582 47354 2588 47356
rect 2644 47354 2668 47356
rect 2724 47354 2748 47356
rect 2804 47354 2828 47356
rect 2884 47354 2890 47356
rect 2644 47302 2646 47354
rect 2826 47302 2828 47354
rect 2582 47300 2588 47302
rect 2644 47300 2668 47302
rect 2724 47300 2748 47302
rect 2804 47300 2828 47302
rect 2884 47300 2890 47302
rect 2582 47280 2890 47300
rect 2424 47110 2544 47138
rect 2688 47116 2740 47122
rect 2318 46608 2374 46617
rect 2318 46543 2374 46552
rect 2318 46472 2374 46481
rect 2318 46407 2374 46416
rect 2332 45626 2360 46407
rect 2320 45620 2372 45626
rect 2320 45562 2372 45568
rect 2318 45520 2374 45529
rect 2318 45455 2374 45464
rect 2332 44946 2360 45455
rect 2320 44940 2372 44946
rect 2320 44882 2372 44888
rect 2318 44840 2374 44849
rect 2318 44775 2374 44784
rect 2332 42158 2360 44775
rect 2320 42152 2372 42158
rect 2320 42094 2372 42100
rect 2320 42016 2372 42022
rect 2320 41958 2372 41964
rect 2332 41682 2360 41958
rect 2320 41676 2372 41682
rect 2424 41664 2452 47110
rect 2608 47076 2688 47104
rect 2504 47048 2556 47054
rect 2608 47036 2636 47076
rect 2688 47058 2740 47064
rect 2976 47054 3004 48311
rect 2556 47008 2636 47036
rect 2964 47048 3016 47054
rect 2504 46990 2556 46996
rect 2964 46990 3016 46996
rect 2516 46481 2544 46990
rect 2502 46472 2558 46481
rect 2502 46407 2558 46416
rect 2504 46368 2556 46374
rect 2504 46310 2556 46316
rect 2516 46073 2544 46310
rect 2582 46268 2890 46288
rect 2582 46266 2588 46268
rect 2644 46266 2668 46268
rect 2724 46266 2748 46268
rect 2804 46266 2828 46268
rect 2884 46266 2890 46268
rect 2644 46214 2646 46266
rect 2826 46214 2828 46266
rect 2582 46212 2588 46214
rect 2644 46212 2668 46214
rect 2724 46212 2748 46214
rect 2804 46212 2828 46214
rect 2884 46212 2890 46214
rect 2582 46192 2890 46212
rect 2502 46064 2558 46073
rect 2976 46034 3004 46990
rect 3056 46708 3108 46714
rect 3056 46650 3108 46656
rect 2502 45999 2558 46008
rect 2964 46028 3016 46034
rect 2964 45970 3016 45976
rect 2872 45960 2924 45966
rect 2502 45928 2558 45937
rect 2502 45863 2558 45872
rect 2870 45928 2872 45937
rect 2924 45928 2926 45937
rect 2870 45863 2926 45872
rect 2516 42129 2544 45863
rect 2870 45520 2926 45529
rect 2870 45455 2872 45464
rect 2924 45455 2926 45464
rect 2872 45426 2924 45432
rect 2594 45384 2650 45393
rect 2594 45319 2596 45328
rect 2648 45319 2650 45328
rect 2596 45290 2648 45296
rect 2976 45268 3004 45970
rect 3068 45966 3096 46650
rect 3056 45960 3108 45966
rect 3056 45902 3108 45908
rect 3056 45824 3108 45830
rect 3054 45792 3056 45801
rect 3108 45792 3110 45801
rect 3054 45727 3110 45736
rect 2976 45240 3096 45268
rect 2582 45180 2890 45200
rect 2582 45178 2588 45180
rect 2644 45178 2668 45180
rect 2724 45178 2748 45180
rect 2804 45178 2828 45180
rect 2884 45178 2890 45180
rect 2644 45126 2646 45178
rect 2826 45126 2828 45178
rect 2582 45124 2588 45126
rect 2644 45124 2668 45126
rect 2724 45124 2748 45126
rect 2804 45124 2828 45126
rect 2884 45124 2890 45126
rect 2582 45104 2890 45124
rect 2964 44736 3016 44742
rect 2962 44704 2964 44713
rect 3016 44704 3018 44713
rect 2962 44639 3018 44648
rect 2964 44532 3016 44538
rect 2964 44474 3016 44480
rect 2582 44092 2890 44112
rect 2582 44090 2588 44092
rect 2644 44090 2668 44092
rect 2724 44090 2748 44092
rect 2804 44090 2828 44092
rect 2884 44090 2890 44092
rect 2644 44038 2646 44090
rect 2826 44038 2828 44090
rect 2582 44036 2588 44038
rect 2644 44036 2668 44038
rect 2724 44036 2748 44038
rect 2804 44036 2828 44038
rect 2884 44036 2890 44038
rect 2582 44016 2890 44036
rect 2976 43976 3004 44474
rect 2884 43948 3004 43976
rect 2596 43784 2648 43790
rect 2596 43726 2648 43732
rect 2608 43178 2636 43726
rect 2596 43172 2648 43178
rect 2596 43114 2648 43120
rect 2884 43092 2912 43948
rect 3068 43790 3096 45240
rect 3160 44305 3188 48690
rect 3146 44296 3202 44305
rect 3146 44231 3202 44240
rect 3148 44192 3200 44198
rect 3148 44134 3200 44140
rect 3160 43897 3188 44134
rect 3146 43888 3202 43897
rect 3146 43823 3202 43832
rect 3056 43784 3108 43790
rect 3056 43726 3108 43732
rect 3148 43784 3200 43790
rect 3148 43726 3200 43732
rect 3054 43480 3110 43489
rect 3160 43450 3188 43726
rect 3054 43415 3110 43424
rect 3148 43444 3200 43450
rect 3068 43330 3096 43415
rect 3148 43386 3200 43392
rect 3068 43314 3188 43330
rect 2964 43308 3016 43314
rect 3068 43308 3200 43314
rect 3068 43302 3148 43308
rect 2964 43250 3016 43256
rect 3148 43250 3200 43256
rect 2976 43160 3004 43250
rect 2976 43132 3096 43160
rect 2884 43064 3004 43092
rect 2582 43004 2890 43024
rect 2582 43002 2588 43004
rect 2644 43002 2668 43004
rect 2724 43002 2748 43004
rect 2804 43002 2828 43004
rect 2884 43002 2890 43004
rect 2644 42950 2646 43002
rect 2826 42950 2828 43002
rect 2582 42948 2588 42950
rect 2644 42948 2668 42950
rect 2724 42948 2748 42950
rect 2804 42948 2828 42950
rect 2884 42948 2890 42950
rect 2582 42928 2890 42948
rect 2976 42945 3004 43064
rect 2962 42936 3018 42945
rect 2962 42871 3018 42880
rect 2870 42800 2926 42809
rect 2870 42735 2926 42744
rect 2780 42560 2832 42566
rect 2780 42502 2832 42508
rect 2792 42265 2820 42502
rect 2778 42256 2834 42265
rect 2884 42226 2912 42735
rect 2778 42191 2834 42200
rect 2872 42220 2924 42226
rect 2872 42162 2924 42168
rect 2502 42120 2558 42129
rect 3068 42106 3096 43132
rect 3148 42696 3200 42702
rect 3148 42638 3200 42644
rect 2502 42055 2558 42064
rect 2976 42078 3096 42106
rect 2582 41916 2890 41936
rect 2582 41914 2588 41916
rect 2644 41914 2668 41916
rect 2724 41914 2748 41916
rect 2804 41914 2828 41916
rect 2884 41914 2890 41916
rect 2644 41862 2646 41914
rect 2826 41862 2828 41914
rect 2582 41860 2588 41862
rect 2644 41860 2668 41862
rect 2724 41860 2748 41862
rect 2804 41860 2828 41862
rect 2884 41860 2890 41862
rect 2582 41840 2890 41860
rect 2872 41676 2924 41682
rect 2424 41636 2636 41664
rect 2320 41618 2372 41624
rect 2410 41576 2466 41585
rect 2410 41511 2466 41520
rect 2320 41472 2372 41478
rect 2318 41440 2320 41449
rect 2372 41440 2374 41449
rect 2318 41375 2374 41384
rect 2226 41304 2282 41313
rect 2424 41290 2452 41511
rect 2226 41239 2282 41248
rect 2332 41262 2452 41290
rect 2226 41168 2282 41177
rect 2226 41103 2282 41112
rect 2136 40656 2188 40662
rect 2136 40598 2188 40604
rect 2136 40520 2188 40526
rect 2136 40462 2188 40468
rect 2148 40186 2176 40462
rect 2136 40180 2188 40186
rect 2136 40122 2188 40128
rect 2134 40080 2190 40089
rect 2134 40015 2190 40024
rect 2148 35698 2176 40015
rect 2136 35692 2188 35698
rect 2136 35634 2188 35640
rect 2136 35556 2188 35562
rect 2136 35498 2188 35504
rect 2044 35080 2096 35086
rect 2044 35022 2096 35028
rect 2148 34474 2176 35498
rect 2240 34542 2268 41103
rect 2332 35034 2360 41262
rect 2608 41120 2636 41636
rect 2872 41618 2924 41624
rect 2688 41608 2740 41614
rect 2688 41550 2740 41556
rect 2700 41274 2728 41550
rect 2884 41274 2912 41618
rect 2688 41268 2740 41274
rect 2688 41210 2740 41216
rect 2872 41268 2924 41274
rect 2872 41210 2924 41216
rect 2780 41132 2832 41138
rect 2608 41092 2780 41120
rect 2780 41074 2832 41080
rect 2778 41032 2834 41041
rect 2778 40967 2780 40976
rect 2832 40967 2834 40976
rect 2780 40938 2832 40944
rect 2582 40828 2890 40848
rect 2582 40826 2588 40828
rect 2644 40826 2668 40828
rect 2724 40826 2748 40828
rect 2804 40826 2828 40828
rect 2884 40826 2890 40828
rect 2644 40774 2646 40826
rect 2826 40774 2828 40826
rect 2582 40772 2588 40774
rect 2644 40772 2668 40774
rect 2724 40772 2748 40774
rect 2804 40772 2828 40774
rect 2884 40772 2890 40774
rect 2582 40752 2890 40772
rect 2872 40656 2924 40662
rect 2872 40598 2924 40604
rect 2778 40080 2834 40089
rect 2412 40044 2464 40050
rect 2412 39986 2464 39992
rect 2504 40044 2556 40050
rect 2778 40015 2780 40024
rect 2504 39986 2556 39992
rect 2832 40015 2834 40024
rect 2780 39986 2832 39992
rect 2424 39284 2452 39986
rect 2516 39438 2544 39986
rect 2884 39953 2912 40598
rect 2976 40118 3004 42078
rect 3056 42016 3108 42022
rect 3056 41958 3108 41964
rect 3068 41721 3096 41958
rect 3054 41712 3110 41721
rect 3054 41647 3110 41656
rect 3056 41608 3108 41614
rect 3056 41550 3108 41556
rect 3068 41070 3096 41550
rect 3056 41064 3108 41070
rect 3054 41032 3056 41041
rect 3108 41032 3110 41041
rect 3054 40967 3110 40976
rect 3056 40928 3108 40934
rect 3056 40870 3108 40876
rect 2964 40112 3016 40118
rect 2964 40054 3016 40060
rect 2870 39944 2926 39953
rect 2870 39879 2872 39888
rect 2924 39879 2926 39888
rect 2872 39850 2924 39856
rect 2582 39740 2890 39760
rect 2582 39738 2588 39740
rect 2644 39738 2668 39740
rect 2724 39738 2748 39740
rect 2804 39738 2828 39740
rect 2884 39738 2890 39740
rect 2644 39686 2646 39738
rect 2826 39686 2828 39738
rect 2582 39684 2588 39686
rect 2644 39684 2668 39686
rect 2724 39684 2748 39686
rect 2804 39684 2828 39686
rect 2884 39684 2890 39686
rect 2582 39664 2890 39684
rect 2504 39432 2556 39438
rect 2504 39374 2556 39380
rect 2872 39432 2924 39438
rect 2872 39374 2924 39380
rect 2780 39364 2832 39370
rect 2780 39306 2832 39312
rect 2424 39256 2544 39284
rect 2412 39092 2464 39098
rect 2412 39034 2464 39040
rect 2424 38554 2452 39034
rect 2412 38548 2464 38554
rect 2412 38490 2464 38496
rect 2424 37398 2452 38490
rect 2412 37392 2464 37398
rect 2412 37334 2464 37340
rect 2412 37188 2464 37194
rect 2412 37130 2464 37136
rect 2424 36922 2452 37130
rect 2412 36916 2464 36922
rect 2412 36858 2464 36864
rect 2412 36712 2464 36718
rect 2412 36654 2464 36660
rect 2424 35562 2452 36654
rect 2412 35556 2464 35562
rect 2412 35498 2464 35504
rect 2332 35006 2452 35034
rect 2320 34944 2372 34950
rect 2320 34886 2372 34892
rect 2228 34536 2280 34542
rect 2228 34478 2280 34484
rect 2136 34468 2188 34474
rect 2136 34410 2188 34416
rect 2228 34400 2280 34406
rect 2228 34342 2280 34348
rect 2136 33924 2188 33930
rect 2136 33866 2188 33872
rect 2148 33658 2176 33866
rect 2136 33652 2188 33658
rect 1964 33612 2084 33640
rect 1860 33594 1912 33600
rect 1952 33516 2004 33522
rect 1872 33476 1952 33504
rect 1872 33386 1900 33476
rect 1952 33458 2004 33464
rect 1860 33380 1912 33386
rect 1860 33322 1912 33328
rect 1952 33380 2004 33386
rect 1952 33322 2004 33328
rect 1412 32184 1532 32212
rect 1688 32558 1808 32586
rect 1412 29646 1440 32184
rect 1582 32056 1638 32065
rect 1582 31991 1638 32000
rect 1492 31816 1544 31822
rect 1492 31758 1544 31764
rect 1504 30802 1532 31758
rect 1492 30796 1544 30802
rect 1492 30738 1544 30744
rect 1492 30660 1544 30666
rect 1492 30602 1544 30608
rect 1504 29889 1532 30602
rect 1490 29880 1546 29889
rect 1490 29815 1546 29824
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1492 29572 1544 29578
rect 1492 29514 1544 29520
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1412 27849 1440 29106
rect 1504 28257 1532 29514
rect 1490 28248 1546 28257
rect 1490 28183 1546 28192
rect 1490 28112 1546 28121
rect 1490 28047 1546 28056
rect 1398 27840 1454 27849
rect 1398 27775 1454 27784
rect 1400 27464 1452 27470
rect 1398 27432 1400 27441
rect 1452 27432 1454 27441
rect 1398 27367 1454 27376
rect 1504 27282 1532 28047
rect 1412 27254 1532 27282
rect 1412 23474 1440 27254
rect 1492 26376 1544 26382
rect 1492 26318 1544 26324
rect 1504 23610 1532 26318
rect 1596 23730 1624 31991
rect 1688 31958 1716 32558
rect 1872 32434 1900 33322
rect 1768 32428 1820 32434
rect 1768 32370 1820 32376
rect 1860 32428 1912 32434
rect 1860 32370 1912 32376
rect 1780 32026 1808 32370
rect 1768 32020 1820 32026
rect 1768 31962 1820 31968
rect 1676 31952 1728 31958
rect 1676 31894 1728 31900
rect 1872 31822 1900 32370
rect 1964 32201 1992 33322
rect 1950 32192 2006 32201
rect 1950 32127 2006 32136
rect 2056 31958 2084 33612
rect 2136 33594 2188 33600
rect 2240 33289 2268 34342
rect 2332 34241 2360 34886
rect 2318 34232 2374 34241
rect 2318 34167 2374 34176
rect 2424 33946 2452 35006
rect 2332 33918 2452 33946
rect 2226 33280 2282 33289
rect 2226 33215 2282 33224
rect 2332 32994 2360 33918
rect 2412 33856 2464 33862
rect 2412 33798 2464 33804
rect 2424 33590 2452 33798
rect 2412 33584 2464 33590
rect 2410 33552 2412 33561
rect 2464 33552 2466 33561
rect 2410 33487 2466 33496
rect 2412 33380 2464 33386
rect 2412 33322 2464 33328
rect 2148 32966 2360 32994
rect 2044 31952 2096 31958
rect 2044 31894 2096 31900
rect 1860 31816 1912 31822
rect 1860 31758 1912 31764
rect 2148 31754 2176 32966
rect 2320 32904 2372 32910
rect 2320 32846 2372 32852
rect 1676 31748 1728 31754
rect 1676 31690 1728 31696
rect 2136 31748 2188 31754
rect 2136 31690 2188 31696
rect 1688 26976 1716 31690
rect 1768 31680 1820 31686
rect 1768 31622 1820 31628
rect 1860 31680 1912 31686
rect 1860 31622 1912 31628
rect 1780 29102 1808 31622
rect 1872 30802 1900 31622
rect 2134 31376 2190 31385
rect 2044 31340 2096 31346
rect 2332 31346 2360 32846
rect 2424 32026 2452 33322
rect 2412 32020 2464 32026
rect 2412 31962 2464 31968
rect 2412 31816 2464 31822
rect 2412 31758 2464 31764
rect 2134 31311 2190 31320
rect 2320 31340 2372 31346
rect 2044 31282 2096 31288
rect 2056 30938 2084 31282
rect 2044 30932 2096 30938
rect 2044 30874 2096 30880
rect 1860 30796 1912 30802
rect 1860 30738 1912 30744
rect 2044 30796 2096 30802
rect 2044 30738 2096 30744
rect 1860 30252 1912 30258
rect 1860 30194 1912 30200
rect 1872 29481 1900 30194
rect 2056 30025 2084 30738
rect 2042 30016 2098 30025
rect 2042 29951 2098 29960
rect 2042 29880 2098 29889
rect 2042 29815 2098 29824
rect 2056 29782 2084 29815
rect 2044 29776 2096 29782
rect 2044 29718 2096 29724
rect 2044 29640 2096 29646
rect 2044 29582 2096 29588
rect 1858 29472 1914 29481
rect 1858 29407 1914 29416
rect 1858 29336 1914 29345
rect 1858 29271 1914 29280
rect 1768 29096 1820 29102
rect 1768 29038 1820 29044
rect 1872 28994 1900 29271
rect 1780 28966 1900 28994
rect 1780 28778 1808 28966
rect 1950 28928 2006 28937
rect 2056 28914 2084 29582
rect 2148 28937 2176 31311
rect 2320 31282 2372 31288
rect 2228 31136 2280 31142
rect 2228 31078 2280 31084
rect 2318 31104 2374 31113
rect 2006 28886 2084 28914
rect 2134 28928 2190 28937
rect 1950 28863 2006 28872
rect 2134 28863 2190 28872
rect 2240 28778 2268 31078
rect 2318 31039 2374 31048
rect 2332 28937 2360 31039
rect 2318 28928 2374 28937
rect 2318 28863 2374 28872
rect 2318 28792 2374 28801
rect 1780 28750 1900 28778
rect 2240 28750 2318 28778
rect 1768 28688 1820 28694
rect 1766 28656 1768 28665
rect 1820 28656 1822 28665
rect 1766 28591 1822 28600
rect 1768 28484 1820 28490
rect 1768 28426 1820 28432
rect 1780 28218 1808 28426
rect 1768 28212 1820 28218
rect 1768 28154 1820 28160
rect 1688 26948 1808 26976
rect 1674 26888 1730 26897
rect 1674 26823 1676 26832
rect 1728 26823 1730 26832
rect 1676 26794 1728 26800
rect 1676 26512 1728 26518
rect 1676 26454 1728 26460
rect 1584 23724 1636 23730
rect 1584 23666 1636 23672
rect 1504 23582 1624 23610
rect 1412 23446 1532 23474
rect 1400 23112 1452 23118
rect 1398 23080 1400 23089
rect 1452 23080 1454 23089
rect 1398 23015 1454 23024
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1412 21865 1440 21966
rect 1398 21856 1454 21865
rect 1398 21791 1454 21800
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 21049 1440 21422
rect 1398 21040 1454 21049
rect 1398 20975 1454 20984
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1412 20233 1440 20334
rect 1398 20224 1454 20233
rect 1398 20159 1454 20168
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1412 19689 1440 19790
rect 1398 19680 1454 19689
rect 1398 19615 1454 19624
rect 1504 19378 1532 23446
rect 1596 19922 1624 23582
rect 1688 20466 1716 26454
rect 1780 23882 1808 26948
rect 1872 25498 1900 28750
rect 2318 28727 2374 28736
rect 2424 28676 2452 31758
rect 2516 31754 2544 39256
rect 2792 38826 2820 39306
rect 2884 38865 2912 39374
rect 2976 38876 3004 40054
rect 3068 39506 3096 40870
rect 3056 39500 3108 39506
rect 3056 39442 3108 39448
rect 3056 39364 3108 39370
rect 3056 39306 3108 39312
rect 3068 39001 3096 39306
rect 3054 38992 3110 39001
rect 3054 38927 3110 38936
rect 2870 38856 2926 38865
rect 2780 38820 2832 38826
rect 2976 38848 3096 38876
rect 2870 38791 2926 38800
rect 2780 38762 2832 38768
rect 2964 38752 3016 38758
rect 2964 38694 3016 38700
rect 2582 38652 2890 38672
rect 2582 38650 2588 38652
rect 2644 38650 2668 38652
rect 2724 38650 2748 38652
rect 2804 38650 2828 38652
rect 2884 38650 2890 38652
rect 2644 38598 2646 38650
rect 2826 38598 2828 38650
rect 2582 38596 2588 38598
rect 2644 38596 2668 38598
rect 2724 38596 2748 38598
rect 2804 38596 2828 38598
rect 2884 38596 2890 38598
rect 2582 38576 2890 38596
rect 2778 38312 2834 38321
rect 2688 38276 2740 38282
rect 2778 38247 2834 38256
rect 2688 38218 2740 38224
rect 2594 38176 2650 38185
rect 2594 38111 2650 38120
rect 2608 37874 2636 38111
rect 2700 38010 2728 38218
rect 2688 38004 2740 38010
rect 2688 37946 2740 37952
rect 2792 37942 2820 38247
rect 2976 38049 3004 38694
rect 2962 38040 3018 38049
rect 2962 37975 3018 37984
rect 2780 37936 2832 37942
rect 2780 37878 2832 37884
rect 2596 37868 2648 37874
rect 2596 37810 2648 37816
rect 2964 37868 3016 37874
rect 2964 37810 3016 37816
rect 2582 37564 2890 37584
rect 2582 37562 2588 37564
rect 2644 37562 2668 37564
rect 2724 37562 2748 37564
rect 2804 37562 2828 37564
rect 2884 37562 2890 37564
rect 2644 37510 2646 37562
rect 2826 37510 2828 37562
rect 2582 37508 2588 37510
rect 2644 37508 2668 37510
rect 2724 37508 2748 37510
rect 2804 37508 2828 37510
rect 2884 37508 2890 37510
rect 2582 37488 2890 37508
rect 2686 37360 2742 37369
rect 2686 37295 2742 37304
rect 2596 37256 2648 37262
rect 2596 37198 2648 37204
rect 2608 36786 2636 37198
rect 2700 37126 2728 37295
rect 2976 37262 3004 37810
rect 2964 37256 3016 37262
rect 2964 37198 3016 37204
rect 2688 37120 2740 37126
rect 2688 37062 2740 37068
rect 2596 36780 2648 36786
rect 2596 36722 2648 36728
rect 2582 36476 2890 36496
rect 2582 36474 2588 36476
rect 2644 36474 2668 36476
rect 2724 36474 2748 36476
rect 2804 36474 2828 36476
rect 2884 36474 2890 36476
rect 2644 36422 2646 36474
rect 2826 36422 2828 36474
rect 2582 36420 2588 36422
rect 2644 36420 2668 36422
rect 2724 36420 2748 36422
rect 2804 36420 2828 36422
rect 2884 36420 2890 36422
rect 2582 36400 2890 36420
rect 2780 36032 2832 36038
rect 2780 35974 2832 35980
rect 2792 35873 2820 35974
rect 2778 35864 2834 35873
rect 2778 35799 2834 35808
rect 2964 35692 3016 35698
rect 3068 35680 3096 38848
rect 3160 36786 3188 42638
rect 3148 36780 3200 36786
rect 3148 36722 3200 36728
rect 3016 35652 3096 35680
rect 2964 35634 3016 35640
rect 2582 35388 2890 35408
rect 2582 35386 2588 35388
rect 2644 35386 2668 35388
rect 2724 35386 2748 35388
rect 2804 35386 2828 35388
rect 2884 35386 2890 35388
rect 2644 35334 2646 35386
rect 2826 35334 2828 35386
rect 2582 35332 2588 35334
rect 2644 35332 2668 35334
rect 2724 35332 2748 35334
rect 2804 35332 2828 35334
rect 2884 35332 2890 35334
rect 2582 35312 2890 35332
rect 2596 35216 2648 35222
rect 2596 35158 2648 35164
rect 2608 34610 2636 35158
rect 2596 34604 2648 34610
rect 2596 34546 2648 34552
rect 2582 34300 2890 34320
rect 2582 34298 2588 34300
rect 2644 34298 2668 34300
rect 2724 34298 2748 34300
rect 2804 34298 2828 34300
rect 2884 34298 2890 34300
rect 2644 34246 2646 34298
rect 2826 34246 2828 34298
rect 2582 34244 2588 34246
rect 2644 34244 2668 34246
rect 2724 34244 2748 34246
rect 2804 34244 2828 34246
rect 2884 34244 2890 34246
rect 2582 34224 2890 34244
rect 2976 34184 3004 35634
rect 3148 35080 3200 35086
rect 3148 35022 3200 35028
rect 3056 34400 3108 34406
rect 3056 34342 3108 34348
rect 2884 34156 3004 34184
rect 2884 33300 2912 34156
rect 2964 33924 3016 33930
rect 2964 33866 3016 33872
rect 2976 33658 3004 33866
rect 3068 33833 3096 34342
rect 3054 33824 3110 33833
rect 3054 33759 3110 33768
rect 2964 33652 3016 33658
rect 2964 33594 3016 33600
rect 3054 33552 3110 33561
rect 3054 33487 3110 33496
rect 2964 33312 3016 33318
rect 2884 33272 2964 33300
rect 2964 33254 3016 33260
rect 2582 33212 2890 33232
rect 2582 33210 2588 33212
rect 2644 33210 2668 33212
rect 2724 33210 2748 33212
rect 2804 33210 2828 33212
rect 2884 33210 2890 33212
rect 2644 33158 2646 33210
rect 2826 33158 2828 33210
rect 2582 33156 2588 33158
rect 2644 33156 2668 33158
rect 2724 33156 2748 33158
rect 2804 33156 2828 33158
rect 2884 33156 2890 33158
rect 2582 33136 2890 33156
rect 2976 32910 3004 33254
rect 2964 32904 3016 32910
rect 2964 32846 3016 32852
rect 2596 32836 2648 32842
rect 2596 32778 2648 32784
rect 2608 32570 2636 32778
rect 2596 32564 2648 32570
rect 2596 32506 2648 32512
rect 2582 32124 2890 32144
rect 2582 32122 2588 32124
rect 2644 32122 2668 32124
rect 2724 32122 2748 32124
rect 2804 32122 2828 32124
rect 2884 32122 2890 32124
rect 2644 32070 2646 32122
rect 2826 32070 2828 32122
rect 2582 32068 2588 32070
rect 2644 32068 2668 32070
rect 2724 32068 2748 32070
rect 2804 32068 2828 32070
rect 2884 32068 2890 32070
rect 2582 32048 2890 32068
rect 2688 31952 2740 31958
rect 2688 31894 2740 31900
rect 2516 31726 2636 31754
rect 2608 31346 2636 31726
rect 2596 31340 2648 31346
rect 2596 31282 2648 31288
rect 2700 31226 2728 31894
rect 2780 31816 2832 31822
rect 2976 31804 3004 32846
rect 3068 32065 3096 33487
rect 3160 33114 3188 35022
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3252 32570 3280 49302
rect 3330 49263 3386 49272
rect 3344 48822 3372 49263
rect 3332 48816 3384 48822
rect 3332 48758 3384 48764
rect 3436 48754 3464 51002
rect 3528 49434 3556 51190
rect 3516 49428 3568 49434
rect 3516 49370 3568 49376
rect 3620 48890 3648 70858
rect 3700 67856 3752 67862
rect 3700 67798 3752 67804
rect 3712 65142 3740 67798
rect 3700 65136 3752 65142
rect 3700 65078 3752 65084
rect 3700 65000 3752 65006
rect 3700 64942 3752 64948
rect 3712 62966 3740 64942
rect 3700 62960 3752 62966
rect 3700 62902 3752 62908
rect 3698 62792 3754 62801
rect 3698 62727 3700 62736
rect 3752 62727 3754 62736
rect 3700 62698 3752 62704
rect 3698 62656 3754 62665
rect 3698 62591 3754 62600
rect 3608 48884 3660 48890
rect 3608 48826 3660 48832
rect 3712 48770 3740 62591
rect 3804 50930 3832 76502
rect 3896 65686 3924 76622
rect 3988 74934 4016 76894
rect 4068 76832 4120 76838
rect 4068 76774 4120 76780
rect 4080 76362 4108 76774
rect 5846 76732 6154 76752
rect 5846 76730 5852 76732
rect 5908 76730 5932 76732
rect 5988 76730 6012 76732
rect 6068 76730 6092 76732
rect 6148 76730 6154 76732
rect 5908 76678 5910 76730
rect 6090 76678 6092 76730
rect 5846 76676 5852 76678
rect 5908 76676 5932 76678
rect 5988 76676 6012 76678
rect 6068 76676 6092 76678
rect 6148 76676 6154 76678
rect 5846 76656 6154 76676
rect 4068 76356 4120 76362
rect 4068 76298 4120 76304
rect 4214 76188 4522 76208
rect 4214 76186 4220 76188
rect 4276 76186 4300 76188
rect 4356 76186 4380 76188
rect 4436 76186 4460 76188
rect 4516 76186 4522 76188
rect 4276 76134 4278 76186
rect 4458 76134 4460 76186
rect 4214 76132 4220 76134
rect 4276 76132 4300 76134
rect 4356 76132 4380 76134
rect 4436 76132 4460 76134
rect 4516 76132 4522 76134
rect 4214 76112 4522 76132
rect 7478 76188 7786 76208
rect 7478 76186 7484 76188
rect 7540 76186 7564 76188
rect 7620 76186 7644 76188
rect 7700 76186 7724 76188
rect 7780 76186 7786 76188
rect 7540 76134 7542 76186
rect 7722 76134 7724 76186
rect 7478 76132 7484 76134
rect 7540 76132 7564 76134
rect 7620 76132 7644 76134
rect 7700 76132 7724 76134
rect 7780 76132 7786 76134
rect 7478 76112 7786 76132
rect 5846 75644 6154 75664
rect 5846 75642 5852 75644
rect 5908 75642 5932 75644
rect 5988 75642 6012 75644
rect 6068 75642 6092 75644
rect 6148 75642 6154 75644
rect 5908 75590 5910 75642
rect 6090 75590 6092 75642
rect 5846 75588 5852 75590
rect 5908 75588 5932 75590
rect 5988 75588 6012 75590
rect 6068 75588 6092 75590
rect 6148 75588 6154 75590
rect 5846 75568 6154 75588
rect 4214 75100 4522 75120
rect 4214 75098 4220 75100
rect 4276 75098 4300 75100
rect 4356 75098 4380 75100
rect 4436 75098 4460 75100
rect 4516 75098 4522 75100
rect 4276 75046 4278 75098
rect 4458 75046 4460 75098
rect 4214 75044 4220 75046
rect 4276 75044 4300 75046
rect 4356 75044 4380 75046
rect 4436 75044 4460 75046
rect 4516 75044 4522 75046
rect 4214 75024 4522 75044
rect 7478 75100 7786 75120
rect 7478 75098 7484 75100
rect 7540 75098 7564 75100
rect 7620 75098 7644 75100
rect 7700 75098 7724 75100
rect 7780 75098 7786 75100
rect 7540 75046 7542 75098
rect 7722 75046 7724 75098
rect 7478 75044 7484 75046
rect 7540 75044 7564 75046
rect 7620 75044 7644 75046
rect 7700 75044 7724 75046
rect 7780 75044 7786 75046
rect 7478 75024 7786 75044
rect 3976 74928 4028 74934
rect 3976 74870 4028 74876
rect 8312 74798 8340 77318
rect 9416 77217 9444 77454
rect 9402 77208 9458 77217
rect 9402 77143 9458 77152
rect 9508 77042 9536 77959
rect 9600 77042 9628 78639
rect 9968 77518 9996 79455
rect 9956 77512 10008 77518
rect 9956 77454 10008 77460
rect 9496 77036 9548 77042
rect 9496 76978 9548 76984
rect 9588 77036 9640 77042
rect 9588 76978 9640 76984
rect 9772 76832 9824 76838
rect 9772 76774 9824 76780
rect 9110 76732 9418 76752
rect 9110 76730 9116 76732
rect 9172 76730 9196 76732
rect 9252 76730 9276 76732
rect 9332 76730 9356 76732
rect 9412 76730 9418 76732
rect 9172 76678 9174 76730
rect 9354 76678 9356 76730
rect 9110 76676 9116 76678
rect 9172 76676 9196 76678
rect 9252 76676 9276 76678
rect 9332 76676 9356 76678
rect 9412 76676 9418 76678
rect 9110 76656 9418 76676
rect 9110 75644 9418 75664
rect 9110 75642 9116 75644
rect 9172 75642 9196 75644
rect 9252 75642 9276 75644
rect 9332 75642 9356 75644
rect 9412 75642 9418 75644
rect 9172 75590 9174 75642
rect 9354 75590 9356 75642
rect 9110 75588 9116 75590
rect 9172 75588 9196 75590
rect 9252 75588 9276 75590
rect 9332 75588 9356 75590
rect 9412 75588 9418 75590
rect 9110 75568 9418 75588
rect 8300 74792 8352 74798
rect 8300 74734 8352 74740
rect 5846 74556 6154 74576
rect 5846 74554 5852 74556
rect 5908 74554 5932 74556
rect 5988 74554 6012 74556
rect 6068 74554 6092 74556
rect 6148 74554 6154 74556
rect 5908 74502 5910 74554
rect 6090 74502 6092 74554
rect 5846 74500 5852 74502
rect 5908 74500 5932 74502
rect 5988 74500 6012 74502
rect 6068 74500 6092 74502
rect 6148 74500 6154 74502
rect 5846 74480 6154 74500
rect 9110 74556 9418 74576
rect 9110 74554 9116 74556
rect 9172 74554 9196 74556
rect 9252 74554 9276 74556
rect 9332 74554 9356 74556
rect 9412 74554 9418 74556
rect 9172 74502 9174 74554
rect 9354 74502 9356 74554
rect 9110 74500 9116 74502
rect 9172 74500 9196 74502
rect 9252 74500 9276 74502
rect 9332 74500 9356 74502
rect 9412 74500 9418 74502
rect 9110 74480 9418 74500
rect 4214 74012 4522 74032
rect 4214 74010 4220 74012
rect 4276 74010 4300 74012
rect 4356 74010 4380 74012
rect 4436 74010 4460 74012
rect 4516 74010 4522 74012
rect 4276 73958 4278 74010
rect 4458 73958 4460 74010
rect 4214 73956 4220 73958
rect 4276 73956 4300 73958
rect 4356 73956 4380 73958
rect 4436 73956 4460 73958
rect 4516 73956 4522 73958
rect 4214 73936 4522 73956
rect 7478 74012 7786 74032
rect 7478 74010 7484 74012
rect 7540 74010 7564 74012
rect 7620 74010 7644 74012
rect 7700 74010 7724 74012
rect 7780 74010 7786 74012
rect 7540 73958 7542 74010
rect 7722 73958 7724 74010
rect 7478 73956 7484 73958
rect 7540 73956 7564 73958
rect 7620 73956 7644 73958
rect 7700 73956 7724 73958
rect 7780 73956 7786 73958
rect 7478 73936 7786 73956
rect 5846 73468 6154 73488
rect 5846 73466 5852 73468
rect 5908 73466 5932 73468
rect 5988 73466 6012 73468
rect 6068 73466 6092 73468
rect 6148 73466 6154 73468
rect 5908 73414 5910 73466
rect 6090 73414 6092 73466
rect 5846 73412 5852 73414
rect 5908 73412 5932 73414
rect 5988 73412 6012 73414
rect 6068 73412 6092 73414
rect 6148 73412 6154 73414
rect 5846 73392 6154 73412
rect 9110 73468 9418 73488
rect 9110 73466 9116 73468
rect 9172 73466 9196 73468
rect 9252 73466 9276 73468
rect 9332 73466 9356 73468
rect 9412 73466 9418 73468
rect 9172 73414 9174 73466
rect 9354 73414 9356 73466
rect 9110 73412 9116 73414
rect 9172 73412 9196 73414
rect 9252 73412 9276 73414
rect 9332 73412 9356 73414
rect 9412 73412 9418 73414
rect 9110 73392 9418 73412
rect 4712 73024 4764 73030
rect 4712 72966 4764 72972
rect 4214 72924 4522 72944
rect 4214 72922 4220 72924
rect 4276 72922 4300 72924
rect 4356 72922 4380 72924
rect 4436 72922 4460 72924
rect 4516 72922 4522 72924
rect 4276 72870 4278 72922
rect 4458 72870 4460 72922
rect 4214 72868 4220 72870
rect 4276 72868 4300 72870
rect 4356 72868 4380 72870
rect 4436 72868 4460 72870
rect 4516 72868 4522 72870
rect 4214 72848 4522 72868
rect 4214 71836 4522 71856
rect 4214 71834 4220 71836
rect 4276 71834 4300 71836
rect 4356 71834 4380 71836
rect 4436 71834 4460 71836
rect 4516 71834 4522 71836
rect 4276 71782 4278 71834
rect 4458 71782 4460 71834
rect 4214 71780 4220 71782
rect 4276 71780 4300 71782
rect 4356 71780 4380 71782
rect 4436 71780 4460 71782
rect 4516 71780 4522 71782
rect 4214 71760 4522 71780
rect 3976 71392 4028 71398
rect 3976 71334 4028 71340
rect 3884 65680 3936 65686
rect 3884 65622 3936 65628
rect 3988 65532 4016 71334
rect 4214 70748 4522 70768
rect 4214 70746 4220 70748
rect 4276 70746 4300 70748
rect 4356 70746 4380 70748
rect 4436 70746 4460 70748
rect 4516 70746 4522 70748
rect 4276 70694 4278 70746
rect 4458 70694 4460 70746
rect 4214 70692 4220 70694
rect 4276 70692 4300 70694
rect 4356 70692 4380 70694
rect 4436 70692 4460 70694
rect 4516 70692 4522 70694
rect 4214 70672 4522 70692
rect 4214 69660 4522 69680
rect 4214 69658 4220 69660
rect 4276 69658 4300 69660
rect 4356 69658 4380 69660
rect 4436 69658 4460 69660
rect 4516 69658 4522 69660
rect 4276 69606 4278 69658
rect 4458 69606 4460 69658
rect 4214 69604 4220 69606
rect 4276 69604 4300 69606
rect 4356 69604 4380 69606
rect 4436 69604 4460 69606
rect 4516 69604 4522 69606
rect 4214 69584 4522 69604
rect 4214 68572 4522 68592
rect 4214 68570 4220 68572
rect 4276 68570 4300 68572
rect 4356 68570 4380 68572
rect 4436 68570 4460 68572
rect 4516 68570 4522 68572
rect 4276 68518 4278 68570
rect 4458 68518 4460 68570
rect 4214 68516 4220 68518
rect 4276 68516 4300 68518
rect 4356 68516 4380 68518
rect 4436 68516 4460 68518
rect 4516 68516 4522 68518
rect 4214 68496 4522 68516
rect 4620 68196 4672 68202
rect 4620 68138 4672 68144
rect 4214 67484 4522 67504
rect 4214 67482 4220 67484
rect 4276 67482 4300 67484
rect 4356 67482 4380 67484
rect 4436 67482 4460 67484
rect 4516 67482 4522 67484
rect 4276 67430 4278 67482
rect 4458 67430 4460 67482
rect 4214 67428 4220 67430
rect 4276 67428 4300 67430
rect 4356 67428 4380 67430
rect 4436 67428 4460 67430
rect 4516 67428 4522 67430
rect 4214 67408 4522 67428
rect 4214 66396 4522 66416
rect 4214 66394 4220 66396
rect 4276 66394 4300 66396
rect 4356 66394 4380 66396
rect 4436 66394 4460 66396
rect 4516 66394 4522 66396
rect 4276 66342 4278 66394
rect 4458 66342 4460 66394
rect 4214 66340 4220 66342
rect 4276 66340 4300 66342
rect 4356 66340 4380 66342
rect 4436 66340 4460 66342
rect 4516 66340 4522 66342
rect 4214 66320 4522 66340
rect 3896 65504 4016 65532
rect 4068 65544 4120 65550
rect 3792 50924 3844 50930
rect 3792 50866 3844 50872
rect 3896 49473 3924 65504
rect 4068 65486 4120 65492
rect 3976 65408 4028 65414
rect 3976 65350 4028 65356
rect 3988 65249 4016 65350
rect 3974 65240 4030 65249
rect 3974 65175 4030 65184
rect 3976 65136 4028 65142
rect 3976 65078 4028 65084
rect 3988 62665 4016 65078
rect 3974 62656 4030 62665
rect 3974 62591 4030 62600
rect 3976 62484 4028 62490
rect 3976 62426 4028 62432
rect 3988 60897 4016 62426
rect 3974 60888 4030 60897
rect 3974 60823 4030 60832
rect 3974 60752 4030 60761
rect 3974 60687 3976 60696
rect 4028 60687 4030 60696
rect 3976 60658 4028 60664
rect 3974 60616 4030 60625
rect 3974 60551 4030 60560
rect 3988 56930 4016 60551
rect 4080 57050 4108 65486
rect 4214 65308 4522 65328
rect 4214 65306 4220 65308
rect 4276 65306 4300 65308
rect 4356 65306 4380 65308
rect 4436 65306 4460 65308
rect 4516 65306 4522 65308
rect 4276 65254 4278 65306
rect 4458 65254 4460 65306
rect 4214 65252 4220 65254
rect 4276 65252 4300 65254
rect 4356 65252 4380 65254
rect 4436 65252 4460 65254
rect 4516 65252 4522 65254
rect 4214 65232 4522 65252
rect 4214 64220 4522 64240
rect 4214 64218 4220 64220
rect 4276 64218 4300 64220
rect 4356 64218 4380 64220
rect 4436 64218 4460 64220
rect 4516 64218 4522 64220
rect 4276 64166 4278 64218
rect 4458 64166 4460 64218
rect 4214 64164 4220 64166
rect 4276 64164 4300 64166
rect 4356 64164 4380 64166
rect 4436 64164 4460 64166
rect 4516 64164 4522 64166
rect 4214 64144 4522 64164
rect 4214 63132 4522 63152
rect 4214 63130 4220 63132
rect 4276 63130 4300 63132
rect 4356 63130 4380 63132
rect 4436 63130 4460 63132
rect 4516 63130 4522 63132
rect 4276 63078 4278 63130
rect 4458 63078 4460 63130
rect 4214 63076 4220 63078
rect 4276 63076 4300 63078
rect 4356 63076 4380 63078
rect 4436 63076 4460 63078
rect 4516 63076 4522 63078
rect 4214 63056 4522 63076
rect 4214 62044 4522 62064
rect 4214 62042 4220 62044
rect 4276 62042 4300 62044
rect 4356 62042 4380 62044
rect 4436 62042 4460 62044
rect 4516 62042 4522 62044
rect 4276 61990 4278 62042
rect 4458 61990 4460 62042
rect 4214 61988 4220 61990
rect 4276 61988 4300 61990
rect 4356 61988 4380 61990
rect 4436 61988 4460 61990
rect 4516 61988 4522 61990
rect 4214 61968 4522 61988
rect 4214 60956 4522 60976
rect 4214 60954 4220 60956
rect 4276 60954 4300 60956
rect 4356 60954 4380 60956
rect 4436 60954 4460 60956
rect 4516 60954 4522 60956
rect 4276 60902 4278 60954
rect 4458 60902 4460 60954
rect 4214 60900 4220 60902
rect 4276 60900 4300 60902
rect 4356 60900 4380 60902
rect 4436 60900 4460 60902
rect 4516 60900 4522 60902
rect 4214 60880 4522 60900
rect 4214 59868 4522 59888
rect 4214 59866 4220 59868
rect 4276 59866 4300 59868
rect 4356 59866 4380 59868
rect 4436 59866 4460 59868
rect 4516 59866 4522 59868
rect 4276 59814 4278 59866
rect 4458 59814 4460 59866
rect 4214 59812 4220 59814
rect 4276 59812 4300 59814
rect 4356 59812 4380 59814
rect 4436 59812 4460 59814
rect 4516 59812 4522 59814
rect 4214 59792 4522 59812
rect 4214 58780 4522 58800
rect 4214 58778 4220 58780
rect 4276 58778 4300 58780
rect 4356 58778 4380 58780
rect 4436 58778 4460 58780
rect 4516 58778 4522 58780
rect 4276 58726 4278 58778
rect 4458 58726 4460 58778
rect 4214 58724 4220 58726
rect 4276 58724 4300 58726
rect 4356 58724 4380 58726
rect 4436 58724 4460 58726
rect 4516 58724 4522 58726
rect 4214 58704 4522 58724
rect 4214 57692 4522 57712
rect 4214 57690 4220 57692
rect 4276 57690 4300 57692
rect 4356 57690 4380 57692
rect 4436 57690 4460 57692
rect 4516 57690 4522 57692
rect 4276 57638 4278 57690
rect 4458 57638 4460 57690
rect 4214 57636 4220 57638
rect 4276 57636 4300 57638
rect 4356 57636 4380 57638
rect 4436 57636 4460 57638
rect 4516 57636 4522 57638
rect 4214 57616 4522 57636
rect 4068 57044 4120 57050
rect 4068 56986 4120 56992
rect 3988 56902 4108 56930
rect 3976 56840 4028 56846
rect 3976 56782 4028 56788
rect 3988 56506 4016 56782
rect 3976 56500 4028 56506
rect 3976 56442 4028 56448
rect 3976 55888 4028 55894
rect 3976 55830 4028 55836
rect 3988 55457 4016 55830
rect 3974 55448 4030 55457
rect 3974 55383 4030 55392
rect 3976 53168 4028 53174
rect 3976 53110 4028 53116
rect 3988 51066 4016 53110
rect 3976 51060 4028 51066
rect 4080 51048 4108 56902
rect 4214 56604 4522 56624
rect 4214 56602 4220 56604
rect 4276 56602 4300 56604
rect 4356 56602 4380 56604
rect 4436 56602 4460 56604
rect 4516 56602 4522 56604
rect 4276 56550 4278 56602
rect 4458 56550 4460 56602
rect 4214 56548 4220 56550
rect 4276 56548 4300 56550
rect 4356 56548 4380 56550
rect 4436 56548 4460 56550
rect 4516 56548 4522 56550
rect 4214 56528 4522 56548
rect 4160 56432 4212 56438
rect 4160 56374 4212 56380
rect 4172 55865 4200 56374
rect 4632 55865 4660 68138
rect 4724 56438 4752 72966
rect 7478 72924 7786 72944
rect 7478 72922 7484 72924
rect 7540 72922 7564 72924
rect 7620 72922 7644 72924
rect 7700 72922 7724 72924
rect 7780 72922 7786 72924
rect 7540 72870 7542 72922
rect 7722 72870 7724 72922
rect 7478 72868 7484 72870
rect 7540 72868 7564 72870
rect 7620 72868 7644 72870
rect 7700 72868 7724 72870
rect 7780 72868 7786 72870
rect 7478 72848 7786 72868
rect 8300 72480 8352 72486
rect 8300 72422 8352 72428
rect 5846 72380 6154 72400
rect 5846 72378 5852 72380
rect 5908 72378 5932 72380
rect 5988 72378 6012 72380
rect 6068 72378 6092 72380
rect 6148 72378 6154 72380
rect 5908 72326 5910 72378
rect 6090 72326 6092 72378
rect 5846 72324 5852 72326
rect 5908 72324 5932 72326
rect 5988 72324 6012 72326
rect 6068 72324 6092 72326
rect 6148 72324 6154 72326
rect 5846 72304 6154 72324
rect 7478 71836 7786 71856
rect 7478 71834 7484 71836
rect 7540 71834 7564 71836
rect 7620 71834 7644 71836
rect 7700 71834 7724 71836
rect 7780 71834 7786 71836
rect 7540 71782 7542 71834
rect 7722 71782 7724 71834
rect 7478 71780 7484 71782
rect 7540 71780 7564 71782
rect 7620 71780 7644 71782
rect 7700 71780 7724 71782
rect 7780 71780 7786 71782
rect 7478 71760 7786 71780
rect 8312 71534 8340 72422
rect 9110 72380 9418 72400
rect 9110 72378 9116 72380
rect 9172 72378 9196 72380
rect 9252 72378 9276 72380
rect 9332 72378 9356 72380
rect 9412 72378 9418 72380
rect 9172 72326 9174 72378
rect 9354 72326 9356 72378
rect 9110 72324 9116 72326
rect 9172 72324 9196 72326
rect 9252 72324 9276 72326
rect 9332 72324 9356 72326
rect 9412 72324 9418 72326
rect 9110 72304 9418 72324
rect 8300 71528 8352 71534
rect 8300 71470 8352 71476
rect 5846 71292 6154 71312
rect 5846 71290 5852 71292
rect 5908 71290 5932 71292
rect 5988 71290 6012 71292
rect 6068 71290 6092 71292
rect 6148 71290 6154 71292
rect 5908 71238 5910 71290
rect 6090 71238 6092 71290
rect 5846 71236 5852 71238
rect 5908 71236 5932 71238
rect 5988 71236 6012 71238
rect 6068 71236 6092 71238
rect 6148 71236 6154 71238
rect 5846 71216 6154 71236
rect 9110 71292 9418 71312
rect 9110 71290 9116 71292
rect 9172 71290 9196 71292
rect 9252 71290 9276 71292
rect 9332 71290 9356 71292
rect 9412 71290 9418 71292
rect 9172 71238 9174 71290
rect 9354 71238 9356 71290
rect 9110 71236 9116 71238
rect 9172 71236 9196 71238
rect 9252 71236 9276 71238
rect 9332 71236 9356 71238
rect 9412 71236 9418 71238
rect 9110 71216 9418 71236
rect 7478 70748 7786 70768
rect 7478 70746 7484 70748
rect 7540 70746 7564 70748
rect 7620 70746 7644 70748
rect 7700 70746 7724 70748
rect 7780 70746 7786 70748
rect 7540 70694 7542 70746
rect 7722 70694 7724 70746
rect 7478 70692 7484 70694
rect 7540 70692 7564 70694
rect 7620 70692 7644 70694
rect 7700 70692 7724 70694
rect 7780 70692 7786 70694
rect 7478 70672 7786 70692
rect 5846 70204 6154 70224
rect 5846 70202 5852 70204
rect 5908 70202 5932 70204
rect 5988 70202 6012 70204
rect 6068 70202 6092 70204
rect 6148 70202 6154 70204
rect 5908 70150 5910 70202
rect 6090 70150 6092 70202
rect 5846 70148 5852 70150
rect 5908 70148 5932 70150
rect 5988 70148 6012 70150
rect 6068 70148 6092 70150
rect 6148 70148 6154 70150
rect 5846 70128 6154 70148
rect 9110 70204 9418 70224
rect 9110 70202 9116 70204
rect 9172 70202 9196 70204
rect 9252 70202 9276 70204
rect 9332 70202 9356 70204
rect 9412 70202 9418 70204
rect 9172 70150 9174 70202
rect 9354 70150 9356 70202
rect 9110 70148 9116 70150
rect 9172 70148 9196 70150
rect 9252 70148 9276 70150
rect 9332 70148 9356 70150
rect 9412 70148 9418 70150
rect 9110 70128 9418 70148
rect 7478 69660 7786 69680
rect 7478 69658 7484 69660
rect 7540 69658 7564 69660
rect 7620 69658 7644 69660
rect 7700 69658 7724 69660
rect 7780 69658 7786 69660
rect 7540 69606 7542 69658
rect 7722 69606 7724 69658
rect 7478 69604 7484 69606
rect 7540 69604 7564 69606
rect 7620 69604 7644 69606
rect 7700 69604 7724 69606
rect 7780 69604 7786 69606
rect 7478 69584 7786 69604
rect 5846 69116 6154 69136
rect 5846 69114 5852 69116
rect 5908 69114 5932 69116
rect 5988 69114 6012 69116
rect 6068 69114 6092 69116
rect 6148 69114 6154 69116
rect 5908 69062 5910 69114
rect 6090 69062 6092 69114
rect 5846 69060 5852 69062
rect 5908 69060 5932 69062
rect 5988 69060 6012 69062
rect 6068 69060 6092 69062
rect 6148 69060 6154 69062
rect 5846 69040 6154 69060
rect 9110 69116 9418 69136
rect 9110 69114 9116 69116
rect 9172 69114 9196 69116
rect 9252 69114 9276 69116
rect 9332 69114 9356 69116
rect 9412 69114 9418 69116
rect 9172 69062 9174 69114
rect 9354 69062 9356 69114
rect 9110 69060 9116 69062
rect 9172 69060 9196 69062
rect 9252 69060 9276 69062
rect 9332 69060 9356 69062
rect 9412 69060 9418 69062
rect 9110 69040 9418 69060
rect 4896 69012 4948 69018
rect 4896 68954 4948 68960
rect 4804 64592 4856 64598
rect 4804 64534 4856 64540
rect 4712 56432 4764 56438
rect 4712 56374 4764 56380
rect 4816 55978 4844 64534
rect 4724 55950 4844 55978
rect 4158 55856 4214 55865
rect 4158 55791 4214 55800
rect 4618 55856 4674 55865
rect 4618 55791 4674 55800
rect 4172 55758 4200 55791
rect 4160 55752 4212 55758
rect 4160 55694 4212 55700
rect 4620 55752 4672 55758
rect 4620 55694 4672 55700
rect 4214 55516 4522 55536
rect 4214 55514 4220 55516
rect 4276 55514 4300 55516
rect 4356 55514 4380 55516
rect 4436 55514 4460 55516
rect 4516 55514 4522 55516
rect 4276 55462 4278 55514
rect 4458 55462 4460 55514
rect 4214 55460 4220 55462
rect 4276 55460 4300 55462
rect 4356 55460 4380 55462
rect 4436 55460 4460 55462
rect 4516 55460 4522 55462
rect 4214 55440 4522 55460
rect 4158 55312 4214 55321
rect 4158 55247 4160 55256
rect 4212 55247 4214 55256
rect 4160 55218 4212 55224
rect 4214 54428 4522 54448
rect 4214 54426 4220 54428
rect 4276 54426 4300 54428
rect 4356 54426 4380 54428
rect 4436 54426 4460 54428
rect 4516 54426 4522 54428
rect 4276 54374 4278 54426
rect 4458 54374 4460 54426
rect 4214 54372 4220 54374
rect 4276 54372 4300 54374
rect 4356 54372 4380 54374
rect 4436 54372 4460 54374
rect 4516 54372 4522 54374
rect 4214 54352 4522 54372
rect 4436 54120 4488 54126
rect 4436 54062 4488 54068
rect 4448 53689 4476 54062
rect 4528 54052 4580 54058
rect 4528 53994 4580 54000
rect 4434 53680 4490 53689
rect 4434 53615 4490 53624
rect 4540 53553 4568 53994
rect 4526 53544 4582 53553
rect 4526 53479 4582 53488
rect 4214 53340 4522 53360
rect 4214 53338 4220 53340
rect 4276 53338 4300 53340
rect 4356 53338 4380 53340
rect 4436 53338 4460 53340
rect 4516 53338 4522 53340
rect 4276 53286 4278 53338
rect 4458 53286 4460 53338
rect 4214 53284 4220 53286
rect 4276 53284 4300 53286
rect 4356 53284 4380 53286
rect 4436 53284 4460 53286
rect 4516 53284 4522 53286
rect 4214 53264 4522 53284
rect 4214 52252 4522 52272
rect 4214 52250 4220 52252
rect 4276 52250 4300 52252
rect 4356 52250 4380 52252
rect 4436 52250 4460 52252
rect 4516 52250 4522 52252
rect 4276 52198 4278 52250
rect 4458 52198 4460 52250
rect 4214 52196 4220 52198
rect 4276 52196 4300 52198
rect 4356 52196 4380 52198
rect 4436 52196 4460 52198
rect 4516 52196 4522 52198
rect 4214 52176 4522 52196
rect 4214 51164 4522 51184
rect 4214 51162 4220 51164
rect 4276 51162 4300 51164
rect 4356 51162 4380 51164
rect 4436 51162 4460 51164
rect 4516 51162 4522 51164
rect 4276 51110 4278 51162
rect 4458 51110 4460 51162
rect 4214 51108 4220 51110
rect 4276 51108 4300 51110
rect 4356 51108 4380 51110
rect 4436 51108 4460 51110
rect 4516 51108 4522 51110
rect 4214 51088 4522 51108
rect 4080 51020 4292 51048
rect 3976 51002 4028 51008
rect 4068 50924 4120 50930
rect 4068 50866 4120 50872
rect 3882 49464 3938 49473
rect 3882 49399 3938 49408
rect 3884 49360 3936 49366
rect 3884 49302 3936 49308
rect 3424 48748 3476 48754
rect 3424 48690 3476 48696
rect 3620 48742 3740 48770
rect 3332 48680 3384 48686
rect 3384 48628 3556 48634
rect 3332 48622 3556 48628
rect 3344 48606 3556 48622
rect 3332 48544 3384 48550
rect 3332 48486 3384 48492
rect 3424 48544 3476 48550
rect 3424 48486 3476 48492
rect 3344 46102 3372 48486
rect 3436 46714 3464 48486
rect 3424 46708 3476 46714
rect 3424 46650 3476 46656
rect 3424 46572 3476 46578
rect 3424 46514 3476 46520
rect 3436 46481 3464 46514
rect 3422 46472 3478 46481
rect 3422 46407 3478 46416
rect 3528 46186 3556 48606
rect 3436 46158 3556 46186
rect 3332 46096 3384 46102
rect 3332 46038 3384 46044
rect 3332 45960 3384 45966
rect 3332 45902 3384 45908
rect 3344 44538 3372 45902
rect 3332 44532 3384 44538
rect 3332 44474 3384 44480
rect 3332 44328 3384 44334
rect 3332 44270 3384 44276
rect 3344 43994 3372 44270
rect 3332 43988 3384 43994
rect 3332 43930 3384 43936
rect 3332 43784 3384 43790
rect 3332 43726 3384 43732
rect 3344 43450 3372 43726
rect 3332 43444 3384 43450
rect 3332 43386 3384 43392
rect 3332 43308 3384 43314
rect 3332 43250 3384 43256
rect 3344 42906 3372 43250
rect 3332 42900 3384 42906
rect 3332 42842 3384 42848
rect 3344 42362 3372 42842
rect 3332 42356 3384 42362
rect 3332 42298 3384 42304
rect 3330 42256 3386 42265
rect 3330 42191 3386 42200
rect 3240 32564 3292 32570
rect 3240 32506 3292 32512
rect 3240 32360 3292 32366
rect 3240 32302 3292 32308
rect 3054 32056 3110 32065
rect 3054 31991 3110 32000
rect 2832 31776 3004 31804
rect 2780 31758 2832 31764
rect 2792 31385 2820 31758
rect 3252 31482 3280 32302
rect 3344 31822 3372 42191
rect 3436 37942 3464 46158
rect 3516 46096 3568 46102
rect 3516 46038 3568 46044
rect 3528 42702 3556 46038
rect 3620 43178 3648 48742
rect 3792 48544 3844 48550
rect 3896 48532 3924 49302
rect 3976 49224 4028 49230
rect 3974 49192 3976 49201
rect 4028 49192 4030 49201
rect 3974 49127 4030 49136
rect 3976 49088 4028 49094
rect 3974 49056 3976 49065
rect 4028 49056 4030 49065
rect 3974 48991 4030 49000
rect 3974 48920 4030 48929
rect 3974 48855 4030 48864
rect 4080 48872 4108 50866
rect 4264 50425 4292 51020
rect 4250 50416 4306 50425
rect 4250 50351 4306 50360
rect 4214 50076 4522 50096
rect 4214 50074 4220 50076
rect 4276 50074 4300 50076
rect 4356 50074 4380 50076
rect 4436 50074 4460 50076
rect 4516 50074 4522 50076
rect 4276 50022 4278 50074
rect 4458 50022 4460 50074
rect 4214 50020 4220 50022
rect 4276 50020 4300 50022
rect 4356 50020 4380 50022
rect 4436 50020 4460 50022
rect 4516 50020 4522 50022
rect 4214 50000 4522 50020
rect 4528 49904 4580 49910
rect 4528 49846 4580 49852
rect 4540 49201 4568 49846
rect 4526 49192 4582 49201
rect 4526 49127 4582 49136
rect 4214 48988 4522 49008
rect 4214 48986 4220 48988
rect 4276 48986 4300 48988
rect 4356 48986 4380 48988
rect 4436 48986 4460 48988
rect 4516 48986 4522 48988
rect 4276 48934 4278 48986
rect 4458 48934 4460 48986
rect 4214 48932 4220 48934
rect 4276 48932 4300 48934
rect 4356 48932 4380 48934
rect 4436 48932 4460 48934
rect 4516 48932 4522 48934
rect 4214 48912 4522 48932
rect 3988 48657 4016 48855
rect 4080 48844 4384 48872
rect 4068 48748 4120 48754
rect 4068 48690 4120 48696
rect 3974 48648 4030 48657
rect 3974 48583 4030 48592
rect 3896 48504 4016 48532
rect 3792 48486 3844 48492
rect 3700 48272 3752 48278
rect 3804 48249 3832 48486
rect 3882 48376 3938 48385
rect 3882 48311 3938 48320
rect 3700 48214 3752 48220
rect 3790 48240 3846 48249
rect 3712 43314 3740 48214
rect 3790 48175 3846 48184
rect 3790 48104 3846 48113
rect 3790 48039 3846 48048
rect 3804 47666 3832 48039
rect 3792 47660 3844 47666
rect 3792 47602 3844 47608
rect 3792 47456 3844 47462
rect 3792 47398 3844 47404
rect 3804 45665 3832 47398
rect 3790 45656 3846 45665
rect 3790 45591 3846 45600
rect 3792 45552 3844 45558
rect 3792 45494 3844 45500
rect 3804 44402 3832 45494
rect 3792 44396 3844 44402
rect 3792 44338 3844 44344
rect 3792 43988 3844 43994
rect 3792 43930 3844 43936
rect 3700 43308 3752 43314
rect 3700 43250 3752 43256
rect 3804 43194 3832 43930
rect 3608 43172 3660 43178
rect 3608 43114 3660 43120
rect 3712 43166 3832 43194
rect 3606 43072 3662 43081
rect 3606 43007 3662 43016
rect 3516 42696 3568 42702
rect 3516 42638 3568 42644
rect 3620 41721 3648 43007
rect 3606 41712 3662 41721
rect 3712 41682 3740 43166
rect 3792 43104 3844 43110
rect 3792 43046 3844 43052
rect 3606 41647 3662 41656
rect 3700 41676 3752 41682
rect 3700 41618 3752 41624
rect 3516 41200 3568 41206
rect 3516 41142 3568 41148
rect 3606 41168 3662 41177
rect 3528 38282 3556 41142
rect 3606 41103 3662 41112
rect 3516 38276 3568 38282
rect 3516 38218 3568 38224
rect 3424 37936 3476 37942
rect 3424 37878 3476 37884
rect 3528 37754 3556 38218
rect 3436 37726 3556 37754
rect 3436 32366 3464 37726
rect 3516 36780 3568 36786
rect 3516 36722 3568 36728
rect 3424 32360 3476 32366
rect 3528 32337 3556 36722
rect 3424 32302 3476 32308
rect 3514 32328 3570 32337
rect 3514 32263 3570 32272
rect 3422 32192 3478 32201
rect 3478 32150 3556 32178
rect 3422 32127 3478 32136
rect 3424 31952 3476 31958
rect 3424 31894 3476 31900
rect 3332 31816 3384 31822
rect 3332 31758 3384 31764
rect 3332 31680 3384 31686
rect 3330 31648 3332 31657
rect 3384 31648 3386 31657
rect 3330 31583 3386 31592
rect 3330 31512 3386 31521
rect 3056 31476 3108 31482
rect 3056 31418 3108 31424
rect 3240 31476 3292 31482
rect 3330 31447 3386 31456
rect 3240 31418 3292 31424
rect 2778 31376 2834 31385
rect 2778 31311 2834 31320
rect 2516 31198 2728 31226
rect 2516 28966 2544 31198
rect 2964 31136 3016 31142
rect 2964 31078 3016 31084
rect 2582 31036 2890 31056
rect 2582 31034 2588 31036
rect 2644 31034 2668 31036
rect 2724 31034 2748 31036
rect 2804 31034 2828 31036
rect 2884 31034 2890 31036
rect 2644 30982 2646 31034
rect 2826 30982 2828 31034
rect 2582 30980 2588 30982
rect 2644 30980 2668 30982
rect 2724 30980 2748 30982
rect 2804 30980 2828 30982
rect 2884 30980 2890 30982
rect 2582 30960 2890 30980
rect 2976 30841 3004 31078
rect 2962 30832 3018 30841
rect 2962 30767 3018 30776
rect 3068 30682 3096 31418
rect 2976 30654 3096 30682
rect 2778 30424 2834 30433
rect 2778 30359 2834 30368
rect 2594 30288 2650 30297
rect 2594 30223 2596 30232
rect 2648 30223 2650 30232
rect 2596 30194 2648 30200
rect 2792 30122 2820 30359
rect 2780 30116 2832 30122
rect 2780 30058 2832 30064
rect 2582 29948 2890 29968
rect 2582 29946 2588 29948
rect 2644 29946 2668 29948
rect 2724 29946 2748 29948
rect 2804 29946 2828 29948
rect 2884 29946 2890 29948
rect 2644 29894 2646 29946
rect 2826 29894 2828 29946
rect 2582 29892 2588 29894
rect 2644 29892 2668 29894
rect 2724 29892 2748 29894
rect 2804 29892 2828 29894
rect 2884 29892 2890 29894
rect 2582 29872 2890 29892
rect 2976 29730 3004 30654
rect 3146 30560 3202 30569
rect 3146 30495 3202 30504
rect 3054 30424 3110 30433
rect 3054 30359 3110 30368
rect 2884 29702 3004 29730
rect 2884 29034 2912 29702
rect 2964 29164 3016 29170
rect 2964 29106 3016 29112
rect 2872 29028 2924 29034
rect 2872 28970 2924 28976
rect 2504 28960 2556 28966
rect 2504 28902 2556 28908
rect 2582 28860 2890 28880
rect 2582 28858 2588 28860
rect 2644 28858 2668 28860
rect 2724 28858 2748 28860
rect 2804 28858 2828 28860
rect 2884 28858 2890 28860
rect 2644 28806 2646 28858
rect 2826 28806 2828 28858
rect 2582 28804 2588 28806
rect 2644 28804 2668 28806
rect 2724 28804 2748 28806
rect 2804 28804 2828 28806
rect 2884 28804 2890 28806
rect 2582 28784 2890 28804
rect 2504 28756 2556 28762
rect 2504 28698 2556 28704
rect 2240 28648 2452 28676
rect 2240 28540 2268 28648
rect 2148 28529 2268 28540
rect 2134 28520 2268 28529
rect 1952 28484 2004 28490
rect 2190 28512 2268 28520
rect 2412 28552 2464 28558
rect 2412 28494 2464 28500
rect 2134 28455 2190 28464
rect 2320 28484 2372 28490
rect 1952 28426 2004 28432
rect 2320 28426 2372 28432
rect 1964 28121 1992 28426
rect 2226 28384 2282 28393
rect 2226 28319 2282 28328
rect 2134 28248 2190 28257
rect 2134 28183 2190 28192
rect 1950 28112 2006 28121
rect 1950 28047 2006 28056
rect 1950 27976 2006 27985
rect 1950 27911 2006 27920
rect 1860 25492 1912 25498
rect 1860 25434 1912 25440
rect 1860 25220 1912 25226
rect 1860 25162 1912 25168
rect 1872 24041 1900 25162
rect 1858 24032 1914 24041
rect 1858 23967 1914 23976
rect 1780 23854 1900 23882
rect 1768 22976 1820 22982
rect 1768 22918 1820 22924
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 1780 19922 1808 22918
rect 1584 19916 1636 19922
rect 1584 19858 1636 19864
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1492 19372 1544 19378
rect 1872 19334 1900 23854
rect 1964 22098 1992 27911
rect 2044 26988 2096 26994
rect 2044 26930 2096 26936
rect 2056 26586 2084 26930
rect 2148 26926 2176 28183
rect 2136 26920 2188 26926
rect 2136 26862 2188 26868
rect 2044 26580 2096 26586
rect 2044 26522 2096 26528
rect 2148 26518 2176 26862
rect 2136 26512 2188 26518
rect 2136 26454 2188 26460
rect 2044 25900 2096 25906
rect 2044 25842 2096 25848
rect 1952 22092 2004 22098
rect 1952 22034 2004 22040
rect 1952 20936 2004 20942
rect 1952 20878 2004 20884
rect 1492 19314 1544 19320
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1780 19306 1900 19334
rect 1412 18873 1440 19246
rect 1398 18864 1454 18873
rect 1398 18799 1454 18808
rect 1780 18408 1808 19306
rect 1780 18380 1900 18408
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1596 16697 1624 17614
rect 1676 17604 1728 17610
rect 1676 17546 1728 17552
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 14657 1440 16050
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1398 14648 1454 14657
rect 1398 14583 1454 14592
rect 1504 14482 1532 15846
rect 1596 15502 1624 16390
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1688 14906 1716 17546
rect 1596 14878 1716 14906
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1596 14278 1624 14878
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1688 14414 1716 14758
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1400 13728 1452 13734
rect 1400 13670 1452 13676
rect 1412 12918 1440 13670
rect 1400 12912 1452 12918
rect 1400 12854 1452 12860
rect 1504 12481 1532 13874
rect 1780 13870 1808 14554
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1490 12472 1546 12481
rect 1490 12407 1546 12416
rect 1596 12073 1624 13262
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1688 12850 1716 13126
rect 1768 12912 1820 12918
rect 1768 12854 1820 12860
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1582 12064 1638 12073
rect 1582 11999 1638 12008
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 10849 1440 11630
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1398 10840 1454 10849
rect 1398 10775 1454 10784
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1412 9897 1440 10542
rect 1504 10441 1532 11086
rect 1490 10432 1546 10441
rect 1490 10367 1546 10376
rect 1780 10130 1808 12854
rect 1768 10124 1820 10130
rect 1768 10066 1820 10072
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1398 9888 1454 9897
rect 1398 9823 1454 9832
rect 1400 9512 1452 9518
rect 1504 9489 1532 9998
rect 1400 9454 1452 9460
rect 1490 9480 1546 9489
rect 1412 9081 1440 9454
rect 1490 9415 1546 9424
rect 1398 9072 1454 9081
rect 1398 9007 1454 9016
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 8673 1440 8910
rect 1398 8664 1454 8673
rect 1398 8599 1454 8608
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8265 1440 8366
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1400 7880 1452 7886
rect 1398 7848 1400 7857
rect 1584 7880 1636 7886
rect 1452 7848 1454 7857
rect 1584 7822 1636 7828
rect 1398 7783 1454 7792
rect 1228 6886 1348 6914
rect 1228 4010 1256 6886
rect 1400 5704 1452 5710
rect 1306 5672 1362 5681
rect 1400 5646 1452 5652
rect 1306 5607 1362 5616
rect 1320 5234 1348 5607
rect 1412 5273 1440 5646
rect 1398 5264 1454 5273
rect 1308 5228 1360 5234
rect 1398 5199 1454 5208
rect 1308 5170 1360 5176
rect 1490 4040 1546 4049
rect 1216 4004 1268 4010
rect 1490 3975 1546 3984
rect 1216 3946 1268 3952
rect 1398 3632 1454 3641
rect 1398 3567 1454 3576
rect 1412 3058 1440 3567
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1504 2446 1532 3975
rect 1596 3618 1624 7822
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1688 6322 1716 6598
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1780 4078 1808 6734
rect 1872 6458 1900 18380
rect 1964 18358 1992 20878
rect 1952 18352 2004 18358
rect 1952 18294 2004 18300
rect 1964 17882 1992 18294
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 2056 17218 2084 25842
rect 2136 24744 2188 24750
rect 2136 24686 2188 24692
rect 2148 23118 2176 24686
rect 2240 24342 2268 28319
rect 2332 24886 2360 28426
rect 2320 24880 2372 24886
rect 2320 24822 2372 24828
rect 2228 24336 2280 24342
rect 2228 24278 2280 24284
rect 2424 24256 2452 28494
rect 2332 24228 2452 24256
rect 2136 23112 2188 23118
rect 2136 23054 2188 23060
rect 2148 22098 2176 23054
rect 2332 22982 2360 24228
rect 2410 24168 2466 24177
rect 2410 24103 2466 24112
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2320 22568 2372 22574
rect 2320 22510 2372 22516
rect 2332 22234 2360 22510
rect 2320 22228 2372 22234
rect 2320 22170 2372 22176
rect 2228 22160 2280 22166
rect 2228 22102 2280 22108
rect 2136 22092 2188 22098
rect 2136 22034 2188 22040
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2148 18970 2176 19858
rect 2136 18964 2188 18970
rect 2136 18906 2188 18912
rect 1964 17190 2084 17218
rect 1964 14362 1992 17190
rect 2240 16454 2268 22102
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2332 18222 2360 22034
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2424 18034 2452 24103
rect 2516 18834 2544 28698
rect 2976 28694 3004 29106
rect 2964 28688 3016 28694
rect 2594 28656 2650 28665
rect 2964 28630 3016 28636
rect 2594 28591 2650 28600
rect 2608 28558 2636 28591
rect 2596 28552 2648 28558
rect 2596 28494 2648 28500
rect 3068 28150 3096 30359
rect 3056 28144 3108 28150
rect 3056 28086 3108 28092
rect 2964 28076 3016 28082
rect 2964 28018 3016 28024
rect 2582 27772 2890 27792
rect 2582 27770 2588 27772
rect 2644 27770 2668 27772
rect 2724 27770 2748 27772
rect 2804 27770 2828 27772
rect 2884 27770 2890 27772
rect 2644 27718 2646 27770
rect 2826 27718 2828 27770
rect 2582 27716 2588 27718
rect 2644 27716 2668 27718
rect 2724 27716 2748 27718
rect 2804 27716 2828 27718
rect 2884 27716 2890 27718
rect 2582 27696 2890 27716
rect 2976 27554 3004 28018
rect 3056 28008 3108 28014
rect 3054 27976 3056 27985
rect 3108 27976 3110 27985
rect 3054 27911 3110 27920
rect 2884 27526 3004 27554
rect 2884 27033 2912 27526
rect 3056 27396 3108 27402
rect 3056 27338 3108 27344
rect 2870 27024 2926 27033
rect 2870 26959 2926 26968
rect 2582 26684 2890 26704
rect 2582 26682 2588 26684
rect 2644 26682 2668 26684
rect 2724 26682 2748 26684
rect 2804 26682 2828 26684
rect 2884 26682 2890 26684
rect 2644 26630 2646 26682
rect 2826 26630 2828 26682
rect 2582 26628 2588 26630
rect 2644 26628 2668 26630
rect 2724 26628 2748 26630
rect 2804 26628 2828 26630
rect 2884 26628 2890 26630
rect 2582 26608 2890 26628
rect 3068 26489 3096 27338
rect 3160 26518 3188 30495
rect 3240 29640 3292 29646
rect 3240 29582 3292 29588
rect 3148 26512 3200 26518
rect 3054 26480 3110 26489
rect 3148 26454 3200 26460
rect 3054 26415 3110 26424
rect 3146 26344 3202 26353
rect 2596 26308 2648 26314
rect 3146 26279 3202 26288
rect 2596 26250 2648 26256
rect 2608 26081 2636 26250
rect 3056 26240 3108 26246
rect 3056 26182 3108 26188
rect 2594 26072 2650 26081
rect 2594 26007 2650 26016
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 2582 25596 2890 25616
rect 2582 25594 2588 25596
rect 2644 25594 2668 25596
rect 2724 25594 2748 25596
rect 2804 25594 2828 25596
rect 2884 25594 2890 25596
rect 2644 25542 2646 25594
rect 2826 25542 2828 25594
rect 2582 25540 2588 25542
rect 2644 25540 2668 25542
rect 2724 25540 2748 25542
rect 2804 25540 2828 25542
rect 2884 25540 2890 25542
rect 2582 25520 2890 25540
rect 2976 25265 3004 25842
rect 3068 25430 3096 26182
rect 3056 25424 3108 25430
rect 3056 25366 3108 25372
rect 2962 25256 3018 25265
rect 2962 25191 3018 25200
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2884 24721 2912 25094
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2870 24712 2926 24721
rect 2870 24647 2926 24656
rect 2582 24508 2890 24528
rect 2582 24506 2588 24508
rect 2644 24506 2668 24508
rect 2724 24506 2748 24508
rect 2804 24506 2828 24508
rect 2884 24506 2890 24508
rect 2644 24454 2646 24506
rect 2826 24454 2828 24506
rect 2582 24452 2588 24454
rect 2644 24452 2668 24454
rect 2724 24452 2748 24454
rect 2804 24452 2828 24454
rect 2884 24452 2890 24454
rect 2582 24432 2890 24452
rect 2976 24206 3004 24754
rect 2688 24200 2740 24206
rect 2964 24200 3016 24206
rect 2740 24148 2820 24154
rect 2688 24142 2820 24148
rect 2964 24142 3016 24148
rect 2700 24126 2820 24142
rect 2792 23662 2820 24126
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2582 23420 2890 23440
rect 2582 23418 2588 23420
rect 2644 23418 2668 23420
rect 2724 23418 2748 23420
rect 2804 23418 2828 23420
rect 2884 23418 2890 23420
rect 2644 23366 2646 23418
rect 2826 23366 2828 23418
rect 2582 23364 2588 23366
rect 2644 23364 2668 23366
rect 2724 23364 2748 23366
rect 2804 23364 2828 23366
rect 2884 23364 2890 23366
rect 2582 23344 2890 23364
rect 2976 22574 3004 24142
rect 3056 24132 3108 24138
rect 3056 24074 3108 24080
rect 3068 23866 3096 24074
rect 3056 23860 3108 23866
rect 3056 23802 3108 23808
rect 3056 23724 3108 23730
rect 3056 23666 3108 23672
rect 3068 23186 3096 23666
rect 3056 23180 3108 23186
rect 3056 23122 3108 23128
rect 3068 22778 3096 23122
rect 3056 22772 3108 22778
rect 3056 22714 3108 22720
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 2582 22332 2890 22352
rect 2582 22330 2588 22332
rect 2644 22330 2668 22332
rect 2724 22330 2748 22332
rect 2804 22330 2828 22332
rect 2884 22330 2890 22332
rect 2644 22278 2646 22330
rect 2826 22278 2828 22330
rect 2582 22276 2588 22278
rect 2644 22276 2668 22278
rect 2724 22276 2748 22278
rect 2804 22276 2828 22278
rect 2884 22276 2890 22278
rect 2582 22256 2890 22276
rect 2582 21244 2890 21264
rect 2582 21242 2588 21244
rect 2644 21242 2668 21244
rect 2724 21242 2748 21244
rect 2804 21242 2828 21244
rect 2884 21242 2890 21244
rect 2644 21190 2646 21242
rect 2826 21190 2828 21242
rect 2582 21188 2588 21190
rect 2644 21188 2668 21190
rect 2724 21188 2748 21190
rect 2804 21188 2828 21190
rect 2884 21188 2890 21190
rect 2582 21168 2890 21188
rect 2976 20942 3004 22510
rect 3056 22500 3108 22506
rect 3056 22442 3108 22448
rect 3068 22030 3096 22442
rect 3160 22438 3188 26279
rect 3252 25650 3280 29582
rect 3344 27538 3372 31447
rect 3332 27532 3384 27538
rect 3332 27474 3384 27480
rect 3330 27432 3386 27441
rect 3330 27367 3386 27376
rect 3344 26246 3372 27367
rect 3332 26240 3384 26246
rect 3332 26182 3384 26188
rect 3436 26042 3464 31894
rect 3424 26036 3476 26042
rect 3424 25978 3476 25984
rect 3332 25900 3384 25906
rect 3332 25842 3384 25848
rect 3344 25809 3372 25842
rect 3330 25800 3386 25809
rect 3330 25735 3386 25744
rect 3252 25622 3464 25650
rect 3240 24744 3292 24750
rect 3240 24686 3292 24692
rect 3252 23526 3280 24686
rect 3332 23656 3384 23662
rect 3332 23598 3384 23604
rect 3240 23520 3292 23526
rect 3240 23462 3292 23468
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 3148 22432 3200 22438
rect 3148 22374 3200 22380
rect 3148 22228 3200 22234
rect 3148 22170 3200 22176
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 2964 20936 3016 20942
rect 2964 20878 3016 20884
rect 2778 20632 2834 20641
rect 2778 20567 2834 20576
rect 2792 20466 2820 20567
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 2582 20156 2890 20176
rect 2582 20154 2588 20156
rect 2644 20154 2668 20156
rect 2724 20154 2748 20156
rect 2804 20154 2828 20156
rect 2884 20154 2890 20156
rect 2644 20102 2646 20154
rect 2826 20102 2828 20154
rect 2582 20100 2588 20102
rect 2644 20100 2668 20102
rect 2724 20100 2748 20102
rect 2804 20100 2828 20102
rect 2884 20100 2890 20102
rect 2582 20080 2890 20100
rect 3068 20058 3096 21490
rect 3160 20466 3188 22170
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3252 19854 3280 22714
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 2582 19068 2890 19088
rect 2582 19066 2588 19068
rect 2644 19066 2668 19068
rect 2724 19066 2748 19068
rect 2804 19066 2828 19068
rect 2884 19066 2890 19068
rect 2644 19014 2646 19066
rect 2826 19014 2828 19066
rect 2582 19012 2588 19014
rect 2644 19012 2668 19014
rect 2724 19012 2748 19014
rect 2804 19012 2828 19014
rect 2884 19012 2890 19014
rect 2582 18992 2890 19012
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2792 18442 2820 18770
rect 2700 18414 2820 18442
rect 2976 18426 3004 19314
rect 3252 18834 3280 19790
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 2964 18420 3016 18426
rect 2700 18290 2728 18414
rect 2964 18362 3016 18368
rect 3148 18352 3200 18358
rect 3148 18294 3200 18300
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2332 18006 2452 18034
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2136 15904 2188 15910
rect 2136 15846 2188 15852
rect 2056 15570 2084 15846
rect 2148 15706 2176 15846
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 2240 15473 2268 16050
rect 2226 15464 2282 15473
rect 2226 15399 2282 15408
rect 2136 15360 2188 15366
rect 2332 15314 2360 18006
rect 2516 17678 2544 18090
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2582 17980 2890 18000
rect 2582 17978 2588 17980
rect 2644 17978 2668 17980
rect 2724 17978 2748 17980
rect 2804 17978 2828 17980
rect 2884 17978 2890 17980
rect 2644 17926 2646 17978
rect 2826 17926 2828 17978
rect 2582 17924 2588 17926
rect 2644 17924 2668 17926
rect 2724 17924 2748 17926
rect 2804 17924 2828 17926
rect 2884 17924 2890 17926
rect 2582 17904 2890 17924
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2410 17232 2466 17241
rect 2410 17167 2466 17176
rect 2424 16590 2452 17167
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2136 15302 2188 15308
rect 2148 14482 2176 15302
rect 2240 15286 2360 15314
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 1964 14334 2176 14362
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1964 10674 1992 14214
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 2056 9042 2084 13398
rect 2148 12238 2176 14334
rect 2240 14006 2268 15286
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2148 7410 2176 11154
rect 2240 7954 2268 13262
rect 2332 12986 2360 14350
rect 2424 13818 2452 15302
rect 2516 14618 2544 17614
rect 2976 17202 3004 18022
rect 3068 17746 3096 18158
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 3160 17678 3188 18294
rect 3148 17672 3200 17678
rect 3054 17640 3110 17649
rect 3148 17614 3200 17620
rect 3054 17575 3110 17584
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2582 16892 2890 16912
rect 2582 16890 2588 16892
rect 2644 16890 2668 16892
rect 2724 16890 2748 16892
rect 2804 16890 2828 16892
rect 2884 16890 2890 16892
rect 2644 16838 2646 16890
rect 2826 16838 2828 16890
rect 2582 16836 2588 16838
rect 2644 16836 2668 16838
rect 2724 16836 2748 16838
rect 2804 16836 2828 16838
rect 2884 16836 2890 16838
rect 2582 16816 2890 16836
rect 3068 16590 3096 17575
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2884 16017 2912 16050
rect 2870 16008 2926 16017
rect 2870 15943 2926 15952
rect 2582 15804 2890 15824
rect 2582 15802 2588 15804
rect 2644 15802 2668 15804
rect 2724 15802 2748 15804
rect 2804 15802 2828 15804
rect 2884 15802 2890 15804
rect 2644 15750 2646 15802
rect 2826 15750 2828 15802
rect 2582 15748 2588 15750
rect 2644 15748 2668 15750
rect 2724 15748 2748 15750
rect 2804 15748 2828 15750
rect 2884 15748 2890 15750
rect 2582 15728 2890 15748
rect 3056 15088 3108 15094
rect 3056 15030 3108 15036
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 2582 14716 2890 14736
rect 2582 14714 2588 14716
rect 2644 14714 2668 14716
rect 2724 14714 2748 14716
rect 2804 14714 2828 14716
rect 2884 14714 2890 14716
rect 2644 14662 2646 14714
rect 2826 14662 2828 14714
rect 2582 14660 2588 14662
rect 2644 14660 2668 14662
rect 2724 14660 2748 14662
rect 2804 14660 2828 14662
rect 2884 14660 2890 14662
rect 2582 14640 2890 14660
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2976 13841 3004 14962
rect 2962 13832 3018 13841
rect 2424 13790 2544 13818
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2424 13190 2452 13670
rect 2516 13462 2544 13790
rect 2962 13767 3018 13776
rect 3068 13716 3096 15030
rect 2976 13688 3096 13716
rect 2582 13628 2890 13648
rect 2582 13626 2588 13628
rect 2644 13626 2668 13628
rect 2724 13626 2748 13628
rect 2804 13626 2828 13628
rect 2884 13626 2890 13628
rect 2644 13574 2646 13626
rect 2826 13574 2828 13626
rect 2582 13572 2588 13574
rect 2644 13572 2668 13574
rect 2724 13572 2748 13574
rect 2804 13572 2828 13574
rect 2884 13572 2890 13574
rect 2582 13552 2890 13572
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2424 8498 2452 13126
rect 2976 12866 3004 13688
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3068 12986 3096 13466
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2976 12838 3096 12866
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2582 12540 2890 12560
rect 2582 12538 2588 12540
rect 2644 12538 2668 12540
rect 2724 12538 2748 12540
rect 2804 12538 2828 12540
rect 2884 12538 2890 12540
rect 2644 12486 2646 12538
rect 2826 12486 2828 12538
rect 2582 12484 2588 12486
rect 2644 12484 2668 12486
rect 2724 12484 2748 12486
rect 2804 12484 2828 12486
rect 2884 12484 2890 12486
rect 2582 12464 2890 12484
rect 2976 11626 3004 12650
rect 3068 11898 3096 12838
rect 3160 12714 3188 17614
rect 3252 17134 3280 18634
rect 3240 17128 3292 17134
rect 3238 17096 3240 17105
rect 3292 17096 3294 17105
rect 3238 17031 3294 17040
rect 3344 16522 3372 23598
rect 3436 21146 3464 25622
rect 3528 22778 3556 32150
rect 3620 31346 3648 41103
rect 3698 41032 3754 41041
rect 3698 40967 3754 40976
rect 3712 39030 3740 40967
rect 3700 39024 3752 39030
rect 3700 38966 3752 38972
rect 3700 38752 3752 38758
rect 3700 38694 3752 38700
rect 3712 38457 3740 38694
rect 3698 38448 3754 38457
rect 3698 38383 3754 38392
rect 3700 38344 3752 38350
rect 3700 38286 3752 38292
rect 3712 35873 3740 38286
rect 3804 37262 3832 43046
rect 3896 40594 3924 48311
rect 3988 47462 4016 48504
rect 3976 47456 4028 47462
rect 3976 47398 4028 47404
rect 3976 47184 4028 47190
rect 3976 47126 4028 47132
rect 3988 47025 4016 47126
rect 3974 47016 4030 47025
rect 3974 46951 4030 46960
rect 4080 46866 4108 48690
rect 4356 48278 4384 48844
rect 4528 48612 4580 48618
rect 4528 48554 4580 48560
rect 4344 48272 4396 48278
rect 4344 48214 4396 48220
rect 4540 48210 4568 48554
rect 4528 48204 4580 48210
rect 4528 48146 4580 48152
rect 4214 47900 4522 47920
rect 4214 47898 4220 47900
rect 4276 47898 4300 47900
rect 4356 47898 4380 47900
rect 4436 47898 4460 47900
rect 4516 47898 4522 47900
rect 4276 47846 4278 47898
rect 4458 47846 4460 47898
rect 4214 47844 4220 47846
rect 4276 47844 4300 47846
rect 4356 47844 4380 47846
rect 4436 47844 4460 47846
rect 4516 47844 4522 47846
rect 4214 47824 4522 47844
rect 4436 47184 4488 47190
rect 4436 47126 4488 47132
rect 4448 47054 4476 47126
rect 4436 47048 4488 47054
rect 4250 47016 4306 47025
rect 4436 46990 4488 46996
rect 4250 46951 4252 46960
rect 4304 46951 4306 46960
rect 4252 46922 4304 46928
rect 3988 46838 4108 46866
rect 3988 45778 4016 46838
rect 4214 46812 4522 46832
rect 4214 46810 4220 46812
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4516 46810 4522 46812
rect 4276 46758 4278 46810
rect 4458 46758 4460 46810
rect 4214 46756 4220 46758
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4516 46756 4522 46758
rect 4214 46736 4522 46756
rect 4068 46504 4120 46510
rect 4068 46446 4120 46452
rect 4080 45898 4108 46446
rect 4528 46368 4580 46374
rect 4528 46310 4580 46316
rect 4540 45898 4568 46310
rect 4068 45892 4120 45898
rect 4068 45834 4120 45840
rect 4528 45892 4580 45898
rect 4528 45834 4580 45840
rect 3988 45750 4108 45778
rect 3974 45656 4030 45665
rect 3974 45591 4030 45600
rect 3988 43994 4016 45591
rect 3976 43988 4028 43994
rect 3976 43930 4028 43936
rect 3976 43648 4028 43654
rect 3974 43616 3976 43625
rect 4028 43616 4030 43625
rect 3974 43551 4030 43560
rect 3974 43208 4030 43217
rect 3974 43143 3976 43152
rect 4028 43143 4030 43152
rect 3976 43114 4028 43120
rect 3974 42664 4030 42673
rect 3974 42599 4030 42608
rect 3988 42566 4016 42599
rect 3976 42560 4028 42566
rect 3976 42502 4028 42508
rect 3976 42356 4028 42362
rect 3976 42298 4028 42304
rect 3884 40588 3936 40594
rect 3884 40530 3936 40536
rect 3988 40474 4016 42298
rect 3896 40446 4016 40474
rect 3792 37256 3844 37262
rect 3792 37198 3844 37204
rect 3792 36916 3844 36922
rect 3792 36858 3844 36864
rect 3804 36281 3832 36858
rect 3790 36272 3846 36281
rect 3790 36207 3846 36216
rect 3896 36122 3924 40446
rect 3976 40384 4028 40390
rect 3976 40326 4028 40332
rect 3988 40225 4016 40326
rect 3974 40216 4030 40225
rect 3974 40151 4030 40160
rect 3976 39840 4028 39846
rect 3976 39782 4028 39788
rect 3988 39545 4016 39782
rect 3974 39536 4030 39545
rect 3974 39471 4030 39480
rect 4080 39438 4108 45750
rect 4214 45724 4522 45744
rect 4214 45722 4220 45724
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4516 45722 4522 45724
rect 4276 45670 4278 45722
rect 4458 45670 4460 45722
rect 4214 45668 4220 45670
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4516 45668 4522 45670
rect 4214 45648 4522 45668
rect 4160 45416 4212 45422
rect 4160 45358 4212 45364
rect 4172 44849 4200 45358
rect 4158 44840 4214 44849
rect 4158 44775 4214 44784
rect 4214 44636 4522 44656
rect 4214 44634 4220 44636
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4516 44634 4522 44636
rect 4276 44582 4278 44634
rect 4458 44582 4460 44634
rect 4214 44580 4220 44582
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4516 44580 4522 44582
rect 4214 44560 4522 44580
rect 4214 43548 4522 43568
rect 4214 43546 4220 43548
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4516 43546 4522 43548
rect 4276 43494 4278 43546
rect 4458 43494 4460 43546
rect 4214 43492 4220 43494
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4516 43492 4522 43494
rect 4214 43472 4522 43492
rect 4158 43344 4214 43353
rect 4158 43279 4214 43288
rect 4172 42702 4200 43279
rect 4160 42696 4212 42702
rect 4160 42638 4212 42644
rect 4214 42460 4522 42480
rect 4214 42458 4220 42460
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4516 42458 4522 42460
rect 4276 42406 4278 42458
rect 4458 42406 4460 42458
rect 4214 42404 4220 42406
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4516 42404 4522 42406
rect 4214 42384 4522 42404
rect 4436 42288 4488 42294
rect 4436 42230 4488 42236
rect 4448 41585 4476 42230
rect 4434 41576 4490 41585
rect 4434 41511 4490 41520
rect 4214 41372 4522 41392
rect 4214 41370 4220 41372
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4516 41370 4522 41372
rect 4276 41318 4278 41370
rect 4458 41318 4460 41370
rect 4214 41316 4220 41318
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4516 41316 4522 41318
rect 4214 41296 4522 41316
rect 4436 41064 4488 41070
rect 4436 41006 4488 41012
rect 4448 40662 4476 41006
rect 4436 40656 4488 40662
rect 4436 40598 4488 40604
rect 4214 40284 4522 40304
rect 4214 40282 4220 40284
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4516 40282 4522 40284
rect 4276 40230 4278 40282
rect 4458 40230 4460 40282
rect 4214 40228 4220 40230
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4516 40228 4522 40230
rect 4214 40208 4522 40228
rect 4068 39432 4120 39438
rect 4068 39374 4120 39380
rect 3976 39296 4028 39302
rect 3974 39264 3976 39273
rect 4028 39264 4030 39273
rect 3974 39199 4030 39208
rect 4214 39196 4522 39216
rect 4214 39194 4220 39196
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4516 39194 4522 39196
rect 4276 39142 4278 39194
rect 4458 39142 4460 39194
rect 4214 39140 4220 39142
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4516 39140 4522 39142
rect 4214 39120 4522 39140
rect 4632 39080 4660 55694
rect 4724 50522 4752 55950
rect 4802 55856 4858 55865
rect 4802 55791 4858 55800
rect 4712 50516 4764 50522
rect 4712 50458 4764 50464
rect 4712 50380 4764 50386
rect 4712 50322 4764 50328
rect 4724 46374 4752 50322
rect 4712 46368 4764 46374
rect 4712 46310 4764 46316
rect 4712 46164 4764 46170
rect 4712 46106 4764 46112
rect 4540 39052 4660 39080
rect 4436 39024 4488 39030
rect 4158 38992 4214 39001
rect 4436 38966 4488 38972
rect 4158 38927 4214 38936
rect 3974 38856 4030 38865
rect 3974 38791 4030 38800
rect 3988 37777 4016 38791
rect 4172 38654 4200 38927
rect 4344 38888 4396 38894
rect 4344 38830 4396 38836
rect 4252 38820 4304 38826
rect 4252 38762 4304 38768
rect 4080 38626 4200 38654
rect 3974 37768 4030 37777
rect 3974 37703 4030 37712
rect 3974 37224 4030 37233
rect 3974 37159 4030 37168
rect 3988 37126 4016 37159
rect 3976 37120 4028 37126
rect 3976 37062 4028 37068
rect 4080 36904 4108 38626
rect 4264 38350 4292 38762
rect 4252 38344 4304 38350
rect 4356 38321 4384 38830
rect 4448 38418 4476 38966
rect 4540 38826 4568 39052
rect 4724 38962 4752 46106
rect 4816 42294 4844 55791
rect 4908 46170 4936 68954
rect 7478 68572 7786 68592
rect 7478 68570 7484 68572
rect 7540 68570 7564 68572
rect 7620 68570 7644 68572
rect 7700 68570 7724 68572
rect 7780 68570 7786 68572
rect 7540 68518 7542 68570
rect 7722 68518 7724 68570
rect 7478 68516 7484 68518
rect 7540 68516 7564 68518
rect 7620 68516 7644 68518
rect 7700 68516 7724 68518
rect 7780 68516 7786 68518
rect 7478 68496 7786 68516
rect 5846 68028 6154 68048
rect 5846 68026 5852 68028
rect 5908 68026 5932 68028
rect 5988 68026 6012 68028
rect 6068 68026 6092 68028
rect 6148 68026 6154 68028
rect 5908 67974 5910 68026
rect 6090 67974 6092 68026
rect 5846 67972 5852 67974
rect 5908 67972 5932 67974
rect 5988 67972 6012 67974
rect 6068 67972 6092 67974
rect 6148 67972 6154 67974
rect 5846 67952 6154 67972
rect 9110 68028 9418 68048
rect 9110 68026 9116 68028
rect 9172 68026 9196 68028
rect 9252 68026 9276 68028
rect 9332 68026 9356 68028
rect 9412 68026 9418 68028
rect 9172 67974 9174 68026
rect 9354 67974 9356 68026
rect 9110 67972 9116 67974
rect 9172 67972 9196 67974
rect 9252 67972 9276 67974
rect 9332 67972 9356 67974
rect 9412 67972 9418 67974
rect 9110 67952 9418 67972
rect 7478 67484 7786 67504
rect 7478 67482 7484 67484
rect 7540 67482 7564 67484
rect 7620 67482 7644 67484
rect 7700 67482 7724 67484
rect 7780 67482 7786 67484
rect 7540 67430 7542 67482
rect 7722 67430 7724 67482
rect 7478 67428 7484 67430
rect 7540 67428 7564 67430
rect 7620 67428 7644 67430
rect 7700 67428 7724 67430
rect 7780 67428 7786 67430
rect 7478 67408 7786 67428
rect 9680 67380 9732 67386
rect 9680 67322 9732 67328
rect 8484 67040 8536 67046
rect 8484 66982 8536 66988
rect 5846 66940 6154 66960
rect 5846 66938 5852 66940
rect 5908 66938 5932 66940
rect 5988 66938 6012 66940
rect 6068 66938 6092 66940
rect 6148 66938 6154 66940
rect 5908 66886 5910 66938
rect 6090 66886 6092 66938
rect 5846 66884 5852 66886
rect 5908 66884 5932 66886
rect 5988 66884 6012 66886
rect 6068 66884 6092 66886
rect 6148 66884 6154 66886
rect 5846 66864 6154 66884
rect 7478 66396 7786 66416
rect 7478 66394 7484 66396
rect 7540 66394 7564 66396
rect 7620 66394 7644 66396
rect 7700 66394 7724 66396
rect 7780 66394 7786 66396
rect 7540 66342 7542 66394
rect 7722 66342 7724 66394
rect 7478 66340 7484 66342
rect 7540 66340 7564 66342
rect 7620 66340 7644 66342
rect 7700 66340 7724 66342
rect 7780 66340 7786 66342
rect 7478 66320 7786 66340
rect 8300 65952 8352 65958
rect 8300 65894 8352 65900
rect 5846 65852 6154 65872
rect 5846 65850 5852 65852
rect 5908 65850 5932 65852
rect 5988 65850 6012 65852
rect 6068 65850 6092 65852
rect 6148 65850 6154 65852
rect 5908 65798 5910 65850
rect 6090 65798 6092 65850
rect 5846 65796 5852 65798
rect 5908 65796 5932 65798
rect 5988 65796 6012 65798
rect 6068 65796 6092 65798
rect 6148 65796 6154 65798
rect 5846 65776 6154 65796
rect 4988 65680 5040 65686
rect 4988 65622 5040 65628
rect 5000 63034 5028 65622
rect 7478 65308 7786 65328
rect 7478 65306 7484 65308
rect 7540 65306 7564 65308
rect 7620 65306 7644 65308
rect 7700 65306 7724 65308
rect 7780 65306 7786 65308
rect 7540 65254 7542 65306
rect 7722 65254 7724 65306
rect 7478 65252 7484 65254
rect 7540 65252 7564 65254
rect 7620 65252 7644 65254
rect 7700 65252 7724 65254
rect 7780 65252 7786 65254
rect 7478 65232 7786 65252
rect 5846 64764 6154 64784
rect 5846 64762 5852 64764
rect 5908 64762 5932 64764
rect 5988 64762 6012 64764
rect 6068 64762 6092 64764
rect 6148 64762 6154 64764
rect 5908 64710 5910 64762
rect 6090 64710 6092 64762
rect 5846 64708 5852 64710
rect 5908 64708 5932 64710
rect 5988 64708 6012 64710
rect 6068 64708 6092 64710
rect 6148 64708 6154 64710
rect 5846 64688 6154 64708
rect 8312 64666 8340 65894
rect 8392 64932 8444 64938
rect 8392 64874 8444 64880
rect 8300 64660 8352 64666
rect 8300 64602 8352 64608
rect 8300 64320 8352 64326
rect 8300 64262 8352 64268
rect 7478 64220 7786 64240
rect 7478 64218 7484 64220
rect 7540 64218 7564 64220
rect 7620 64218 7644 64220
rect 7700 64218 7724 64220
rect 7780 64218 7786 64220
rect 7540 64166 7542 64218
rect 7722 64166 7724 64218
rect 7478 64164 7484 64166
rect 7540 64164 7564 64166
rect 7620 64164 7644 64166
rect 7700 64164 7724 64166
rect 7780 64164 7786 64166
rect 7478 64144 7786 64164
rect 5172 63776 5224 63782
rect 5172 63718 5224 63724
rect 4988 63028 5040 63034
rect 4988 62970 5040 62976
rect 5080 59016 5132 59022
rect 5080 58958 5132 58964
rect 4988 56432 5040 56438
rect 4988 56374 5040 56380
rect 5000 50386 5028 56374
rect 5092 53145 5120 58958
rect 5078 53136 5134 53145
rect 5078 53071 5134 53080
rect 5080 52964 5132 52970
rect 5080 52906 5132 52912
rect 5092 51241 5120 52906
rect 5078 51232 5134 51241
rect 5078 51167 5134 51176
rect 5078 51096 5134 51105
rect 5184 51066 5212 63718
rect 5846 63676 6154 63696
rect 5846 63674 5852 63676
rect 5908 63674 5932 63676
rect 5988 63674 6012 63676
rect 6068 63674 6092 63676
rect 6148 63674 6154 63676
rect 5908 63622 5910 63674
rect 6090 63622 6092 63674
rect 5846 63620 5852 63622
rect 5908 63620 5932 63622
rect 5988 63620 6012 63622
rect 6068 63620 6092 63622
rect 6148 63620 6154 63622
rect 5846 63600 6154 63620
rect 8312 63510 8340 64262
rect 8404 63918 8432 64874
rect 8392 63912 8444 63918
rect 8392 63854 8444 63860
rect 8300 63504 8352 63510
rect 8300 63446 8352 63452
rect 7478 63132 7786 63152
rect 7478 63130 7484 63132
rect 7540 63130 7564 63132
rect 7620 63130 7644 63132
rect 7700 63130 7724 63132
rect 7780 63130 7786 63132
rect 7540 63078 7542 63130
rect 7722 63078 7724 63130
rect 7478 63076 7484 63078
rect 7540 63076 7564 63078
rect 7620 63076 7644 63078
rect 7700 63076 7724 63078
rect 7780 63076 7786 63078
rect 7478 63056 7786 63076
rect 5356 62892 5408 62898
rect 5356 62834 5408 62840
rect 5264 62688 5316 62694
rect 5264 62630 5316 62636
rect 5078 51031 5134 51040
rect 5172 51060 5224 51066
rect 4988 50380 5040 50386
rect 4988 50322 5040 50328
rect 4986 50280 5042 50289
rect 4986 50215 5042 50224
rect 4896 46164 4948 46170
rect 4896 46106 4948 46112
rect 5000 46050 5028 50215
rect 4908 46022 5028 46050
rect 4804 42288 4856 42294
rect 4804 42230 4856 42236
rect 4802 42120 4858 42129
rect 4802 42055 4858 42064
rect 4712 38956 4764 38962
rect 4712 38898 4764 38904
rect 4528 38820 4580 38826
rect 4528 38762 4580 38768
rect 4712 38820 4764 38826
rect 4712 38762 4764 38768
rect 4620 38752 4672 38758
rect 4620 38694 4672 38700
rect 4436 38412 4488 38418
rect 4436 38354 4488 38360
rect 4252 38286 4304 38292
rect 4342 38312 4398 38321
rect 4342 38247 4398 38256
rect 4214 38108 4522 38128
rect 4214 38106 4220 38108
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4516 38106 4522 38108
rect 4276 38054 4278 38106
rect 4458 38054 4460 38106
rect 4214 38052 4220 38054
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4516 38052 4522 38054
rect 4214 38032 4522 38052
rect 4214 37020 4522 37040
rect 4214 37018 4220 37020
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4516 37018 4522 37020
rect 4276 36966 4278 37018
rect 4458 36966 4460 37018
rect 4214 36964 4220 36966
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4516 36964 4522 36966
rect 4214 36944 4522 36964
rect 4080 36876 4200 36904
rect 3974 36680 4030 36689
rect 3974 36615 4030 36624
rect 4068 36644 4120 36650
rect 3988 36378 4016 36615
rect 4068 36586 4120 36592
rect 3976 36372 4028 36378
rect 3976 36314 4028 36320
rect 4080 36258 4108 36586
rect 3804 36094 3924 36122
rect 3988 36230 4108 36258
rect 3698 35864 3754 35873
rect 3698 35799 3754 35808
rect 3700 33040 3752 33046
rect 3700 32982 3752 32988
rect 3712 32881 3740 32982
rect 3698 32872 3754 32881
rect 3698 32807 3754 32816
rect 3700 32428 3752 32434
rect 3700 32370 3752 32376
rect 3608 31340 3660 31346
rect 3608 31282 3660 31288
rect 3606 31240 3662 31249
rect 3606 31175 3608 31184
rect 3660 31175 3662 31184
rect 3608 31146 3660 31152
rect 3606 30696 3662 30705
rect 3606 30631 3662 30640
rect 3620 25974 3648 30631
rect 3608 25968 3660 25974
rect 3608 25910 3660 25916
rect 3606 25800 3662 25809
rect 3606 25735 3662 25744
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3528 22545 3556 22578
rect 3514 22536 3570 22545
rect 3514 22471 3570 22480
rect 3620 22234 3648 25735
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3424 20936 3476 20942
rect 3424 20878 3476 20884
rect 3332 16516 3384 16522
rect 3332 16458 3384 16464
rect 3240 16448 3292 16454
rect 3240 16390 3292 16396
rect 3252 15502 3280 16390
rect 3436 15745 3464 20878
rect 3608 19440 3660 19446
rect 3608 19382 3660 19388
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3528 17610 3556 19314
rect 3620 17882 3648 19382
rect 3712 18442 3740 32370
rect 3804 25498 3832 36094
rect 3988 35986 4016 36230
rect 4172 36145 4200 36876
rect 4632 36650 4660 38694
rect 4620 36644 4672 36650
rect 4620 36586 4672 36592
rect 4724 36530 4752 38762
rect 4632 36502 4752 36530
rect 4158 36136 4214 36145
rect 4158 36071 4214 36080
rect 3896 35958 4016 35986
rect 3896 31958 3924 35958
rect 4214 35932 4522 35952
rect 4214 35930 4220 35932
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4516 35930 4522 35932
rect 4276 35878 4278 35930
rect 4458 35878 4460 35930
rect 4214 35876 4220 35878
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4516 35876 4522 35878
rect 3974 35864 4030 35873
rect 4214 35856 4522 35876
rect 3974 35799 4030 35808
rect 3988 35698 4016 35799
rect 4632 35714 4660 36502
rect 4712 36168 4764 36174
rect 4712 36110 4764 36116
rect 4724 35834 4752 36110
rect 4712 35828 4764 35834
rect 4712 35770 4764 35776
rect 3976 35692 4028 35698
rect 4632 35686 4752 35714
rect 3976 35634 4028 35640
rect 3988 34592 4016 35634
rect 4620 35624 4672 35630
rect 4620 35566 4672 35572
rect 4068 35080 4120 35086
rect 4068 35022 4120 35028
rect 4080 34746 4108 35022
rect 4214 34844 4522 34864
rect 4214 34842 4220 34844
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4516 34842 4522 34844
rect 4276 34790 4278 34842
rect 4458 34790 4460 34842
rect 4214 34788 4220 34790
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4516 34788 4522 34790
rect 4214 34768 4522 34788
rect 4068 34740 4120 34746
rect 4068 34682 4120 34688
rect 3988 34564 4108 34592
rect 3976 34468 4028 34474
rect 3976 34410 4028 34416
rect 3988 33658 4016 34410
rect 3976 33652 4028 33658
rect 3976 33594 4028 33600
rect 3976 32768 4028 32774
rect 3976 32710 4028 32716
rect 3988 32473 4016 32710
rect 3974 32464 4030 32473
rect 3974 32399 4030 32408
rect 3976 32224 4028 32230
rect 3976 32166 4028 32172
rect 3884 31952 3936 31958
rect 3988 31929 4016 32166
rect 3884 31894 3936 31900
rect 3974 31920 4030 31929
rect 3974 31855 4030 31864
rect 3882 31784 3938 31793
rect 3882 31719 3938 31728
rect 3896 31634 3924 31719
rect 3896 31606 4016 31634
rect 3882 31512 3938 31521
rect 3882 31447 3938 31456
rect 3896 29238 3924 31447
rect 3988 30977 4016 31606
rect 3974 30968 4030 30977
rect 3974 30903 4030 30912
rect 4080 30818 4108 34564
rect 4214 33756 4522 33776
rect 4214 33754 4220 33756
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4516 33754 4522 33756
rect 4276 33702 4278 33754
rect 4458 33702 4460 33754
rect 4214 33700 4220 33702
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4516 33700 4522 33702
rect 4214 33680 4522 33700
rect 4632 33572 4660 35566
rect 4540 33544 4660 33572
rect 4540 33017 4568 33544
rect 4620 33448 4672 33454
rect 4620 33390 4672 33396
rect 4526 33008 4582 33017
rect 4526 32943 4582 32952
rect 4214 32668 4522 32688
rect 4214 32666 4220 32668
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4516 32666 4522 32668
rect 4276 32614 4278 32666
rect 4458 32614 4460 32666
rect 4214 32612 4220 32614
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4516 32612 4522 32614
rect 4214 32592 4522 32612
rect 4436 32496 4488 32502
rect 4436 32438 4488 32444
rect 4526 32464 4582 32473
rect 4448 31890 4476 32438
rect 4526 32399 4582 32408
rect 4436 31884 4488 31890
rect 4436 31826 4488 31832
rect 4540 31668 4568 32399
rect 4632 32026 4660 33390
rect 4724 32065 4752 35686
rect 4816 32502 4844 42055
rect 4804 32496 4856 32502
rect 4804 32438 4856 32444
rect 4710 32056 4766 32065
rect 4620 32020 4672 32026
rect 4908 32026 4936 46022
rect 4988 45892 5040 45898
rect 4988 45834 5040 45840
rect 5000 40934 5028 45834
rect 5092 41585 5120 51031
rect 5172 51002 5224 51008
rect 5276 50998 5304 62630
rect 5368 53174 5396 62834
rect 5846 62588 6154 62608
rect 5846 62586 5852 62588
rect 5908 62586 5932 62588
rect 5988 62586 6012 62588
rect 6068 62586 6092 62588
rect 6148 62586 6154 62588
rect 5908 62534 5910 62586
rect 6090 62534 6092 62586
rect 5846 62532 5852 62534
rect 5908 62532 5932 62534
rect 5988 62532 6012 62534
rect 6068 62532 6092 62534
rect 6148 62532 6154 62534
rect 5846 62512 6154 62532
rect 8300 62144 8352 62150
rect 8300 62086 8352 62092
rect 7478 62044 7786 62064
rect 7478 62042 7484 62044
rect 7540 62042 7564 62044
rect 7620 62042 7644 62044
rect 7700 62042 7724 62044
rect 7780 62042 7786 62044
rect 7540 61990 7542 62042
rect 7722 61990 7724 62042
rect 7478 61988 7484 61990
rect 7540 61988 7564 61990
rect 7620 61988 7644 61990
rect 7700 61988 7724 61990
rect 7780 61988 7786 61990
rect 7478 61968 7786 61988
rect 8312 61878 8340 62086
rect 8300 61872 8352 61878
rect 8300 61814 8352 61820
rect 5846 61500 6154 61520
rect 5846 61498 5852 61500
rect 5908 61498 5932 61500
rect 5988 61498 6012 61500
rect 6068 61498 6092 61500
rect 6148 61498 6154 61500
rect 5908 61446 5910 61498
rect 6090 61446 6092 61498
rect 5846 61444 5852 61446
rect 5908 61444 5932 61446
rect 5988 61444 6012 61446
rect 6068 61444 6092 61446
rect 6148 61444 6154 61446
rect 5846 61424 6154 61444
rect 7478 60956 7786 60976
rect 7478 60954 7484 60956
rect 7540 60954 7564 60956
rect 7620 60954 7644 60956
rect 7700 60954 7724 60956
rect 7780 60954 7786 60956
rect 7540 60902 7542 60954
rect 7722 60902 7724 60954
rect 7478 60900 7484 60902
rect 7540 60900 7564 60902
rect 7620 60900 7644 60902
rect 7700 60900 7724 60902
rect 7780 60900 7786 60902
rect 7478 60880 7786 60900
rect 6920 60512 6972 60518
rect 6920 60454 6972 60460
rect 5846 60412 6154 60432
rect 5846 60410 5852 60412
rect 5908 60410 5932 60412
rect 5988 60410 6012 60412
rect 6068 60410 6092 60412
rect 6148 60410 6154 60412
rect 5908 60358 5910 60410
rect 6090 60358 6092 60410
rect 5846 60356 5852 60358
rect 5908 60356 5932 60358
rect 5988 60356 6012 60358
rect 6068 60356 6092 60358
rect 6148 60356 6154 60358
rect 5846 60336 6154 60356
rect 5846 59324 6154 59344
rect 5846 59322 5852 59324
rect 5908 59322 5932 59324
rect 5988 59322 6012 59324
rect 6068 59322 6092 59324
rect 6148 59322 6154 59324
rect 5908 59270 5910 59322
rect 6090 59270 6092 59322
rect 5846 59268 5852 59270
rect 5908 59268 5932 59270
rect 5988 59268 6012 59270
rect 6068 59268 6092 59270
rect 6148 59268 6154 59270
rect 5846 59248 6154 59268
rect 5846 58236 6154 58256
rect 5846 58234 5852 58236
rect 5908 58234 5932 58236
rect 5988 58234 6012 58236
rect 6068 58234 6092 58236
rect 6148 58234 6154 58236
rect 5908 58182 5910 58234
rect 6090 58182 6092 58234
rect 5846 58180 5852 58182
rect 5908 58180 5932 58182
rect 5988 58180 6012 58182
rect 6068 58180 6092 58182
rect 6148 58180 6154 58182
rect 5846 58160 6154 58180
rect 6932 57497 6960 60454
rect 7478 59868 7786 59888
rect 7478 59866 7484 59868
rect 7540 59866 7564 59868
rect 7620 59866 7644 59868
rect 7700 59866 7724 59868
rect 7780 59866 7786 59868
rect 7540 59814 7542 59866
rect 7722 59814 7724 59866
rect 7478 59812 7484 59814
rect 7540 59812 7564 59814
rect 7620 59812 7644 59814
rect 7700 59812 7724 59814
rect 7780 59812 7786 59814
rect 7478 59792 7786 59812
rect 8300 59628 8352 59634
rect 8300 59570 8352 59576
rect 7478 58780 7786 58800
rect 7478 58778 7484 58780
rect 7540 58778 7564 58780
rect 7620 58778 7644 58780
rect 7700 58778 7724 58780
rect 7780 58778 7786 58780
rect 7540 58726 7542 58778
rect 7722 58726 7724 58778
rect 7478 58724 7484 58726
rect 7540 58724 7564 58726
rect 7620 58724 7644 58726
rect 7700 58724 7724 58726
rect 7780 58724 7786 58726
rect 7478 58704 7786 58724
rect 7478 57692 7786 57712
rect 7478 57690 7484 57692
rect 7540 57690 7564 57692
rect 7620 57690 7644 57692
rect 7700 57690 7724 57692
rect 7780 57690 7786 57692
rect 7540 57638 7542 57690
rect 7722 57638 7724 57690
rect 7478 57636 7484 57638
rect 7540 57636 7564 57638
rect 7620 57636 7644 57638
rect 7700 57636 7724 57638
rect 7780 57636 7786 57638
rect 7478 57616 7786 57636
rect 6918 57488 6974 57497
rect 6918 57423 6974 57432
rect 6276 57316 6328 57322
rect 6276 57258 6328 57264
rect 5846 57148 6154 57168
rect 5846 57146 5852 57148
rect 5908 57146 5932 57148
rect 5988 57146 6012 57148
rect 6068 57146 6092 57148
rect 6148 57146 6154 57148
rect 5908 57094 5910 57146
rect 6090 57094 6092 57146
rect 5846 57092 5852 57094
rect 5908 57092 5932 57094
rect 5988 57092 6012 57094
rect 6068 57092 6092 57094
rect 6148 57092 6154 57094
rect 5846 57072 6154 57092
rect 5846 56060 6154 56080
rect 5846 56058 5852 56060
rect 5908 56058 5932 56060
rect 5988 56058 6012 56060
rect 6068 56058 6092 56060
rect 6148 56058 6154 56060
rect 5908 56006 5910 56058
rect 6090 56006 6092 56058
rect 5846 56004 5852 56006
rect 5908 56004 5932 56006
rect 5988 56004 6012 56006
rect 6068 56004 6092 56006
rect 6148 56004 6154 56006
rect 5846 55984 6154 56004
rect 5448 55820 5500 55826
rect 5448 55762 5500 55768
rect 5356 53168 5408 53174
rect 5356 53110 5408 53116
rect 5460 51490 5488 55762
rect 5722 55720 5778 55729
rect 5722 55655 5778 55664
rect 5540 55412 5592 55418
rect 5540 55354 5592 55360
rect 5552 54874 5580 55354
rect 5540 54868 5592 54874
rect 5540 54810 5592 54816
rect 5632 52488 5684 52494
rect 5632 52430 5684 52436
rect 5460 51462 5580 51490
rect 5446 51096 5502 51105
rect 5446 51031 5502 51040
rect 5264 50992 5316 50998
rect 5170 50960 5226 50969
rect 5264 50934 5316 50940
rect 5170 50895 5226 50904
rect 5078 41576 5134 41585
rect 5078 41511 5134 41520
rect 5080 41472 5132 41478
rect 5080 41414 5132 41420
rect 4988 40928 5040 40934
rect 4988 40870 5040 40876
rect 4988 40656 5040 40662
rect 4988 40598 5040 40604
rect 5000 36394 5028 40598
rect 5092 36582 5120 41414
rect 5080 36576 5132 36582
rect 5080 36518 5132 36524
rect 5000 36366 5120 36394
rect 4986 36272 5042 36281
rect 4986 36207 5042 36216
rect 4710 31991 4766 32000
rect 4896 32020 4948 32026
rect 4620 31962 4672 31968
rect 4896 31962 4948 31968
rect 5000 31872 5028 36207
rect 4908 31844 5028 31872
rect 4804 31816 4856 31822
rect 4804 31758 4856 31764
rect 4712 31680 4764 31686
rect 4540 31640 4660 31668
rect 4214 31580 4522 31600
rect 4214 31578 4220 31580
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4516 31578 4522 31580
rect 4276 31526 4278 31578
rect 4458 31526 4460 31578
rect 4214 31524 4220 31526
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4516 31524 4522 31526
rect 4214 31504 4522 31524
rect 4158 31376 4214 31385
rect 4158 31311 4214 31320
rect 3988 30790 4108 30818
rect 3884 29232 3936 29238
rect 3884 29174 3936 29180
rect 3884 29028 3936 29034
rect 3884 28970 3936 28976
rect 3792 25492 3844 25498
rect 3792 25434 3844 25440
rect 3896 25378 3924 28970
rect 3804 25350 3924 25378
rect 3804 24698 3832 25350
rect 3884 25220 3936 25226
rect 3884 25162 3936 25168
rect 3896 24857 3924 25162
rect 3882 24848 3938 24857
rect 3882 24783 3938 24792
rect 3804 24670 3924 24698
rect 3792 24608 3844 24614
rect 3792 24550 3844 24556
rect 3804 24274 3832 24550
rect 3792 24268 3844 24274
rect 3792 24210 3844 24216
rect 3792 24064 3844 24070
rect 3792 24006 3844 24012
rect 3804 23730 3832 24006
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3792 23588 3844 23594
rect 3792 23530 3844 23536
rect 3804 18578 3832 23530
rect 3896 23202 3924 24670
rect 3988 23866 4016 30790
rect 4172 30682 4200 31311
rect 4080 30654 4200 30682
rect 4080 30274 4108 30654
rect 4214 30492 4522 30512
rect 4214 30490 4220 30492
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4516 30490 4522 30492
rect 4276 30438 4278 30490
rect 4458 30438 4460 30490
rect 4214 30436 4220 30438
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4516 30436 4522 30438
rect 4214 30416 4522 30436
rect 4080 30246 4200 30274
rect 4172 29594 4200 30246
rect 4080 29566 4200 29594
rect 4080 29186 4108 29566
rect 4214 29404 4522 29424
rect 4214 29402 4220 29404
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4516 29402 4522 29404
rect 4276 29350 4278 29402
rect 4458 29350 4460 29402
rect 4214 29348 4220 29350
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4516 29348 4522 29350
rect 4214 29328 4522 29348
rect 4080 29158 4200 29186
rect 4068 29096 4120 29102
rect 4066 29064 4068 29073
rect 4120 29064 4122 29073
rect 4066 28999 4122 29008
rect 4172 28506 4200 29158
rect 4080 28478 4200 28506
rect 4080 28098 4108 28478
rect 4214 28316 4522 28336
rect 4214 28314 4220 28316
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4516 28314 4522 28316
rect 4276 28262 4278 28314
rect 4458 28262 4460 28314
rect 4214 28260 4220 28262
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4516 28260 4522 28262
rect 4214 28240 4522 28260
rect 4080 28070 4200 28098
rect 4172 27316 4200 28070
rect 4080 27288 4200 27316
rect 4080 27112 4108 27288
rect 4214 27228 4522 27248
rect 4214 27226 4220 27228
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4516 27226 4522 27228
rect 4276 27174 4278 27226
rect 4458 27174 4460 27226
rect 4214 27172 4220 27174
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4516 27172 4522 27174
rect 4214 27152 4522 27172
rect 4080 27084 4200 27112
rect 4172 26296 4200 27084
rect 4528 27056 4580 27062
rect 4526 27024 4528 27033
rect 4580 27024 4582 27033
rect 4526 26959 4582 26968
rect 4080 26268 4200 26296
rect 4080 25922 4108 26268
rect 4214 26140 4522 26160
rect 4214 26138 4220 26140
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4516 26138 4522 26140
rect 4276 26086 4278 26138
rect 4458 26086 4460 26138
rect 4214 26084 4220 26086
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4516 26084 4522 26086
rect 4214 26064 4522 26084
rect 4080 25894 4200 25922
rect 4172 25242 4200 25894
rect 4080 25214 4200 25242
rect 4080 24834 4108 25214
rect 4214 25052 4522 25072
rect 4214 25050 4220 25052
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4516 25050 4522 25052
rect 4276 24998 4278 25050
rect 4458 24998 4460 25050
rect 4214 24996 4220 24998
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4516 24996 4522 24998
rect 4214 24976 4522 24996
rect 4080 24806 4200 24834
rect 4172 24154 4200 24806
rect 4080 24126 4200 24154
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 4080 23746 4108 24126
rect 4214 23964 4522 23984
rect 4214 23962 4220 23964
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4516 23962 4522 23964
rect 4276 23910 4278 23962
rect 4458 23910 4460 23962
rect 4214 23908 4220 23910
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4516 23908 4522 23910
rect 4214 23888 4522 23908
rect 4528 23792 4580 23798
rect 4080 23718 4200 23746
rect 4528 23734 4580 23740
rect 4068 23520 4120 23526
rect 4068 23462 4120 23468
rect 3896 23174 4016 23202
rect 3884 23112 3936 23118
rect 3884 23054 3936 23060
rect 3896 22681 3924 23054
rect 3882 22672 3938 22681
rect 3882 22607 3938 22616
rect 3988 22556 4016 23174
rect 3896 22528 4016 22556
rect 3896 18698 3924 22528
rect 3976 22432 4028 22438
rect 3976 22374 4028 22380
rect 3988 21486 4016 22374
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3884 18692 3936 18698
rect 3884 18634 3936 18640
rect 3804 18550 3924 18578
rect 3712 18414 3832 18442
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3712 18193 3740 18226
rect 3698 18184 3754 18193
rect 3698 18119 3754 18128
rect 3608 17876 3660 17882
rect 3608 17818 3660 17824
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3422 15736 3478 15745
rect 3422 15671 3478 15680
rect 3528 15620 3556 17546
rect 3436 15592 3556 15620
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3436 14260 3464 15592
rect 3516 15428 3568 15434
rect 3516 15370 3568 15376
rect 3344 14232 3464 14260
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3252 12850 3280 13126
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3344 12730 3372 14232
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3436 13297 3464 13874
rect 3422 13288 3478 13297
rect 3422 13223 3478 13232
rect 3528 13172 3556 15370
rect 3620 14113 3648 17818
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3606 14104 3662 14113
rect 3606 14039 3662 14048
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3252 12702 3372 12730
rect 3436 13144 3556 13172
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 3252 11830 3280 12702
rect 3436 12594 3464 13144
rect 3514 13016 3570 13025
rect 3514 12951 3570 12960
rect 3344 12566 3464 12594
rect 3240 11824 3292 11830
rect 3054 11792 3110 11801
rect 3240 11766 3292 11772
rect 3054 11727 3056 11736
rect 3108 11727 3110 11736
rect 3056 11698 3108 11704
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2962 11520 3018 11529
rect 2582 11452 2890 11472
rect 2962 11455 3018 11464
rect 2582 11450 2588 11452
rect 2644 11450 2668 11452
rect 2724 11450 2748 11452
rect 2804 11450 2828 11452
rect 2884 11450 2890 11452
rect 2644 11398 2646 11450
rect 2826 11398 2828 11450
rect 2582 11396 2588 11398
rect 2644 11396 2668 11398
rect 2724 11396 2748 11398
rect 2804 11396 2828 11398
rect 2884 11396 2890 11398
rect 2582 11376 2890 11396
rect 2582 10364 2890 10384
rect 2582 10362 2588 10364
rect 2644 10362 2668 10364
rect 2724 10362 2748 10364
rect 2804 10362 2828 10364
rect 2884 10362 2890 10364
rect 2644 10310 2646 10362
rect 2826 10310 2828 10362
rect 2582 10308 2588 10310
rect 2644 10308 2668 10310
rect 2724 10308 2748 10310
rect 2804 10308 2828 10310
rect 2884 10308 2890 10310
rect 2582 10288 2890 10308
rect 2582 9276 2890 9296
rect 2582 9274 2588 9276
rect 2644 9274 2668 9276
rect 2724 9274 2748 9276
rect 2804 9274 2828 9276
rect 2884 9274 2890 9276
rect 2644 9222 2646 9274
rect 2826 9222 2828 9274
rect 2582 9220 2588 9222
rect 2644 9220 2668 9222
rect 2724 9220 2748 9222
rect 2804 9220 2828 9222
rect 2884 9220 2890 9222
rect 2582 9200 2890 9220
rect 2976 8650 3004 11455
rect 3068 11218 3096 11698
rect 3344 11354 3372 12566
rect 3422 12472 3478 12481
rect 3422 12407 3478 12416
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3436 11286 3464 12407
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 3068 9178 3096 9386
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2884 8622 3004 8650
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2884 8362 2912 8622
rect 3068 8498 3096 8774
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2582 8188 2890 8208
rect 2582 8186 2588 8188
rect 2644 8186 2668 8188
rect 2724 8186 2748 8188
rect 2804 8186 2828 8188
rect 2884 8186 2890 8188
rect 2644 8134 2646 8186
rect 2826 8134 2828 8186
rect 2582 8132 2588 8134
rect 2644 8132 2668 8134
rect 2724 8132 2748 8134
rect 2804 8132 2828 8134
rect 2884 8132 2890 8134
rect 2582 8112 2890 8132
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2700 7478 2728 7822
rect 2688 7472 2740 7478
rect 2976 7449 3004 8434
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 2688 7414 2740 7420
rect 2962 7440 3018 7449
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2136 7404 2188 7410
rect 2962 7375 3018 7384
rect 2136 7346 2188 7352
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1964 6202 1992 6734
rect 1872 6174 1992 6202
rect 1872 4622 1900 6174
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1964 4826 1992 5170
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1596 3590 1716 3618
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1596 3097 1624 3470
rect 1688 3194 1716 3590
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1582 3088 1638 3097
rect 1582 3023 1638 3032
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 1780 2310 1808 4014
rect 2056 3942 2084 7346
rect 2148 6798 2176 7346
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2424 6322 2452 7142
rect 2582 7100 2890 7120
rect 2582 7098 2588 7100
rect 2644 7098 2668 7100
rect 2724 7098 2748 7100
rect 2804 7098 2828 7100
rect 2884 7098 2890 7100
rect 2644 7046 2646 7098
rect 2826 7046 2828 7098
rect 2582 7044 2588 7046
rect 2644 7044 2668 7046
rect 2724 7044 2748 7046
rect 2804 7044 2828 7046
rect 2884 7044 2890 7046
rect 2582 7024 2890 7044
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2594 6760 2650 6769
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2056 3194 2084 3878
rect 2240 3738 2268 5646
rect 2516 4622 2544 6734
rect 2594 6695 2650 6704
rect 2608 6458 2636 6695
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2976 6225 3004 7278
rect 3068 6390 3096 8298
rect 3160 6866 3188 9998
rect 3252 8974 3280 10610
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 3160 6497 3188 6666
rect 3146 6488 3202 6497
rect 3146 6423 3202 6432
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 2962 6216 3018 6225
rect 2962 6151 3018 6160
rect 2582 6012 2890 6032
rect 2582 6010 2588 6012
rect 2644 6010 2668 6012
rect 2724 6010 2748 6012
rect 2804 6010 2828 6012
rect 2884 6010 2890 6012
rect 2644 5958 2646 6010
rect 2826 5958 2828 6010
rect 2582 5956 2588 5958
rect 2644 5956 2668 5958
rect 2724 5956 2748 5958
rect 2804 5956 2828 5958
rect 2884 5956 2890 5958
rect 2582 5936 2890 5956
rect 2962 5944 3018 5953
rect 2962 5879 2964 5888
rect 3016 5879 3018 5888
rect 2964 5850 3016 5856
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2884 5273 2912 5306
rect 2870 5264 2926 5273
rect 2870 5199 2926 5208
rect 2582 4924 2890 4944
rect 2582 4922 2588 4924
rect 2644 4922 2668 4924
rect 2724 4922 2748 4924
rect 2804 4922 2828 4924
rect 2884 4922 2890 4924
rect 2644 4870 2646 4922
rect 2826 4870 2828 4922
rect 2582 4868 2588 4870
rect 2644 4868 2668 4870
rect 2724 4868 2748 4870
rect 2804 4868 2828 4870
rect 2884 4868 2890 4870
rect 2582 4848 2890 4868
rect 3068 4622 3096 6326
rect 3252 5370 3280 8910
rect 3344 6322 3372 11018
rect 3528 10826 3556 12951
rect 3436 10798 3556 10826
rect 3436 9586 3464 10798
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 2240 1873 2268 2994
rect 2332 2582 2360 4490
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2424 3534 2452 4082
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2424 2650 2452 3470
rect 2516 3194 2544 4558
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 2700 4078 2728 4490
rect 2792 4146 2820 4558
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2582 3836 2890 3856
rect 2582 3834 2588 3836
rect 2644 3834 2668 3836
rect 2724 3834 2748 3836
rect 2804 3834 2828 3836
rect 2884 3834 2890 3836
rect 2644 3782 2646 3834
rect 2826 3782 2828 3834
rect 2582 3780 2588 3782
rect 2644 3780 2668 3782
rect 2724 3780 2748 3782
rect 2804 3780 2828 3782
rect 2884 3780 2890 3782
rect 2582 3760 2890 3780
rect 3344 3194 3372 6258
rect 3436 5778 3464 9522
rect 3528 7546 3556 10610
rect 3620 8634 3648 13942
rect 3712 12714 3740 16050
rect 3804 12850 3832 18414
rect 3896 17814 3924 18550
rect 3988 18465 4016 18702
rect 3974 18456 4030 18465
rect 3974 18391 4030 18400
rect 3884 17808 3936 17814
rect 3884 17750 3936 17756
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 3896 13433 3924 17206
rect 3988 17202 4016 17478
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3988 16289 4016 16526
rect 3974 16280 4030 16289
rect 3974 16215 4030 16224
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 14249 4016 14350
rect 3974 14240 4030 14249
rect 3974 14175 4030 14184
rect 3882 13424 3938 13433
rect 3882 13359 3938 13368
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3884 13252 3936 13258
rect 3884 13194 3936 13200
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3712 11665 3740 11698
rect 3698 11656 3754 11665
rect 3698 11591 3754 11600
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3620 7313 3648 7346
rect 3606 7304 3662 7313
rect 3606 7239 3662 7248
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3620 4457 3648 5170
rect 3712 4690 3740 11494
rect 3804 7546 3832 12786
rect 3896 12306 3924 13194
rect 3988 12889 4016 13262
rect 3974 12880 4030 12889
rect 3974 12815 4030 12824
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3896 11762 3924 12242
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3988 10418 4016 12650
rect 4080 10674 4108 23462
rect 4172 23322 4200 23718
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 4540 23050 4568 23734
rect 4528 23044 4580 23050
rect 4528 22986 4580 22992
rect 4214 22876 4522 22896
rect 4214 22874 4220 22876
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4516 22874 4522 22876
rect 4276 22822 4278 22874
rect 4458 22822 4460 22874
rect 4214 22820 4220 22822
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4516 22820 4522 22822
rect 4214 22800 4522 22820
rect 4214 21788 4522 21808
rect 4214 21786 4220 21788
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4516 21786 4522 21788
rect 4276 21734 4278 21786
rect 4458 21734 4460 21786
rect 4214 21732 4220 21734
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4516 21732 4522 21734
rect 4214 21712 4522 21732
rect 4214 20700 4522 20720
rect 4214 20698 4220 20700
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4516 20698 4522 20700
rect 4276 20646 4278 20698
rect 4458 20646 4460 20698
rect 4214 20644 4220 20646
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4516 20644 4522 20646
rect 4214 20624 4522 20644
rect 4214 19612 4522 19632
rect 4214 19610 4220 19612
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4516 19610 4522 19612
rect 4276 19558 4278 19610
rect 4458 19558 4460 19610
rect 4214 19556 4220 19558
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4516 19556 4522 19558
rect 4214 19536 4522 19556
rect 4214 18524 4522 18544
rect 4214 18522 4220 18524
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4516 18522 4522 18524
rect 4276 18470 4278 18522
rect 4458 18470 4460 18522
rect 4214 18468 4220 18470
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4516 18468 4522 18470
rect 4214 18448 4522 18468
rect 4214 17436 4522 17456
rect 4214 17434 4220 17436
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4516 17434 4522 17436
rect 4276 17382 4278 17434
rect 4458 17382 4460 17434
rect 4214 17380 4220 17382
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4516 17380 4522 17382
rect 4214 17360 4522 17380
rect 4632 17218 4660 31640
rect 4712 31622 4764 31628
rect 4724 23066 4752 31622
rect 4816 23610 4844 31758
rect 4908 23730 4936 31844
rect 4986 31784 5042 31793
rect 4986 31719 5042 31728
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 4816 23582 4936 23610
rect 4724 23038 4844 23066
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4724 17338 4752 22918
rect 4816 21690 4844 23038
rect 4908 22953 4936 23582
rect 5000 23322 5028 31719
rect 5092 31482 5120 36366
rect 5080 31476 5132 31482
rect 5080 31418 5132 31424
rect 5080 31340 5132 31346
rect 5080 31282 5132 31288
rect 5092 23866 5120 31282
rect 5080 23860 5132 23866
rect 5080 23802 5132 23808
rect 5080 23724 5132 23730
rect 5080 23666 5132 23672
rect 4988 23316 5040 23322
rect 4988 23258 5040 23264
rect 4894 22944 4950 22953
rect 4894 22879 4950 22888
rect 4894 22672 4950 22681
rect 4894 22607 4950 22616
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4632 17190 4752 17218
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4214 16348 4522 16368
rect 4214 16346 4220 16348
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4516 16346 4522 16348
rect 4276 16294 4278 16346
rect 4458 16294 4460 16346
rect 4214 16292 4220 16294
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4516 16292 4522 16294
rect 4214 16272 4522 16292
rect 4214 15260 4522 15280
rect 4214 15258 4220 15260
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4516 15258 4522 15260
rect 4276 15206 4278 15258
rect 4458 15206 4460 15258
rect 4214 15204 4220 15206
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4516 15204 4522 15206
rect 4214 15184 4522 15204
rect 4214 14172 4522 14192
rect 4214 14170 4220 14172
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4516 14170 4522 14172
rect 4276 14118 4278 14170
rect 4458 14118 4460 14170
rect 4214 14116 4220 14118
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4516 14116 4522 14118
rect 4214 14096 4522 14116
rect 4214 13084 4522 13104
rect 4214 13082 4220 13084
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4516 13082 4522 13084
rect 4276 13030 4278 13082
rect 4458 13030 4460 13082
rect 4214 13028 4220 13030
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4516 13028 4522 13030
rect 4214 13008 4522 13028
rect 4632 12322 4660 16934
rect 4724 12442 4752 17190
rect 4816 16998 4844 21490
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4632 12294 4844 12322
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4214 11996 4522 12016
rect 4214 11994 4220 11996
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4516 11994 4522 11996
rect 4276 11942 4278 11994
rect 4458 11942 4460 11994
rect 4214 11940 4220 11942
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4516 11940 4522 11942
rect 4214 11920 4522 11940
rect 4214 10908 4522 10928
rect 4214 10906 4220 10908
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4516 10906 4522 10908
rect 4276 10854 4278 10906
rect 4458 10854 4460 10906
rect 4214 10852 4220 10854
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4516 10852 4522 10854
rect 4214 10832 4522 10852
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 3896 10390 4016 10418
rect 3896 9654 3924 10390
rect 3974 10296 4030 10305
rect 3974 10231 3976 10240
rect 4028 10231 4030 10240
rect 3976 10202 4028 10208
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3896 7886 3924 9114
rect 3988 8974 4016 9998
rect 4214 9820 4522 9840
rect 4214 9818 4220 9820
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4516 9818 4522 9820
rect 4276 9766 4278 9818
rect 4458 9766 4460 9818
rect 4214 9764 4220 9766
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4516 9764 4522 9766
rect 4214 9744 4522 9764
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3896 5794 3924 7822
rect 3988 5914 4016 8910
rect 4214 8732 4522 8752
rect 4214 8730 4220 8732
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4516 8730 4522 8732
rect 4276 8678 4278 8730
rect 4458 8678 4460 8730
rect 4214 8676 4220 8678
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4516 8676 4522 8678
rect 4214 8656 4522 8676
rect 4214 7644 4522 7664
rect 4214 7642 4220 7644
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4516 7642 4522 7644
rect 4276 7590 4278 7642
rect 4458 7590 4460 7642
rect 4214 7588 4220 7590
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4516 7588 4522 7590
rect 4214 7568 4522 7588
rect 4632 6866 4660 12174
rect 4724 10198 4752 12174
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4816 10010 4844 12294
rect 4908 10538 4936 22607
rect 5092 22098 5120 23666
rect 5080 22092 5132 22098
rect 5080 22034 5132 22040
rect 5184 19242 5212 50895
rect 5460 50844 5488 51031
rect 5552 50969 5580 51462
rect 5644 51105 5672 52430
rect 5630 51096 5686 51105
rect 5630 51031 5686 51040
rect 5538 50960 5594 50969
rect 5538 50895 5594 50904
rect 5632 50856 5684 50862
rect 5354 50824 5410 50833
rect 5460 50816 5580 50844
rect 5354 50759 5410 50768
rect 5262 50688 5318 50697
rect 5262 50623 5318 50632
rect 5276 49298 5304 50623
rect 5264 49292 5316 49298
rect 5264 49234 5316 49240
rect 5264 48136 5316 48142
rect 5264 48078 5316 48084
rect 5276 41682 5304 48078
rect 5368 45665 5396 50759
rect 5552 50674 5580 50816
rect 5632 50798 5684 50804
rect 5460 50646 5580 50674
rect 5354 45656 5410 45665
rect 5354 45591 5410 45600
rect 5356 45484 5408 45490
rect 5356 45426 5408 45432
rect 5368 45082 5396 45426
rect 5356 45076 5408 45082
rect 5356 45018 5408 45024
rect 5354 44976 5410 44985
rect 5354 44911 5410 44920
rect 5264 41676 5316 41682
rect 5264 41618 5316 41624
rect 5368 41562 5396 44911
rect 5460 41614 5488 50646
rect 5540 50312 5592 50318
rect 5540 50254 5592 50260
rect 5552 48618 5580 50254
rect 5540 48612 5592 48618
rect 5540 48554 5592 48560
rect 5644 48314 5672 50798
rect 5552 48286 5672 48314
rect 5552 45558 5580 48286
rect 5540 45552 5592 45558
rect 5540 45494 5592 45500
rect 5540 44872 5592 44878
rect 5540 44814 5592 44820
rect 5552 43722 5580 44814
rect 5632 44736 5684 44742
rect 5632 44678 5684 44684
rect 5644 43926 5672 44678
rect 5632 43920 5684 43926
rect 5632 43862 5684 43868
rect 5540 43716 5592 43722
rect 5540 43658 5592 43664
rect 5644 41993 5672 43862
rect 5630 41984 5686 41993
rect 5630 41919 5686 41928
rect 5276 41534 5396 41562
rect 5448 41608 5500 41614
rect 5448 41550 5500 41556
rect 5276 31657 5304 41534
rect 5354 41440 5410 41449
rect 5736 41414 5764 55655
rect 5846 54972 6154 54992
rect 5846 54970 5852 54972
rect 5908 54970 5932 54972
rect 5988 54970 6012 54972
rect 6068 54970 6092 54972
rect 6148 54970 6154 54972
rect 5908 54918 5910 54970
rect 6090 54918 6092 54970
rect 5846 54916 5852 54918
rect 5908 54916 5932 54918
rect 5988 54916 6012 54918
rect 6068 54916 6092 54918
rect 6148 54916 6154 54918
rect 5846 54896 6154 54916
rect 5846 53884 6154 53904
rect 5846 53882 5852 53884
rect 5908 53882 5932 53884
rect 5988 53882 6012 53884
rect 6068 53882 6092 53884
rect 6148 53882 6154 53884
rect 5908 53830 5910 53882
rect 6090 53830 6092 53882
rect 5846 53828 5852 53830
rect 5908 53828 5932 53830
rect 5988 53828 6012 53830
rect 6068 53828 6092 53830
rect 6148 53828 6154 53830
rect 5846 53808 6154 53828
rect 6184 53168 6236 53174
rect 6184 53110 6236 53116
rect 5846 52796 6154 52816
rect 5846 52794 5852 52796
rect 5908 52794 5932 52796
rect 5988 52794 6012 52796
rect 6068 52794 6092 52796
rect 6148 52794 6154 52796
rect 5908 52742 5910 52794
rect 6090 52742 6092 52794
rect 5846 52740 5852 52742
rect 5908 52740 5932 52742
rect 5988 52740 6012 52742
rect 6068 52740 6092 52742
rect 6148 52740 6154 52742
rect 5846 52720 6154 52740
rect 5846 51708 6154 51728
rect 5846 51706 5852 51708
rect 5908 51706 5932 51708
rect 5988 51706 6012 51708
rect 6068 51706 6092 51708
rect 6148 51706 6154 51708
rect 5908 51654 5910 51706
rect 6090 51654 6092 51706
rect 5846 51652 5852 51654
rect 5908 51652 5932 51654
rect 5988 51652 6012 51654
rect 6068 51652 6092 51654
rect 6148 51652 6154 51654
rect 5846 51632 6154 51652
rect 5846 50620 6154 50640
rect 5846 50618 5852 50620
rect 5908 50618 5932 50620
rect 5988 50618 6012 50620
rect 6068 50618 6092 50620
rect 6148 50618 6154 50620
rect 5908 50566 5910 50618
rect 6090 50566 6092 50618
rect 5846 50564 5852 50566
rect 5908 50564 5932 50566
rect 5988 50564 6012 50566
rect 6068 50564 6092 50566
rect 6148 50564 6154 50566
rect 5846 50544 6154 50564
rect 5846 49532 6154 49552
rect 5846 49530 5852 49532
rect 5908 49530 5932 49532
rect 5988 49530 6012 49532
rect 6068 49530 6092 49532
rect 6148 49530 6154 49532
rect 5908 49478 5910 49530
rect 6090 49478 6092 49530
rect 5846 49476 5852 49478
rect 5908 49476 5932 49478
rect 5988 49476 6012 49478
rect 6068 49476 6092 49478
rect 6148 49476 6154 49478
rect 5846 49456 6154 49476
rect 5846 48444 6154 48464
rect 5846 48442 5852 48444
rect 5908 48442 5932 48444
rect 5988 48442 6012 48444
rect 6068 48442 6092 48444
rect 6148 48442 6154 48444
rect 5908 48390 5910 48442
rect 6090 48390 6092 48442
rect 5846 48388 5852 48390
rect 5908 48388 5932 48390
rect 5988 48388 6012 48390
rect 6068 48388 6092 48390
rect 6148 48388 6154 48390
rect 5846 48368 6154 48388
rect 5846 47356 6154 47376
rect 5846 47354 5852 47356
rect 5908 47354 5932 47356
rect 5988 47354 6012 47356
rect 6068 47354 6092 47356
rect 6148 47354 6154 47356
rect 5908 47302 5910 47354
rect 6090 47302 6092 47354
rect 5846 47300 5852 47302
rect 5908 47300 5932 47302
rect 5988 47300 6012 47302
rect 6068 47300 6092 47302
rect 6148 47300 6154 47302
rect 5846 47280 6154 47300
rect 5846 46268 6154 46288
rect 5846 46266 5852 46268
rect 5908 46266 5932 46268
rect 5988 46266 6012 46268
rect 6068 46266 6092 46268
rect 6148 46266 6154 46268
rect 5908 46214 5910 46266
rect 6090 46214 6092 46266
rect 5846 46212 5852 46214
rect 5908 46212 5932 46214
rect 5988 46212 6012 46214
rect 6068 46212 6092 46214
rect 6148 46212 6154 46214
rect 5846 46192 6154 46212
rect 5846 45180 6154 45200
rect 5846 45178 5852 45180
rect 5908 45178 5932 45180
rect 5988 45178 6012 45180
rect 6068 45178 6092 45180
rect 6148 45178 6154 45180
rect 5908 45126 5910 45178
rect 6090 45126 6092 45178
rect 5846 45124 5852 45126
rect 5908 45124 5932 45126
rect 5988 45124 6012 45126
rect 6068 45124 6092 45126
rect 6148 45124 6154 45126
rect 5846 45104 6154 45124
rect 6196 44826 6224 53110
rect 6288 49638 6316 57258
rect 6460 56908 6512 56914
rect 6460 56850 6512 56856
rect 6368 55684 6420 55690
rect 6368 55626 6420 55632
rect 6276 49632 6328 49638
rect 6276 49574 6328 49580
rect 6196 44798 6316 44826
rect 6184 44736 6236 44742
rect 6184 44678 6236 44684
rect 5846 44092 6154 44112
rect 5846 44090 5852 44092
rect 5908 44090 5932 44092
rect 5988 44090 6012 44092
rect 6068 44090 6092 44092
rect 6148 44090 6154 44092
rect 5908 44038 5910 44090
rect 6090 44038 6092 44090
rect 5846 44036 5852 44038
rect 5908 44036 5932 44038
rect 5988 44036 6012 44038
rect 6068 44036 6092 44038
rect 6148 44036 6154 44038
rect 5846 44016 6154 44036
rect 5846 43004 6154 43024
rect 5846 43002 5852 43004
rect 5908 43002 5932 43004
rect 5988 43002 6012 43004
rect 6068 43002 6092 43004
rect 6148 43002 6154 43004
rect 5908 42950 5910 43002
rect 6090 42950 6092 43002
rect 5846 42948 5852 42950
rect 5908 42948 5932 42950
rect 5988 42948 6012 42950
rect 6068 42948 6092 42950
rect 6148 42948 6154 42950
rect 5846 42928 6154 42948
rect 5846 41916 6154 41936
rect 5846 41914 5852 41916
rect 5908 41914 5932 41916
rect 5988 41914 6012 41916
rect 6068 41914 6092 41916
rect 6148 41914 6154 41916
rect 5908 41862 5910 41914
rect 6090 41862 6092 41914
rect 5846 41860 5852 41862
rect 5908 41860 5932 41862
rect 5988 41860 6012 41862
rect 6068 41860 6092 41862
rect 6148 41860 6154 41862
rect 5846 41840 6154 41860
rect 5908 41608 5960 41614
rect 5908 41550 5960 41556
rect 5816 41540 5868 41546
rect 5816 41482 5868 41488
rect 5354 41375 5410 41384
rect 5644 41386 5764 41414
rect 5368 40662 5396 41375
rect 5644 41256 5672 41386
rect 5644 41228 5764 41256
rect 5540 41200 5592 41206
rect 5540 41142 5592 41148
rect 5448 40928 5500 40934
rect 5448 40870 5500 40876
rect 5356 40656 5408 40662
rect 5356 40598 5408 40604
rect 5356 40520 5408 40526
rect 5356 40462 5408 40468
rect 5368 38554 5396 40462
rect 5460 40118 5488 40870
rect 5448 40112 5500 40118
rect 5448 40054 5500 40060
rect 5448 39976 5500 39982
rect 5448 39918 5500 39924
rect 5356 38548 5408 38554
rect 5356 38490 5408 38496
rect 5356 38344 5408 38350
rect 5356 38286 5408 38292
rect 5368 37874 5396 38286
rect 5356 37868 5408 37874
rect 5356 37810 5408 37816
rect 5368 36961 5396 37810
rect 5354 36952 5410 36961
rect 5354 36887 5410 36896
rect 5460 36768 5488 39918
rect 5368 36740 5488 36768
rect 5368 36689 5396 36740
rect 5354 36680 5410 36689
rect 5354 36615 5410 36624
rect 5448 36644 5500 36650
rect 5448 36586 5500 36592
rect 5356 36576 5408 36582
rect 5356 36518 5408 36524
rect 5262 31648 5318 31657
rect 5262 31583 5318 31592
rect 5264 31476 5316 31482
rect 5264 31418 5316 31424
rect 5276 23866 5304 31418
rect 5264 23860 5316 23866
rect 5264 23802 5316 23808
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5276 22710 5304 23666
rect 5264 22704 5316 22710
rect 5264 22646 5316 22652
rect 5172 19236 5224 19242
rect 5172 19178 5224 19184
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 5000 15638 5028 17274
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4724 9982 4844 10010
rect 4724 9586 4752 9982
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4214 6556 4522 6576
rect 4214 6554 4220 6556
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4516 6554 4522 6556
rect 4276 6502 4278 6554
rect 4458 6502 4460 6554
rect 4214 6500 4220 6502
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4516 6500 4522 6502
rect 4214 6480 4522 6500
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3896 5766 4016 5794
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3606 4448 3662 4457
rect 3606 4383 3662 4392
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 2582 2748 2890 2768
rect 2582 2746 2588 2748
rect 2644 2746 2668 2748
rect 2724 2746 2748 2748
rect 2804 2746 2828 2748
rect 2884 2746 2890 2748
rect 2644 2694 2646 2746
rect 2826 2694 2828 2746
rect 2582 2692 2588 2694
rect 2644 2692 2668 2694
rect 2724 2692 2748 2694
rect 2804 2692 2828 2694
rect 2884 2692 2890 2694
rect 2582 2672 2890 2692
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 2320 2576 2372 2582
rect 2320 2518 2372 2524
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2226 1864 2282 1873
rect 2226 1799 2282 1808
rect 2792 649 2820 2314
rect 2884 1465 2912 2382
rect 2976 2281 3004 2994
rect 3528 2553 3556 2994
rect 3896 2650 3924 4626
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3988 2582 4016 5766
rect 4160 5704 4212 5710
rect 4080 5652 4160 5658
rect 4080 5646 4212 5652
rect 4080 5630 4200 5646
rect 4080 4729 4108 5630
rect 4214 5468 4522 5488
rect 4214 5466 4220 5468
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4516 5466 4522 5468
rect 4276 5414 4278 5466
rect 4458 5414 4460 5466
rect 4214 5412 4220 5414
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4516 5412 4522 5414
rect 4214 5392 4522 5412
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4540 4826 4568 5170
rect 4724 5166 4752 9522
rect 5368 8090 5396 36518
rect 5460 21622 5488 36586
rect 5552 36582 5580 41142
rect 5632 41132 5684 41138
rect 5632 41074 5684 41080
rect 5644 39982 5672 41074
rect 5632 39976 5684 39982
rect 5632 39918 5684 39924
rect 5632 39432 5684 39438
rect 5632 39374 5684 39380
rect 5644 39030 5672 39374
rect 5632 39024 5684 39030
rect 5632 38966 5684 38972
rect 5736 38400 5764 41228
rect 5828 41070 5856 41482
rect 5920 41138 5948 41550
rect 5908 41132 5960 41138
rect 5908 41074 5960 41080
rect 5816 41064 5868 41070
rect 5816 41006 5868 41012
rect 5846 40828 6154 40848
rect 5846 40826 5852 40828
rect 5908 40826 5932 40828
rect 5988 40826 6012 40828
rect 6068 40826 6092 40828
rect 6148 40826 6154 40828
rect 5908 40774 5910 40826
rect 6090 40774 6092 40826
rect 5846 40772 5852 40774
rect 5908 40772 5932 40774
rect 5988 40772 6012 40774
rect 6068 40772 6092 40774
rect 6148 40772 6154 40774
rect 5846 40752 6154 40772
rect 5846 39740 6154 39760
rect 5846 39738 5852 39740
rect 5908 39738 5932 39740
rect 5988 39738 6012 39740
rect 6068 39738 6092 39740
rect 6148 39738 6154 39740
rect 5908 39686 5910 39738
rect 6090 39686 6092 39738
rect 5846 39684 5852 39686
rect 5908 39684 5932 39686
rect 5988 39684 6012 39686
rect 6068 39684 6092 39686
rect 6148 39684 6154 39686
rect 5846 39664 6154 39684
rect 5846 38652 6154 38672
rect 5846 38650 5852 38652
rect 5908 38650 5932 38652
rect 5988 38650 6012 38652
rect 6068 38650 6092 38652
rect 6148 38650 6154 38652
rect 5908 38598 5910 38650
rect 6090 38598 6092 38650
rect 5846 38596 5852 38598
rect 5908 38596 5932 38598
rect 5988 38596 6012 38598
rect 6068 38596 6092 38598
rect 6148 38596 6154 38598
rect 5846 38576 6154 38596
rect 5644 38372 5764 38400
rect 5540 36576 5592 36582
rect 5540 36518 5592 36524
rect 5538 36408 5594 36417
rect 5538 36343 5594 36352
rect 5552 35698 5580 36343
rect 5540 35692 5592 35698
rect 5540 35634 5592 35640
rect 5540 34604 5592 34610
rect 5540 34546 5592 34552
rect 5552 33658 5580 34546
rect 5644 34134 5672 38372
rect 5724 38276 5776 38282
rect 5724 38218 5776 38224
rect 5736 37330 5764 38218
rect 5846 37564 6154 37584
rect 5846 37562 5852 37564
rect 5908 37562 5932 37564
rect 5988 37562 6012 37564
rect 6068 37562 6092 37564
rect 6148 37562 6154 37564
rect 5908 37510 5910 37562
rect 6090 37510 6092 37562
rect 5846 37508 5852 37510
rect 5908 37508 5932 37510
rect 5988 37508 6012 37510
rect 6068 37508 6092 37510
rect 6148 37508 6154 37510
rect 5846 37488 6154 37508
rect 5724 37324 5776 37330
rect 5724 37266 5776 37272
rect 5632 34128 5684 34134
rect 5632 34070 5684 34076
rect 5632 33992 5684 33998
rect 5632 33934 5684 33940
rect 5540 33652 5592 33658
rect 5540 33594 5592 33600
rect 5644 33522 5672 33934
rect 5632 33516 5684 33522
rect 5632 33458 5684 33464
rect 5632 33380 5684 33386
rect 5632 33322 5684 33328
rect 5644 32298 5672 33322
rect 5632 32292 5684 32298
rect 5632 32234 5684 32240
rect 5736 23254 5764 37266
rect 5846 36476 6154 36496
rect 5846 36474 5852 36476
rect 5908 36474 5932 36476
rect 5988 36474 6012 36476
rect 6068 36474 6092 36476
rect 6148 36474 6154 36476
rect 5908 36422 5910 36474
rect 6090 36422 6092 36474
rect 5846 36420 5852 36422
rect 5908 36420 5932 36422
rect 5988 36420 6012 36422
rect 6068 36420 6092 36422
rect 6148 36420 6154 36422
rect 5846 36400 6154 36420
rect 5846 35388 6154 35408
rect 5846 35386 5852 35388
rect 5908 35386 5932 35388
rect 5988 35386 6012 35388
rect 6068 35386 6092 35388
rect 6148 35386 6154 35388
rect 5908 35334 5910 35386
rect 6090 35334 6092 35386
rect 5846 35332 5852 35334
rect 5908 35332 5932 35334
rect 5988 35332 6012 35334
rect 6068 35332 6092 35334
rect 6148 35332 6154 35334
rect 5846 35312 6154 35332
rect 5846 34300 6154 34320
rect 5846 34298 5852 34300
rect 5908 34298 5932 34300
rect 5988 34298 6012 34300
rect 6068 34298 6092 34300
rect 6148 34298 6154 34300
rect 5908 34246 5910 34298
rect 6090 34246 6092 34298
rect 5846 34244 5852 34246
rect 5908 34244 5932 34246
rect 5988 34244 6012 34246
rect 6068 34244 6092 34246
rect 6148 34244 6154 34246
rect 5846 34224 6154 34244
rect 5816 34128 5868 34134
rect 5816 34070 5868 34076
rect 5828 33386 5856 34070
rect 5816 33380 5868 33386
rect 5816 33322 5868 33328
rect 5846 33212 6154 33232
rect 5846 33210 5852 33212
rect 5908 33210 5932 33212
rect 5988 33210 6012 33212
rect 6068 33210 6092 33212
rect 6148 33210 6154 33212
rect 5908 33158 5910 33210
rect 6090 33158 6092 33210
rect 5846 33156 5852 33158
rect 5908 33156 5932 33158
rect 5988 33156 6012 33158
rect 6068 33156 6092 33158
rect 6148 33156 6154 33158
rect 5846 33136 6154 33156
rect 5846 32124 6154 32144
rect 5846 32122 5852 32124
rect 5908 32122 5932 32124
rect 5988 32122 6012 32124
rect 6068 32122 6092 32124
rect 6148 32122 6154 32124
rect 5908 32070 5910 32122
rect 6090 32070 6092 32122
rect 5846 32068 5852 32070
rect 5908 32068 5932 32070
rect 5988 32068 6012 32070
rect 6068 32068 6092 32070
rect 6148 32068 6154 32070
rect 5846 32048 6154 32068
rect 6196 31414 6224 44678
rect 6288 43058 6316 44798
rect 6380 43450 6408 55626
rect 6472 49162 6500 56850
rect 7478 56604 7786 56624
rect 7478 56602 7484 56604
rect 7540 56602 7564 56604
rect 7620 56602 7644 56604
rect 7700 56602 7724 56604
rect 7780 56602 7786 56604
rect 7540 56550 7542 56602
rect 7722 56550 7724 56602
rect 7478 56548 7484 56550
rect 7540 56548 7564 56550
rect 7620 56548 7644 56550
rect 7700 56548 7724 56550
rect 7780 56548 7786 56550
rect 7478 56528 7786 56548
rect 7478 55516 7786 55536
rect 7478 55514 7484 55516
rect 7540 55514 7564 55516
rect 7620 55514 7644 55516
rect 7700 55514 7724 55516
rect 7780 55514 7786 55516
rect 7540 55462 7542 55514
rect 7722 55462 7724 55514
rect 7478 55460 7484 55462
rect 7540 55460 7564 55462
rect 7620 55460 7644 55462
rect 7700 55460 7724 55462
rect 7780 55460 7786 55462
rect 7478 55440 7786 55460
rect 6552 55072 6604 55078
rect 6552 55014 6604 55020
rect 6564 50454 6592 55014
rect 8312 54738 8340 59570
rect 8496 55944 8524 66982
rect 9110 66940 9418 66960
rect 9110 66938 9116 66940
rect 9172 66938 9196 66940
rect 9252 66938 9276 66940
rect 9332 66938 9356 66940
rect 9412 66938 9418 66940
rect 9172 66886 9174 66938
rect 9354 66886 9356 66938
rect 9110 66884 9116 66886
rect 9172 66884 9196 66886
rect 9252 66884 9276 66886
rect 9332 66884 9356 66886
rect 9412 66884 9418 66886
rect 9110 66864 9418 66884
rect 9692 66842 9720 67322
rect 9680 66836 9732 66842
rect 9680 66778 9732 66784
rect 9110 65852 9418 65872
rect 9110 65850 9116 65852
rect 9172 65850 9196 65852
rect 9252 65850 9276 65852
rect 9332 65850 9356 65852
rect 9412 65850 9418 65852
rect 9172 65798 9174 65850
rect 9354 65798 9356 65850
rect 9110 65796 9116 65798
rect 9172 65796 9196 65798
rect 9252 65796 9276 65798
rect 9332 65796 9356 65798
rect 9412 65796 9418 65798
rect 9110 65776 9418 65796
rect 9110 64764 9418 64784
rect 9110 64762 9116 64764
rect 9172 64762 9196 64764
rect 9252 64762 9276 64764
rect 9332 64762 9356 64764
rect 9412 64762 9418 64764
rect 9172 64710 9174 64762
rect 9354 64710 9356 64762
rect 9110 64708 9116 64710
rect 9172 64708 9196 64710
rect 9252 64708 9276 64710
rect 9332 64708 9356 64710
rect 9412 64708 9418 64710
rect 9110 64688 9418 64708
rect 9110 63676 9418 63696
rect 9110 63674 9116 63676
rect 9172 63674 9196 63676
rect 9252 63674 9276 63676
rect 9332 63674 9356 63676
rect 9412 63674 9418 63676
rect 9172 63622 9174 63674
rect 9354 63622 9356 63674
rect 9110 63620 9116 63622
rect 9172 63620 9196 63622
rect 9252 63620 9276 63622
rect 9332 63620 9356 63622
rect 9412 63620 9418 63622
rect 9110 63600 9418 63620
rect 9312 63368 9364 63374
rect 9310 63336 9312 63345
rect 9588 63368 9640 63374
rect 9364 63336 9366 63345
rect 9588 63310 9640 63316
rect 9310 63271 9366 63280
rect 9110 62588 9418 62608
rect 9110 62586 9116 62588
rect 9172 62586 9196 62588
rect 9252 62586 9276 62588
rect 9332 62586 9356 62588
rect 9412 62586 9418 62588
rect 9172 62534 9174 62586
rect 9354 62534 9356 62586
rect 9110 62532 9116 62534
rect 9172 62532 9196 62534
rect 9252 62532 9276 62534
rect 9332 62532 9356 62534
rect 9412 62532 9418 62534
rect 9110 62512 9418 62532
rect 9110 61500 9418 61520
rect 9110 61498 9116 61500
rect 9172 61498 9196 61500
rect 9252 61498 9276 61500
rect 9332 61498 9356 61500
rect 9412 61498 9418 61500
rect 9172 61446 9174 61498
rect 9354 61446 9356 61498
rect 9110 61444 9116 61446
rect 9172 61444 9196 61446
rect 9252 61444 9276 61446
rect 9332 61444 9356 61446
rect 9412 61444 9418 61446
rect 9110 61424 9418 61444
rect 9110 60412 9418 60432
rect 9110 60410 9116 60412
rect 9172 60410 9196 60412
rect 9252 60410 9276 60412
rect 9332 60410 9356 60412
rect 9412 60410 9418 60412
rect 9172 60358 9174 60410
rect 9354 60358 9356 60410
rect 9110 60356 9116 60358
rect 9172 60356 9196 60358
rect 9252 60356 9276 60358
rect 9332 60356 9356 60358
rect 9412 60356 9418 60358
rect 9110 60336 9418 60356
rect 9312 59560 9364 59566
rect 9310 59528 9312 59537
rect 9364 59528 9366 59537
rect 9310 59463 9366 59472
rect 9110 59324 9418 59344
rect 9110 59322 9116 59324
rect 9172 59322 9196 59324
rect 9252 59322 9276 59324
rect 9332 59322 9356 59324
rect 9412 59322 9418 59324
rect 9172 59270 9174 59322
rect 9354 59270 9356 59322
rect 9110 59268 9116 59270
rect 9172 59268 9196 59270
rect 9252 59268 9276 59270
rect 9332 59268 9356 59270
rect 9412 59268 9418 59270
rect 9110 59248 9418 59268
rect 9600 58410 9628 63310
rect 9588 58404 9640 58410
rect 9588 58346 9640 58352
rect 9680 58336 9732 58342
rect 9680 58278 9732 58284
rect 9110 58236 9418 58256
rect 9110 58234 9116 58236
rect 9172 58234 9196 58236
rect 9252 58234 9276 58236
rect 9332 58234 9356 58236
rect 9412 58234 9418 58236
rect 9172 58182 9174 58234
rect 9354 58182 9356 58234
rect 9110 58180 9116 58182
rect 9172 58180 9196 58182
rect 9252 58180 9276 58182
rect 9332 58180 9356 58182
rect 9412 58180 9418 58182
rect 9110 58160 9418 58180
rect 9496 57384 9548 57390
rect 9496 57326 9548 57332
rect 9508 57225 9536 57326
rect 9494 57216 9550 57225
rect 9110 57148 9418 57168
rect 9494 57151 9550 57160
rect 9110 57146 9116 57148
rect 9172 57146 9196 57148
rect 9252 57146 9276 57148
rect 9332 57146 9356 57148
rect 9412 57146 9418 57148
rect 9172 57094 9174 57146
rect 9354 57094 9356 57146
rect 9110 57092 9116 57094
rect 9172 57092 9196 57094
rect 9252 57092 9276 57094
rect 9332 57092 9356 57094
rect 9412 57092 9418 57094
rect 9110 57072 9418 57092
rect 9312 56840 9364 56846
rect 9312 56782 9364 56788
rect 9324 56409 9352 56782
rect 9310 56400 9366 56409
rect 9310 56335 9366 56344
rect 8576 56296 8628 56302
rect 8576 56238 8628 56244
rect 8404 55916 8524 55944
rect 8300 54732 8352 54738
rect 8300 54674 8352 54680
rect 6644 54664 6696 54670
rect 6644 54606 6696 54612
rect 6552 50448 6604 50454
rect 6552 50390 6604 50396
rect 6460 49156 6512 49162
rect 6460 49098 6512 49104
rect 6460 47184 6512 47190
rect 6460 47126 6512 47132
rect 6368 43444 6420 43450
rect 6368 43386 6420 43392
rect 6288 43030 6408 43058
rect 6276 42764 6328 42770
rect 6276 42706 6328 42712
rect 6288 36242 6316 42706
rect 6380 41750 6408 43030
rect 6472 42786 6500 47126
rect 6552 47116 6604 47122
rect 6552 47058 6604 47064
rect 6564 46578 6592 47058
rect 6552 46572 6604 46578
rect 6552 46514 6604 46520
rect 6564 44810 6592 46514
rect 6552 44804 6604 44810
rect 6552 44746 6604 44752
rect 6564 44554 6592 44746
rect 6656 44742 6684 54606
rect 7478 54428 7786 54448
rect 7478 54426 7484 54428
rect 7540 54426 7564 54428
rect 7620 54426 7644 54428
rect 7700 54426 7724 54428
rect 7780 54426 7786 54428
rect 7540 54374 7542 54426
rect 7722 54374 7724 54426
rect 7478 54372 7484 54374
rect 7540 54372 7564 54374
rect 7620 54372 7644 54374
rect 7700 54372 7724 54374
rect 7780 54372 7786 54374
rect 7478 54352 7786 54372
rect 7478 53340 7786 53360
rect 7478 53338 7484 53340
rect 7540 53338 7564 53340
rect 7620 53338 7644 53340
rect 7700 53338 7724 53340
rect 7780 53338 7786 53340
rect 7540 53286 7542 53338
rect 7722 53286 7724 53338
rect 7478 53284 7484 53286
rect 7540 53284 7564 53286
rect 7620 53284 7644 53286
rect 7700 53284 7724 53286
rect 7780 53284 7786 53286
rect 7478 53264 7786 53284
rect 7478 52252 7786 52272
rect 7478 52250 7484 52252
rect 7540 52250 7564 52252
rect 7620 52250 7644 52252
rect 7700 52250 7724 52252
rect 7780 52250 7786 52252
rect 7540 52198 7542 52250
rect 7722 52198 7724 52250
rect 7478 52196 7484 52198
rect 7540 52196 7564 52198
rect 7620 52196 7644 52198
rect 7700 52196 7724 52198
rect 7780 52196 7786 52198
rect 7478 52176 7786 52196
rect 7478 51164 7786 51184
rect 7478 51162 7484 51164
rect 7540 51162 7564 51164
rect 7620 51162 7644 51164
rect 7700 51162 7724 51164
rect 7780 51162 7786 51164
rect 7540 51110 7542 51162
rect 7722 51110 7724 51162
rect 7478 51108 7484 51110
rect 7540 51108 7564 51110
rect 7620 51108 7644 51110
rect 7700 51108 7724 51110
rect 7780 51108 7786 51110
rect 7478 51088 7786 51108
rect 6736 51060 6788 51066
rect 6736 51002 6788 51008
rect 6644 44736 6696 44742
rect 6644 44678 6696 44684
rect 6564 44526 6684 44554
rect 6552 44396 6604 44402
rect 6552 44338 6604 44344
rect 6564 43994 6592 44338
rect 6552 43988 6604 43994
rect 6552 43930 6604 43936
rect 6656 43790 6684 44526
rect 6644 43784 6696 43790
rect 6644 43726 6696 43732
rect 6472 42758 6592 42786
rect 6460 42696 6512 42702
rect 6460 42638 6512 42644
rect 6368 41744 6420 41750
rect 6368 41686 6420 41692
rect 6368 41608 6420 41614
rect 6368 41550 6420 41556
rect 6380 39574 6408 41550
rect 6472 41274 6500 42638
rect 6564 41449 6592 42758
rect 6656 41546 6684 43726
rect 6644 41540 6696 41546
rect 6644 41482 6696 41488
rect 6550 41440 6606 41449
rect 6748 41414 6776 51002
rect 6828 50516 6880 50522
rect 6828 50458 6880 50464
rect 6550 41375 6606 41384
rect 6656 41386 6776 41414
rect 6460 41268 6512 41274
rect 6460 41210 6512 41216
rect 6460 41064 6512 41070
rect 6460 41006 6512 41012
rect 6368 39568 6420 39574
rect 6368 39510 6420 39516
rect 6472 38962 6500 41006
rect 6460 38956 6512 38962
rect 6460 38898 6512 38904
rect 6368 37188 6420 37194
rect 6368 37130 6420 37136
rect 6380 36922 6408 37130
rect 6368 36916 6420 36922
rect 6368 36858 6420 36864
rect 6552 36780 6604 36786
rect 6552 36722 6604 36728
rect 6460 36576 6512 36582
rect 6460 36518 6512 36524
rect 6276 36236 6328 36242
rect 6276 36178 6328 36184
rect 6276 35692 6328 35698
rect 6276 35634 6328 35640
rect 6288 33998 6316 35634
rect 6368 35624 6420 35630
rect 6368 35566 6420 35572
rect 6276 33992 6328 33998
rect 6276 33934 6328 33940
rect 6380 33862 6408 35566
rect 6368 33856 6420 33862
rect 6368 33798 6420 33804
rect 6184 31408 6236 31414
rect 6184 31350 6236 31356
rect 5846 31036 6154 31056
rect 5846 31034 5852 31036
rect 5908 31034 5932 31036
rect 5988 31034 6012 31036
rect 6068 31034 6092 31036
rect 6148 31034 6154 31036
rect 5908 30982 5910 31034
rect 6090 30982 6092 31034
rect 5846 30980 5852 30982
rect 5908 30980 5932 30982
rect 5988 30980 6012 30982
rect 6068 30980 6092 30982
rect 6148 30980 6154 30982
rect 5846 30960 6154 30980
rect 6472 30666 6500 36518
rect 6564 35834 6592 36722
rect 6656 36310 6684 41386
rect 6736 39432 6788 39438
rect 6736 39374 6788 39380
rect 6748 39098 6776 39374
rect 6736 39092 6788 39098
rect 6736 39034 6788 39040
rect 6840 36854 6868 50458
rect 7478 50076 7786 50096
rect 7478 50074 7484 50076
rect 7540 50074 7564 50076
rect 7620 50074 7644 50076
rect 7700 50074 7724 50076
rect 7780 50074 7786 50076
rect 7540 50022 7542 50074
rect 7722 50022 7724 50074
rect 7478 50020 7484 50022
rect 7540 50020 7564 50022
rect 7620 50020 7644 50022
rect 7700 50020 7724 50022
rect 7780 50020 7786 50022
rect 7478 50000 7786 50020
rect 7478 48988 7786 49008
rect 7478 48986 7484 48988
rect 7540 48986 7564 48988
rect 7620 48986 7644 48988
rect 7700 48986 7724 48988
rect 7780 48986 7786 48988
rect 7540 48934 7542 48986
rect 7722 48934 7724 48986
rect 7478 48932 7484 48934
rect 7540 48932 7564 48934
rect 7620 48932 7644 48934
rect 7700 48932 7724 48934
rect 7780 48932 7786 48934
rect 7478 48912 7786 48932
rect 7104 48204 7156 48210
rect 7104 48146 7156 48152
rect 7012 48068 7064 48074
rect 7012 48010 7064 48016
rect 6920 45960 6972 45966
rect 6920 45902 6972 45908
rect 6932 45354 6960 45902
rect 6920 45348 6972 45354
rect 6920 45290 6972 45296
rect 6920 43444 6972 43450
rect 6920 43386 6972 43392
rect 6932 41206 6960 43386
rect 7024 41478 7052 48010
rect 7012 41472 7064 41478
rect 7012 41414 7064 41420
rect 6920 41200 6972 41206
rect 6920 41142 6972 41148
rect 7012 41132 7064 41138
rect 7012 41074 7064 41080
rect 6920 40112 6972 40118
rect 6920 40054 6972 40060
rect 6932 39642 6960 40054
rect 6920 39636 6972 39642
rect 6920 39578 6972 39584
rect 7024 39574 7052 41074
rect 7012 39568 7064 39574
rect 7012 39510 7064 39516
rect 7116 38758 7144 48146
rect 7478 47900 7786 47920
rect 7478 47898 7484 47900
rect 7540 47898 7564 47900
rect 7620 47898 7644 47900
rect 7700 47898 7724 47900
rect 7780 47898 7786 47900
rect 7540 47846 7542 47898
rect 7722 47846 7724 47898
rect 7478 47844 7484 47846
rect 7540 47844 7564 47846
rect 7620 47844 7644 47846
rect 7700 47844 7724 47846
rect 7780 47844 7786 47846
rect 7478 47824 7786 47844
rect 8300 47660 8352 47666
rect 8300 47602 8352 47608
rect 7478 46812 7786 46832
rect 7478 46810 7484 46812
rect 7540 46810 7564 46812
rect 7620 46810 7644 46812
rect 7700 46810 7724 46812
rect 7780 46810 7786 46812
rect 7540 46758 7542 46810
rect 7722 46758 7724 46810
rect 7478 46756 7484 46758
rect 7540 46756 7564 46758
rect 7620 46756 7644 46758
rect 7700 46756 7724 46758
rect 7780 46756 7786 46758
rect 7478 46736 7786 46756
rect 8312 46714 8340 47602
rect 8300 46708 8352 46714
rect 8300 46650 8352 46656
rect 8116 46572 8168 46578
rect 8116 46514 8168 46520
rect 7478 45724 7786 45744
rect 7478 45722 7484 45724
rect 7540 45722 7564 45724
rect 7620 45722 7644 45724
rect 7700 45722 7724 45724
rect 7780 45722 7786 45724
rect 7540 45670 7542 45722
rect 7722 45670 7724 45722
rect 7478 45668 7484 45670
rect 7540 45668 7564 45670
rect 7620 45668 7644 45670
rect 7700 45668 7724 45670
rect 7780 45668 7786 45670
rect 7478 45648 7786 45668
rect 8128 45082 8156 46514
rect 8116 45076 8168 45082
rect 8116 45018 8168 45024
rect 7478 44636 7786 44656
rect 7478 44634 7484 44636
rect 7540 44634 7564 44636
rect 7620 44634 7644 44636
rect 7700 44634 7724 44636
rect 7780 44634 7786 44636
rect 7540 44582 7542 44634
rect 7722 44582 7724 44634
rect 7478 44580 7484 44582
rect 7540 44580 7564 44582
rect 7620 44580 7644 44582
rect 7700 44580 7724 44582
rect 7780 44580 7786 44582
rect 7478 44560 7786 44580
rect 7478 43548 7786 43568
rect 7478 43546 7484 43548
rect 7540 43546 7564 43548
rect 7620 43546 7644 43548
rect 7700 43546 7724 43548
rect 7780 43546 7786 43548
rect 7540 43494 7542 43546
rect 7722 43494 7724 43546
rect 7478 43492 7484 43494
rect 7540 43492 7564 43494
rect 7620 43492 7644 43494
rect 7700 43492 7724 43494
rect 7780 43492 7786 43494
rect 7478 43472 7786 43492
rect 8404 42770 8432 55916
rect 8588 51074 8616 56238
rect 9110 56060 9418 56080
rect 9110 56058 9116 56060
rect 9172 56058 9196 56060
rect 9252 56058 9276 56060
rect 9332 56058 9356 56060
rect 9412 56058 9418 56060
rect 9172 56006 9174 56058
rect 9354 56006 9356 56058
rect 9110 56004 9116 56006
rect 9172 56004 9196 56006
rect 9252 56004 9276 56006
rect 9332 56004 9356 56006
rect 9412 56004 9418 56006
rect 9110 55984 9418 56004
rect 9312 55752 9364 55758
rect 9310 55720 9312 55729
rect 9364 55720 9366 55729
rect 9310 55655 9366 55664
rect 9692 55418 9720 58278
rect 9680 55412 9732 55418
rect 9680 55354 9732 55360
rect 9496 55276 9548 55282
rect 9496 55218 9548 55224
rect 9110 54972 9418 54992
rect 9110 54970 9116 54972
rect 9172 54970 9196 54972
rect 9252 54970 9276 54972
rect 9332 54970 9356 54972
rect 9412 54970 9418 54972
rect 9172 54918 9174 54970
rect 9354 54918 9356 54970
rect 9110 54916 9116 54918
rect 9172 54916 9196 54918
rect 9252 54916 9276 54918
rect 9332 54916 9356 54918
rect 9412 54916 9418 54918
rect 9110 54896 9418 54916
rect 9508 54913 9536 55218
rect 9494 54904 9550 54913
rect 9494 54839 9550 54848
rect 9110 53884 9418 53904
rect 9110 53882 9116 53884
rect 9172 53882 9196 53884
rect 9252 53882 9276 53884
rect 9332 53882 9356 53884
rect 9412 53882 9418 53884
rect 9172 53830 9174 53882
rect 9354 53830 9356 53882
rect 9110 53828 9116 53830
rect 9172 53828 9196 53830
rect 9252 53828 9276 53830
rect 9332 53828 9356 53830
rect 9412 53828 9418 53830
rect 9110 53808 9418 53828
rect 9110 52796 9418 52816
rect 9110 52794 9116 52796
rect 9172 52794 9196 52796
rect 9252 52794 9276 52796
rect 9332 52794 9356 52796
rect 9412 52794 9418 52796
rect 9172 52742 9174 52794
rect 9354 52742 9356 52794
rect 9110 52740 9116 52742
rect 9172 52740 9196 52742
rect 9252 52740 9276 52742
rect 9332 52740 9356 52742
rect 9412 52740 9418 52742
rect 9110 52720 9418 52740
rect 9110 51708 9418 51728
rect 9110 51706 9116 51708
rect 9172 51706 9196 51708
rect 9252 51706 9276 51708
rect 9332 51706 9356 51708
rect 9412 51706 9418 51708
rect 9172 51654 9174 51706
rect 9354 51654 9356 51706
rect 9110 51652 9116 51654
rect 9172 51652 9196 51654
rect 9252 51652 9276 51654
rect 9332 51652 9356 51654
rect 9412 51652 9418 51654
rect 9110 51632 9418 51652
rect 8588 51046 8708 51074
rect 8484 48544 8536 48550
rect 8484 48486 8536 48492
rect 8392 42764 8444 42770
rect 8392 42706 8444 42712
rect 8496 42650 8524 48486
rect 8576 44940 8628 44946
rect 8576 44882 8628 44888
rect 8312 42622 8524 42650
rect 7478 42460 7786 42480
rect 7478 42458 7484 42460
rect 7540 42458 7564 42460
rect 7620 42458 7644 42460
rect 7700 42458 7724 42460
rect 7780 42458 7786 42460
rect 7540 42406 7542 42458
rect 7722 42406 7724 42458
rect 7478 42404 7484 42406
rect 7540 42404 7564 42406
rect 7620 42404 7644 42406
rect 7700 42404 7724 42406
rect 7780 42404 7786 42406
rect 7478 42384 7786 42404
rect 7478 41372 7786 41392
rect 7478 41370 7484 41372
rect 7540 41370 7564 41372
rect 7620 41370 7644 41372
rect 7700 41370 7724 41372
rect 7780 41370 7786 41372
rect 7540 41318 7542 41370
rect 7722 41318 7724 41370
rect 7478 41316 7484 41318
rect 7540 41316 7564 41318
rect 7620 41316 7644 41318
rect 7700 41316 7724 41318
rect 7780 41316 7786 41318
rect 7478 41296 7786 41316
rect 7478 40284 7786 40304
rect 7478 40282 7484 40284
rect 7540 40282 7564 40284
rect 7620 40282 7644 40284
rect 7700 40282 7724 40284
rect 7780 40282 7786 40284
rect 7540 40230 7542 40282
rect 7722 40230 7724 40282
rect 7478 40228 7484 40230
rect 7540 40228 7564 40230
rect 7620 40228 7644 40230
rect 7700 40228 7724 40230
rect 7780 40228 7786 40230
rect 7478 40208 7786 40228
rect 7478 39196 7786 39216
rect 7478 39194 7484 39196
rect 7540 39194 7564 39196
rect 7620 39194 7644 39196
rect 7700 39194 7724 39196
rect 7780 39194 7786 39196
rect 7540 39142 7542 39194
rect 7722 39142 7724 39194
rect 7478 39140 7484 39142
rect 7540 39140 7564 39142
rect 7620 39140 7644 39142
rect 7700 39140 7724 39142
rect 7780 39140 7786 39142
rect 7478 39120 7786 39140
rect 8208 38956 8260 38962
rect 8208 38898 8260 38904
rect 7104 38752 7156 38758
rect 7104 38694 7156 38700
rect 7478 38108 7786 38128
rect 7478 38106 7484 38108
rect 7540 38106 7564 38108
rect 7620 38106 7644 38108
rect 7700 38106 7724 38108
rect 7780 38106 7786 38108
rect 7540 38054 7542 38106
rect 7722 38054 7724 38106
rect 7478 38052 7484 38054
rect 7540 38052 7564 38054
rect 7620 38052 7644 38054
rect 7700 38052 7724 38054
rect 7780 38052 7786 38054
rect 7478 38032 7786 38052
rect 8220 37126 8248 38898
rect 8208 37120 8260 37126
rect 8208 37062 8260 37068
rect 7478 37020 7786 37040
rect 7478 37018 7484 37020
rect 7540 37018 7564 37020
rect 7620 37018 7644 37020
rect 7700 37018 7724 37020
rect 7780 37018 7786 37020
rect 7540 36966 7542 37018
rect 7722 36966 7724 37018
rect 7478 36964 7484 36966
rect 7540 36964 7564 36966
rect 7620 36964 7644 36966
rect 7700 36964 7724 36966
rect 7780 36964 7786 36966
rect 7478 36944 7786 36964
rect 6828 36848 6880 36854
rect 6828 36790 6880 36796
rect 7196 36780 7248 36786
rect 7196 36722 7248 36728
rect 6644 36304 6696 36310
rect 6644 36246 6696 36252
rect 7208 35834 7236 36722
rect 7478 35932 7786 35952
rect 7478 35930 7484 35932
rect 7540 35930 7564 35932
rect 7620 35930 7644 35932
rect 7700 35930 7724 35932
rect 7780 35930 7786 35932
rect 7540 35878 7542 35930
rect 7722 35878 7724 35930
rect 7478 35876 7484 35878
rect 7540 35876 7564 35878
rect 7620 35876 7644 35878
rect 7700 35876 7724 35878
rect 7780 35876 7786 35878
rect 7478 35856 7786 35876
rect 6552 35828 6604 35834
rect 6552 35770 6604 35776
rect 7196 35828 7248 35834
rect 7196 35770 7248 35776
rect 7478 34844 7786 34864
rect 7478 34842 7484 34844
rect 7540 34842 7564 34844
rect 7620 34842 7644 34844
rect 7700 34842 7724 34844
rect 7780 34842 7786 34844
rect 7540 34790 7542 34842
rect 7722 34790 7724 34842
rect 7478 34788 7484 34790
rect 7540 34788 7564 34790
rect 7620 34788 7644 34790
rect 7700 34788 7724 34790
rect 7780 34788 7786 34790
rect 7478 34768 7786 34788
rect 7478 33756 7786 33776
rect 7478 33754 7484 33756
rect 7540 33754 7564 33756
rect 7620 33754 7644 33756
rect 7700 33754 7724 33756
rect 7780 33754 7786 33756
rect 7540 33702 7542 33754
rect 7722 33702 7724 33754
rect 7478 33700 7484 33702
rect 7540 33700 7564 33702
rect 7620 33700 7644 33702
rect 7700 33700 7724 33702
rect 7780 33700 7786 33702
rect 7478 33680 7786 33700
rect 7840 32904 7892 32910
rect 7840 32846 7892 32852
rect 7478 32668 7786 32688
rect 7478 32666 7484 32668
rect 7540 32666 7564 32668
rect 7620 32666 7644 32668
rect 7700 32666 7724 32668
rect 7780 32666 7786 32668
rect 7540 32614 7542 32666
rect 7722 32614 7724 32666
rect 7478 32612 7484 32614
rect 7540 32612 7564 32614
rect 7620 32612 7644 32614
rect 7700 32612 7724 32614
rect 7780 32612 7786 32614
rect 7478 32592 7786 32612
rect 7478 31580 7786 31600
rect 7478 31578 7484 31580
rect 7540 31578 7564 31580
rect 7620 31578 7644 31580
rect 7700 31578 7724 31580
rect 7780 31578 7786 31580
rect 7540 31526 7542 31578
rect 7722 31526 7724 31578
rect 7478 31524 7484 31526
rect 7540 31524 7564 31526
rect 7620 31524 7644 31526
rect 7700 31524 7724 31526
rect 7780 31524 7786 31526
rect 7478 31504 7786 31524
rect 6460 30660 6512 30666
rect 6460 30602 6512 30608
rect 7478 30492 7786 30512
rect 7478 30490 7484 30492
rect 7540 30490 7564 30492
rect 7620 30490 7644 30492
rect 7700 30490 7724 30492
rect 7780 30490 7786 30492
rect 7540 30438 7542 30490
rect 7722 30438 7724 30490
rect 7478 30436 7484 30438
rect 7540 30436 7564 30438
rect 7620 30436 7644 30438
rect 7700 30436 7724 30438
rect 7780 30436 7786 30438
rect 7478 30416 7786 30436
rect 5846 29948 6154 29968
rect 5846 29946 5852 29948
rect 5908 29946 5932 29948
rect 5988 29946 6012 29948
rect 6068 29946 6092 29948
rect 6148 29946 6154 29948
rect 5908 29894 5910 29946
rect 6090 29894 6092 29946
rect 5846 29892 5852 29894
rect 5908 29892 5932 29894
rect 5988 29892 6012 29894
rect 6068 29892 6092 29894
rect 6148 29892 6154 29894
rect 5846 29872 6154 29892
rect 7478 29404 7786 29424
rect 7478 29402 7484 29404
rect 7540 29402 7564 29404
rect 7620 29402 7644 29404
rect 7700 29402 7724 29404
rect 7780 29402 7786 29404
rect 7540 29350 7542 29402
rect 7722 29350 7724 29402
rect 7478 29348 7484 29350
rect 7540 29348 7564 29350
rect 7620 29348 7644 29350
rect 7700 29348 7724 29350
rect 7780 29348 7786 29350
rect 7478 29328 7786 29348
rect 5846 28860 6154 28880
rect 5846 28858 5852 28860
rect 5908 28858 5932 28860
rect 5988 28858 6012 28860
rect 6068 28858 6092 28860
rect 6148 28858 6154 28860
rect 5908 28806 5910 28858
rect 6090 28806 6092 28858
rect 5846 28804 5852 28806
rect 5908 28804 5932 28806
rect 5988 28804 6012 28806
rect 6068 28804 6092 28806
rect 6148 28804 6154 28806
rect 5846 28784 6154 28804
rect 7478 28316 7786 28336
rect 7478 28314 7484 28316
rect 7540 28314 7564 28316
rect 7620 28314 7644 28316
rect 7700 28314 7724 28316
rect 7780 28314 7786 28316
rect 7540 28262 7542 28314
rect 7722 28262 7724 28314
rect 7478 28260 7484 28262
rect 7540 28260 7564 28262
rect 7620 28260 7644 28262
rect 7700 28260 7724 28262
rect 7780 28260 7786 28262
rect 7478 28240 7786 28260
rect 5846 27772 6154 27792
rect 5846 27770 5852 27772
rect 5908 27770 5932 27772
rect 5988 27770 6012 27772
rect 6068 27770 6092 27772
rect 6148 27770 6154 27772
rect 5908 27718 5910 27770
rect 6090 27718 6092 27770
rect 5846 27716 5852 27718
rect 5908 27716 5932 27718
rect 5988 27716 6012 27718
rect 6068 27716 6092 27718
rect 6148 27716 6154 27718
rect 5846 27696 6154 27716
rect 7478 27228 7786 27248
rect 7478 27226 7484 27228
rect 7540 27226 7564 27228
rect 7620 27226 7644 27228
rect 7700 27226 7724 27228
rect 7780 27226 7786 27228
rect 7540 27174 7542 27226
rect 7722 27174 7724 27226
rect 7478 27172 7484 27174
rect 7540 27172 7564 27174
rect 7620 27172 7644 27174
rect 7700 27172 7724 27174
rect 7780 27172 7786 27174
rect 7478 27152 7786 27172
rect 5846 26684 6154 26704
rect 5846 26682 5852 26684
rect 5908 26682 5932 26684
rect 5988 26682 6012 26684
rect 6068 26682 6092 26684
rect 6148 26682 6154 26684
rect 5908 26630 5910 26682
rect 6090 26630 6092 26682
rect 5846 26628 5852 26630
rect 5908 26628 5932 26630
rect 5988 26628 6012 26630
rect 6068 26628 6092 26630
rect 6148 26628 6154 26630
rect 5846 26608 6154 26628
rect 7478 26140 7786 26160
rect 7478 26138 7484 26140
rect 7540 26138 7564 26140
rect 7620 26138 7644 26140
rect 7700 26138 7724 26140
rect 7780 26138 7786 26140
rect 7540 26086 7542 26138
rect 7722 26086 7724 26138
rect 7478 26084 7484 26086
rect 7540 26084 7564 26086
rect 7620 26084 7644 26086
rect 7700 26084 7724 26086
rect 7780 26084 7786 26086
rect 7478 26064 7786 26084
rect 5846 25596 6154 25616
rect 5846 25594 5852 25596
rect 5908 25594 5932 25596
rect 5988 25594 6012 25596
rect 6068 25594 6092 25596
rect 6148 25594 6154 25596
rect 5908 25542 5910 25594
rect 6090 25542 6092 25594
rect 5846 25540 5852 25542
rect 5908 25540 5932 25542
rect 5988 25540 6012 25542
rect 6068 25540 6092 25542
rect 6148 25540 6154 25542
rect 5846 25520 6154 25540
rect 7478 25052 7786 25072
rect 7478 25050 7484 25052
rect 7540 25050 7564 25052
rect 7620 25050 7644 25052
rect 7700 25050 7724 25052
rect 7780 25050 7786 25052
rect 7540 24998 7542 25050
rect 7722 24998 7724 25050
rect 7478 24996 7484 24998
rect 7540 24996 7564 24998
rect 7620 24996 7644 24998
rect 7700 24996 7724 24998
rect 7780 24996 7786 24998
rect 7478 24976 7786 24996
rect 5846 24508 6154 24528
rect 5846 24506 5852 24508
rect 5908 24506 5932 24508
rect 5988 24506 6012 24508
rect 6068 24506 6092 24508
rect 6148 24506 6154 24508
rect 5908 24454 5910 24506
rect 6090 24454 6092 24506
rect 5846 24452 5852 24454
rect 5908 24452 5932 24454
rect 5988 24452 6012 24454
rect 6068 24452 6092 24454
rect 6148 24452 6154 24454
rect 5846 24432 6154 24452
rect 7852 24274 7880 32846
rect 7932 31816 7984 31822
rect 7932 31758 7984 31764
rect 7840 24268 7892 24274
rect 7840 24210 7892 24216
rect 7478 23964 7786 23984
rect 7478 23962 7484 23964
rect 7540 23962 7564 23964
rect 7620 23962 7644 23964
rect 7700 23962 7724 23964
rect 7780 23962 7786 23964
rect 7540 23910 7542 23962
rect 7722 23910 7724 23962
rect 7478 23908 7484 23910
rect 7540 23908 7564 23910
rect 7620 23908 7644 23910
rect 7700 23908 7724 23910
rect 7780 23908 7786 23910
rect 7478 23888 7786 23908
rect 7944 23662 7972 31758
rect 7932 23656 7984 23662
rect 7932 23598 7984 23604
rect 5846 23420 6154 23440
rect 5846 23418 5852 23420
rect 5908 23418 5932 23420
rect 5988 23418 6012 23420
rect 6068 23418 6092 23420
rect 6148 23418 6154 23420
rect 5908 23366 5910 23418
rect 6090 23366 6092 23418
rect 5846 23364 5852 23366
rect 5908 23364 5932 23366
rect 5988 23364 6012 23366
rect 6068 23364 6092 23366
rect 6148 23364 6154 23366
rect 5846 23344 6154 23364
rect 5724 23248 5776 23254
rect 5724 23190 5776 23196
rect 7478 22876 7786 22896
rect 7478 22874 7484 22876
rect 7540 22874 7564 22876
rect 7620 22874 7644 22876
rect 7700 22874 7724 22876
rect 7780 22874 7786 22876
rect 7540 22822 7542 22874
rect 7722 22822 7724 22874
rect 7478 22820 7484 22822
rect 7540 22820 7564 22822
rect 7620 22820 7644 22822
rect 7700 22820 7724 22822
rect 7780 22820 7786 22822
rect 7478 22800 7786 22820
rect 5846 22332 6154 22352
rect 5846 22330 5852 22332
rect 5908 22330 5932 22332
rect 5988 22330 6012 22332
rect 6068 22330 6092 22332
rect 6148 22330 6154 22332
rect 5908 22278 5910 22330
rect 6090 22278 6092 22330
rect 5846 22276 5852 22278
rect 5908 22276 5932 22278
rect 5988 22276 6012 22278
rect 6068 22276 6092 22278
rect 6148 22276 6154 22278
rect 5846 22256 6154 22276
rect 7478 21788 7786 21808
rect 7478 21786 7484 21788
rect 7540 21786 7564 21788
rect 7620 21786 7644 21788
rect 7700 21786 7724 21788
rect 7780 21786 7786 21788
rect 7540 21734 7542 21786
rect 7722 21734 7724 21786
rect 7478 21732 7484 21734
rect 7540 21732 7564 21734
rect 7620 21732 7644 21734
rect 7700 21732 7724 21734
rect 7780 21732 7786 21734
rect 7478 21712 7786 21732
rect 5448 21616 5500 21622
rect 5448 21558 5500 21564
rect 5846 21244 6154 21264
rect 5846 21242 5852 21244
rect 5908 21242 5932 21244
rect 5988 21242 6012 21244
rect 6068 21242 6092 21244
rect 6148 21242 6154 21244
rect 5908 21190 5910 21242
rect 6090 21190 6092 21242
rect 5846 21188 5852 21190
rect 5908 21188 5932 21190
rect 5988 21188 6012 21190
rect 6068 21188 6092 21190
rect 6148 21188 6154 21190
rect 5846 21168 6154 21188
rect 7478 20700 7786 20720
rect 7478 20698 7484 20700
rect 7540 20698 7564 20700
rect 7620 20698 7644 20700
rect 7700 20698 7724 20700
rect 7780 20698 7786 20700
rect 7540 20646 7542 20698
rect 7722 20646 7724 20698
rect 7478 20644 7484 20646
rect 7540 20644 7564 20646
rect 7620 20644 7644 20646
rect 7700 20644 7724 20646
rect 7780 20644 7786 20646
rect 7478 20624 7786 20644
rect 5846 20156 6154 20176
rect 5846 20154 5852 20156
rect 5908 20154 5932 20156
rect 5988 20154 6012 20156
rect 6068 20154 6092 20156
rect 6148 20154 6154 20156
rect 5908 20102 5910 20154
rect 6090 20102 6092 20154
rect 5846 20100 5852 20102
rect 5908 20100 5932 20102
rect 5988 20100 6012 20102
rect 6068 20100 6092 20102
rect 6148 20100 6154 20102
rect 5846 20080 6154 20100
rect 7478 19612 7786 19632
rect 7478 19610 7484 19612
rect 7540 19610 7564 19612
rect 7620 19610 7644 19612
rect 7700 19610 7724 19612
rect 7780 19610 7786 19612
rect 7540 19558 7542 19610
rect 7722 19558 7724 19610
rect 7478 19556 7484 19558
rect 7540 19556 7564 19558
rect 7620 19556 7644 19558
rect 7700 19556 7724 19558
rect 7780 19556 7786 19558
rect 7478 19536 7786 19556
rect 5846 19068 6154 19088
rect 5846 19066 5852 19068
rect 5908 19066 5932 19068
rect 5988 19066 6012 19068
rect 6068 19066 6092 19068
rect 6148 19066 6154 19068
rect 5908 19014 5910 19066
rect 6090 19014 6092 19066
rect 5846 19012 5852 19014
rect 5908 19012 5932 19014
rect 5988 19012 6012 19014
rect 6068 19012 6092 19014
rect 6148 19012 6154 19014
rect 5846 18992 6154 19012
rect 7478 18524 7786 18544
rect 7478 18522 7484 18524
rect 7540 18522 7564 18524
rect 7620 18522 7644 18524
rect 7700 18522 7724 18524
rect 7780 18522 7786 18524
rect 7540 18470 7542 18522
rect 7722 18470 7724 18522
rect 7478 18468 7484 18470
rect 7540 18468 7564 18470
rect 7620 18468 7644 18470
rect 7700 18468 7724 18470
rect 7780 18468 7786 18470
rect 7478 18448 7786 18468
rect 5846 17980 6154 18000
rect 5846 17978 5852 17980
rect 5908 17978 5932 17980
rect 5988 17978 6012 17980
rect 6068 17978 6092 17980
rect 6148 17978 6154 17980
rect 5908 17926 5910 17978
rect 6090 17926 6092 17978
rect 5846 17924 5852 17926
rect 5908 17924 5932 17926
rect 5988 17924 6012 17926
rect 6068 17924 6092 17926
rect 6148 17924 6154 17926
rect 5846 17904 6154 17924
rect 7478 17436 7786 17456
rect 7478 17434 7484 17436
rect 7540 17434 7564 17436
rect 7620 17434 7644 17436
rect 7700 17434 7724 17436
rect 7780 17434 7786 17436
rect 7540 17382 7542 17434
rect 7722 17382 7724 17434
rect 7478 17380 7484 17382
rect 7540 17380 7564 17382
rect 7620 17380 7644 17382
rect 7700 17380 7724 17382
rect 7780 17380 7786 17382
rect 7478 17360 7786 17380
rect 5846 16892 6154 16912
rect 5846 16890 5852 16892
rect 5908 16890 5932 16892
rect 5988 16890 6012 16892
rect 6068 16890 6092 16892
rect 6148 16890 6154 16892
rect 5908 16838 5910 16890
rect 6090 16838 6092 16890
rect 5846 16836 5852 16838
rect 5908 16836 5932 16838
rect 5988 16836 6012 16838
rect 6068 16836 6092 16838
rect 6148 16836 6154 16838
rect 5846 16816 6154 16836
rect 7478 16348 7786 16368
rect 7478 16346 7484 16348
rect 7540 16346 7564 16348
rect 7620 16346 7644 16348
rect 7700 16346 7724 16348
rect 7780 16346 7786 16348
rect 7540 16294 7542 16346
rect 7722 16294 7724 16346
rect 7478 16292 7484 16294
rect 7540 16292 7564 16294
rect 7620 16292 7644 16294
rect 7700 16292 7724 16294
rect 7780 16292 7786 16294
rect 7478 16272 7786 16292
rect 5846 15804 6154 15824
rect 5846 15802 5852 15804
rect 5908 15802 5932 15804
rect 5988 15802 6012 15804
rect 6068 15802 6092 15804
rect 6148 15802 6154 15804
rect 5908 15750 5910 15802
rect 6090 15750 6092 15802
rect 5846 15748 5852 15750
rect 5908 15748 5932 15750
rect 5988 15748 6012 15750
rect 6068 15748 6092 15750
rect 6148 15748 6154 15750
rect 5846 15728 6154 15748
rect 7478 15260 7786 15280
rect 7478 15258 7484 15260
rect 7540 15258 7564 15260
rect 7620 15258 7644 15260
rect 7700 15258 7724 15260
rect 7780 15258 7786 15260
rect 7540 15206 7542 15258
rect 7722 15206 7724 15258
rect 7478 15204 7484 15206
rect 7540 15204 7564 15206
rect 7620 15204 7644 15206
rect 7700 15204 7724 15206
rect 7780 15204 7786 15206
rect 7478 15184 7786 15204
rect 5846 14716 6154 14736
rect 5846 14714 5852 14716
rect 5908 14714 5932 14716
rect 5988 14714 6012 14716
rect 6068 14714 6092 14716
rect 6148 14714 6154 14716
rect 5908 14662 5910 14714
rect 6090 14662 6092 14714
rect 5846 14660 5852 14662
rect 5908 14660 5932 14662
rect 5988 14660 6012 14662
rect 6068 14660 6092 14662
rect 6148 14660 6154 14662
rect 5846 14640 6154 14660
rect 7478 14172 7786 14192
rect 7478 14170 7484 14172
rect 7540 14170 7564 14172
rect 7620 14170 7644 14172
rect 7700 14170 7724 14172
rect 7780 14170 7786 14172
rect 7540 14118 7542 14170
rect 7722 14118 7724 14170
rect 7478 14116 7484 14118
rect 7540 14116 7564 14118
rect 7620 14116 7644 14118
rect 7700 14116 7724 14118
rect 7780 14116 7786 14118
rect 7478 14096 7786 14116
rect 5846 13628 6154 13648
rect 5846 13626 5852 13628
rect 5908 13626 5932 13628
rect 5988 13626 6012 13628
rect 6068 13626 6092 13628
rect 6148 13626 6154 13628
rect 5908 13574 5910 13626
rect 6090 13574 6092 13626
rect 5846 13572 5852 13574
rect 5908 13572 5932 13574
rect 5988 13572 6012 13574
rect 6068 13572 6092 13574
rect 6148 13572 6154 13574
rect 5846 13552 6154 13572
rect 7478 13084 7786 13104
rect 7478 13082 7484 13084
rect 7540 13082 7564 13084
rect 7620 13082 7644 13084
rect 7700 13082 7724 13084
rect 7780 13082 7786 13084
rect 7540 13030 7542 13082
rect 7722 13030 7724 13082
rect 7478 13028 7484 13030
rect 7540 13028 7564 13030
rect 7620 13028 7644 13030
rect 7700 13028 7724 13030
rect 7780 13028 7786 13030
rect 7478 13008 7786 13028
rect 5846 12540 6154 12560
rect 5846 12538 5852 12540
rect 5908 12538 5932 12540
rect 5988 12538 6012 12540
rect 6068 12538 6092 12540
rect 6148 12538 6154 12540
rect 5908 12486 5910 12538
rect 6090 12486 6092 12538
rect 5846 12484 5852 12486
rect 5908 12484 5932 12486
rect 5988 12484 6012 12486
rect 6068 12484 6092 12486
rect 6148 12484 6154 12486
rect 5846 12464 6154 12484
rect 7478 11996 7786 12016
rect 7478 11994 7484 11996
rect 7540 11994 7564 11996
rect 7620 11994 7644 11996
rect 7700 11994 7724 11996
rect 7780 11994 7786 11996
rect 7540 11942 7542 11994
rect 7722 11942 7724 11994
rect 7478 11940 7484 11942
rect 7540 11940 7564 11942
rect 7620 11940 7644 11942
rect 7700 11940 7724 11942
rect 7780 11940 7786 11942
rect 7478 11920 7786 11940
rect 5846 11452 6154 11472
rect 5846 11450 5852 11452
rect 5908 11450 5932 11452
rect 5988 11450 6012 11452
rect 6068 11450 6092 11452
rect 6148 11450 6154 11452
rect 5908 11398 5910 11450
rect 6090 11398 6092 11450
rect 5846 11396 5852 11398
rect 5908 11396 5932 11398
rect 5988 11396 6012 11398
rect 6068 11396 6092 11398
rect 6148 11396 6154 11398
rect 5846 11376 6154 11396
rect 7478 10908 7786 10928
rect 7478 10906 7484 10908
rect 7540 10906 7564 10908
rect 7620 10906 7644 10908
rect 7700 10906 7724 10908
rect 7780 10906 7786 10908
rect 7540 10854 7542 10906
rect 7722 10854 7724 10906
rect 7478 10852 7484 10854
rect 7540 10852 7564 10854
rect 7620 10852 7644 10854
rect 7700 10852 7724 10854
rect 7780 10852 7786 10854
rect 7478 10832 7786 10852
rect 5846 10364 6154 10384
rect 5846 10362 5852 10364
rect 5908 10362 5932 10364
rect 5988 10362 6012 10364
rect 6068 10362 6092 10364
rect 6148 10362 6154 10364
rect 5908 10310 5910 10362
rect 6090 10310 6092 10362
rect 5846 10308 5852 10310
rect 5908 10308 5932 10310
rect 5988 10308 6012 10310
rect 6068 10308 6092 10310
rect 6148 10308 6154 10310
rect 5846 10288 6154 10308
rect 7478 9820 7786 9840
rect 7478 9818 7484 9820
rect 7540 9818 7564 9820
rect 7620 9818 7644 9820
rect 7700 9818 7724 9820
rect 7780 9818 7786 9820
rect 7540 9766 7542 9818
rect 7722 9766 7724 9818
rect 7478 9764 7484 9766
rect 7540 9764 7564 9766
rect 7620 9764 7644 9766
rect 7700 9764 7724 9766
rect 7780 9764 7786 9766
rect 7478 9744 7786 9764
rect 8312 9382 8340 42622
rect 8588 41414 8616 44882
rect 8404 41386 8616 41414
rect 8404 31754 8432 41386
rect 8484 38344 8536 38350
rect 8484 38286 8536 38292
rect 8496 36922 8524 38286
rect 8576 37256 8628 37262
rect 8576 37198 8628 37204
rect 8484 36916 8536 36922
rect 8484 36858 8536 36864
rect 8588 34202 8616 37198
rect 8576 34196 8628 34202
rect 8576 34138 8628 34144
rect 8404 31726 8616 31754
rect 8392 30728 8444 30734
rect 8392 30670 8444 30676
rect 8404 29850 8432 30670
rect 8392 29844 8444 29850
rect 8392 29786 8444 29792
rect 8588 15162 8616 31726
rect 8680 30190 8708 51046
rect 9110 50620 9418 50640
rect 9110 50618 9116 50620
rect 9172 50618 9196 50620
rect 9252 50618 9276 50620
rect 9332 50618 9356 50620
rect 9412 50618 9418 50620
rect 9172 50566 9174 50618
rect 9354 50566 9356 50618
rect 9110 50564 9116 50566
rect 9172 50564 9196 50566
rect 9252 50564 9276 50566
rect 9332 50564 9356 50566
rect 9412 50564 9418 50566
rect 9110 50544 9418 50564
rect 9588 49972 9640 49978
rect 9588 49914 9640 49920
rect 9110 49532 9418 49552
rect 9110 49530 9116 49532
rect 9172 49530 9196 49532
rect 9252 49530 9276 49532
rect 9332 49530 9356 49532
rect 9412 49530 9418 49532
rect 9172 49478 9174 49530
rect 9354 49478 9356 49530
rect 9110 49476 9116 49478
rect 9172 49476 9196 49478
rect 9252 49476 9276 49478
rect 9332 49476 9356 49478
rect 9412 49476 9418 49478
rect 9110 49456 9418 49476
rect 9600 49473 9628 49914
rect 9680 49836 9732 49842
rect 9680 49778 9732 49784
rect 9586 49464 9642 49473
rect 9586 49399 9642 49408
rect 9110 48444 9418 48464
rect 9110 48442 9116 48444
rect 9172 48442 9196 48444
rect 9252 48442 9276 48444
rect 9332 48442 9356 48444
rect 9412 48442 9418 48444
rect 9172 48390 9174 48442
rect 9354 48390 9356 48442
rect 9110 48388 9116 48390
rect 9172 48388 9196 48390
rect 9252 48388 9276 48390
rect 9332 48388 9356 48390
rect 9412 48388 9418 48390
rect 9110 48368 9418 48388
rect 9692 48278 9720 49778
rect 9680 48272 9732 48278
rect 9680 48214 9732 48220
rect 9496 48136 9548 48142
rect 9496 48078 9548 48084
rect 9110 47356 9418 47376
rect 9110 47354 9116 47356
rect 9172 47354 9196 47356
rect 9252 47354 9276 47356
rect 9332 47354 9356 47356
rect 9412 47354 9418 47356
rect 9172 47302 9174 47354
rect 9354 47302 9356 47354
rect 9110 47300 9116 47302
rect 9172 47300 9196 47302
rect 9252 47300 9276 47302
rect 9332 47300 9356 47302
rect 9412 47300 9418 47302
rect 9110 47280 9418 47300
rect 9508 47258 9536 48078
rect 9496 47252 9548 47258
rect 9496 47194 9548 47200
rect 9110 46268 9418 46288
rect 9110 46266 9116 46268
rect 9172 46266 9196 46268
rect 9252 46266 9276 46268
rect 9332 46266 9356 46268
rect 9412 46266 9418 46268
rect 9172 46214 9174 46266
rect 9354 46214 9356 46266
rect 9110 46212 9116 46214
rect 9172 46212 9196 46214
rect 9252 46212 9276 46214
rect 9332 46212 9356 46214
rect 9412 46212 9418 46214
rect 9110 46192 9418 46212
rect 9110 45180 9418 45200
rect 9110 45178 9116 45180
rect 9172 45178 9196 45180
rect 9252 45178 9276 45180
rect 9332 45178 9356 45180
rect 9412 45178 9418 45180
rect 9172 45126 9174 45178
rect 9354 45126 9356 45178
rect 9110 45124 9116 45126
rect 9172 45124 9196 45126
rect 9252 45124 9276 45126
rect 9332 45124 9356 45126
rect 9412 45124 9418 45126
rect 9110 45104 9418 45124
rect 9110 44092 9418 44112
rect 9110 44090 9116 44092
rect 9172 44090 9196 44092
rect 9252 44090 9276 44092
rect 9332 44090 9356 44092
rect 9412 44090 9418 44092
rect 9172 44038 9174 44090
rect 9354 44038 9356 44090
rect 9110 44036 9116 44038
rect 9172 44036 9196 44038
rect 9252 44036 9276 44038
rect 9332 44036 9356 44038
rect 9412 44036 9418 44038
rect 9110 44016 9418 44036
rect 9680 43308 9732 43314
rect 9680 43250 9732 43256
rect 9110 43004 9418 43024
rect 9110 43002 9116 43004
rect 9172 43002 9196 43004
rect 9252 43002 9276 43004
rect 9332 43002 9356 43004
rect 9412 43002 9418 43004
rect 9172 42950 9174 43002
rect 9354 42950 9356 43002
rect 9110 42948 9116 42950
rect 9172 42948 9196 42950
rect 9252 42948 9276 42950
rect 9332 42948 9356 42950
rect 9412 42948 9418 42950
rect 9110 42928 9418 42948
rect 9496 42220 9548 42226
rect 9496 42162 9548 42168
rect 9110 41916 9418 41936
rect 9110 41914 9116 41916
rect 9172 41914 9196 41916
rect 9252 41914 9276 41916
rect 9332 41914 9356 41916
rect 9412 41914 9418 41916
rect 9172 41862 9174 41914
rect 9354 41862 9356 41914
rect 9110 41860 9116 41862
rect 9172 41860 9196 41862
rect 9252 41860 9276 41862
rect 9332 41860 9356 41862
rect 9412 41860 9418 41862
rect 9110 41840 9418 41860
rect 9110 40828 9418 40848
rect 9110 40826 9116 40828
rect 9172 40826 9196 40828
rect 9252 40826 9276 40828
rect 9332 40826 9356 40828
rect 9412 40826 9418 40828
rect 9172 40774 9174 40826
rect 9354 40774 9356 40826
rect 9110 40772 9116 40774
rect 9172 40772 9196 40774
rect 9252 40772 9276 40774
rect 9332 40772 9356 40774
rect 9412 40772 9418 40774
rect 9110 40752 9418 40772
rect 9508 40730 9536 42162
rect 9692 41818 9720 43250
rect 9784 43246 9812 76774
rect 10140 76424 10192 76430
rect 10138 76392 10140 76401
rect 10192 76392 10194 76401
rect 10138 76327 10194 76336
rect 10140 75948 10192 75954
rect 10140 75890 10192 75896
rect 10152 75721 10180 75890
rect 10138 75712 10194 75721
rect 10138 75647 10194 75656
rect 10140 75336 10192 75342
rect 10140 75278 10192 75284
rect 10152 74905 10180 75278
rect 10138 74896 10194 74905
rect 10138 74831 10194 74840
rect 10140 74248 10192 74254
rect 10140 74190 10192 74196
rect 10152 74089 10180 74190
rect 10138 74080 10194 74089
rect 10138 74015 10194 74024
rect 10140 73772 10192 73778
rect 10140 73714 10192 73720
rect 10152 73409 10180 73714
rect 10138 73400 10194 73409
rect 10138 73335 10194 73344
rect 9956 73160 10008 73166
rect 9956 73102 10008 73108
rect 9968 72282 9996 73102
rect 10140 72684 10192 72690
rect 10140 72626 10192 72632
rect 10152 72593 10180 72626
rect 10138 72584 10194 72593
rect 10138 72519 10194 72528
rect 9956 72276 10008 72282
rect 9956 72218 10008 72224
rect 10140 72072 10192 72078
rect 10140 72014 10192 72020
rect 10152 71777 10180 72014
rect 10138 71768 10194 71777
rect 10138 71703 10194 71712
rect 10140 71596 10192 71602
rect 10140 71538 10192 71544
rect 10152 71097 10180 71538
rect 10138 71088 10194 71097
rect 10138 71023 10194 71032
rect 10140 70508 10192 70514
rect 10140 70450 10192 70456
rect 10152 70281 10180 70450
rect 10138 70272 10194 70281
rect 10138 70207 10194 70216
rect 10140 69896 10192 69902
rect 10140 69838 10192 69844
rect 9956 69760 10008 69766
rect 9956 69702 10008 69708
rect 9968 68882 9996 69702
rect 10152 69465 10180 69838
rect 10138 69456 10194 69465
rect 10138 69391 10194 69400
rect 9956 68876 10008 68882
rect 9956 68818 10008 68824
rect 10140 68808 10192 68814
rect 10138 68776 10140 68785
rect 10192 68776 10194 68785
rect 10138 68711 10194 68720
rect 9956 68672 10008 68678
rect 9956 68614 10008 68620
rect 9968 68270 9996 68614
rect 10140 68332 10192 68338
rect 10140 68274 10192 68280
rect 9956 68264 10008 68270
rect 9956 68206 10008 68212
rect 9864 68128 9916 68134
rect 9864 68070 9916 68076
rect 9876 66094 9904 68070
rect 10152 67969 10180 68274
rect 10138 67960 10194 67969
rect 10138 67895 10194 67904
rect 9956 67788 10008 67794
rect 9956 67730 10008 67736
rect 9968 67386 9996 67730
rect 9956 67380 10008 67386
rect 9956 67322 10008 67328
rect 10140 67244 10192 67250
rect 10140 67186 10192 67192
rect 10152 67153 10180 67186
rect 10138 67144 10194 67153
rect 10138 67079 10194 67088
rect 10140 66632 10192 66638
rect 10140 66574 10192 66580
rect 10152 66473 10180 66574
rect 10138 66464 10194 66473
rect 10138 66399 10194 66408
rect 10140 66156 10192 66162
rect 10140 66098 10192 66104
rect 9864 66088 9916 66094
rect 9864 66030 9916 66036
rect 10152 65657 10180 66098
rect 10138 65648 10194 65657
rect 10138 65583 10194 65592
rect 10140 65068 10192 65074
rect 10140 65010 10192 65016
rect 10152 64841 10180 65010
rect 10138 64832 10194 64841
rect 10138 64767 10194 64776
rect 10140 64456 10192 64462
rect 10140 64398 10192 64404
rect 10152 64161 10180 64398
rect 10138 64152 10194 64161
rect 10138 64087 10194 64096
rect 10140 62892 10192 62898
rect 10140 62834 10192 62840
rect 10152 62529 10180 62834
rect 10138 62520 10194 62529
rect 10138 62455 10194 62464
rect 10140 62280 10192 62286
rect 10140 62222 10192 62228
rect 10152 61849 10180 62222
rect 10138 61840 10194 61849
rect 10138 61775 10194 61784
rect 10140 61192 10192 61198
rect 10140 61134 10192 61140
rect 10152 61033 10180 61134
rect 10138 61024 10194 61033
rect 10138 60959 10194 60968
rect 10140 60716 10192 60722
rect 10140 60658 10192 60664
rect 10152 60353 10180 60658
rect 10138 60344 10194 60353
rect 10138 60279 10194 60288
rect 10140 59016 10192 59022
rect 10140 58958 10192 58964
rect 9956 58880 10008 58886
rect 9956 58822 10008 58828
rect 9968 56982 9996 58822
rect 10152 58721 10180 58958
rect 10138 58712 10194 58721
rect 10138 58647 10194 58656
rect 10140 58540 10192 58546
rect 10140 58482 10192 58488
rect 10152 58041 10180 58482
rect 10138 58032 10194 58041
rect 10138 57967 10194 57976
rect 9956 56976 10008 56982
rect 9956 56918 10008 56924
rect 9956 56160 10008 56166
rect 9956 56102 10008 56108
rect 9864 54528 9916 54534
rect 9864 54470 9916 54476
rect 9876 54194 9904 54470
rect 9864 54188 9916 54194
rect 9864 54130 9916 54136
rect 9968 53582 9996 56102
rect 10140 55616 10192 55622
rect 10140 55558 10192 55564
rect 10152 54670 10180 55558
rect 10140 54664 10192 54670
rect 10140 54606 10192 54612
rect 10232 54256 10284 54262
rect 10232 54198 10284 54204
rect 10046 54088 10102 54097
rect 10046 54023 10048 54032
rect 10100 54023 10102 54032
rect 10048 53994 10100 54000
rect 9956 53576 10008 53582
rect 9956 53518 10008 53524
rect 10048 53440 10100 53446
rect 10046 53408 10048 53417
rect 10100 53408 10102 53417
rect 10046 53343 10102 53352
rect 10048 52896 10100 52902
rect 10048 52838 10100 52844
rect 10060 52601 10088 52838
rect 10046 52592 10102 52601
rect 10046 52527 10102 52536
rect 10140 52488 10192 52494
rect 10140 52430 10192 52436
rect 9864 52352 9916 52358
rect 9864 52294 9916 52300
rect 9876 52018 9904 52294
rect 10152 52154 10180 52430
rect 10140 52148 10192 52154
rect 10140 52090 10192 52096
rect 9864 52012 9916 52018
rect 9864 51954 9916 51960
rect 10140 51876 10192 51882
rect 10140 51818 10192 51824
rect 10048 51808 10100 51814
rect 10046 51776 10048 51785
rect 10100 51776 10102 51785
rect 10046 51711 10102 51720
rect 9864 51400 9916 51406
rect 9864 51342 9916 51348
rect 9876 51066 9904 51342
rect 10048 51264 10100 51270
rect 10048 51206 10100 51212
rect 10060 51105 10088 51206
rect 10046 51096 10102 51105
rect 9864 51060 9916 51066
rect 10046 51031 10102 51040
rect 9864 51002 9916 51008
rect 10152 50930 10180 51818
rect 10140 50924 10192 50930
rect 10140 50866 10192 50872
rect 9864 50312 9916 50318
rect 9864 50254 9916 50260
rect 10046 50280 10102 50289
rect 9876 48890 9904 50254
rect 10046 50215 10102 50224
rect 10060 50182 10088 50215
rect 10048 50176 10100 50182
rect 10048 50118 10100 50124
rect 9956 49224 10008 49230
rect 9956 49166 10008 49172
rect 9864 48884 9916 48890
rect 9864 48826 9916 48832
rect 9968 47258 9996 49166
rect 10048 49088 10100 49094
rect 10048 49030 10100 49036
rect 10060 48793 10088 49030
rect 10046 48784 10102 48793
rect 10046 48719 10102 48728
rect 10048 48000 10100 48006
rect 10046 47968 10048 47977
rect 10100 47968 10102 47977
rect 10046 47903 10102 47912
rect 10048 47456 10100 47462
rect 10048 47398 10100 47404
rect 9956 47252 10008 47258
rect 9956 47194 10008 47200
rect 10060 47161 10088 47398
rect 10046 47152 10102 47161
rect 10046 47087 10102 47096
rect 10046 46472 10102 46481
rect 10046 46407 10048 46416
rect 10100 46407 10102 46416
rect 10048 46378 10100 46384
rect 10048 45824 10100 45830
rect 10048 45766 10100 45772
rect 10060 45665 10088 45766
rect 10046 45656 10102 45665
rect 10046 45591 10102 45600
rect 9864 44872 9916 44878
rect 9864 44814 9916 44820
rect 10046 44840 10102 44849
rect 9876 44538 9904 44814
rect 10046 44775 10102 44784
rect 10060 44742 10088 44775
rect 10048 44736 10100 44742
rect 10048 44678 10100 44684
rect 9864 44532 9916 44538
rect 9864 44474 9916 44480
rect 9864 44396 9916 44402
rect 9864 44338 9916 44344
rect 9772 43240 9824 43246
rect 9772 43182 9824 43188
rect 9876 42566 9904 44338
rect 10048 44192 10100 44198
rect 10046 44160 10048 44169
rect 10100 44160 10102 44169
rect 10046 44095 10102 44104
rect 9956 43784 10008 43790
rect 9956 43726 10008 43732
rect 9968 43450 9996 43726
rect 10048 43648 10100 43654
rect 10048 43590 10100 43596
rect 9956 43444 10008 43450
rect 9956 43386 10008 43392
rect 10060 43353 10088 43590
rect 10046 43344 10102 43353
rect 10046 43279 10102 43288
rect 9956 42696 10008 42702
rect 9956 42638 10008 42644
rect 9864 42560 9916 42566
rect 9864 42502 9916 42508
rect 9968 41818 9996 42638
rect 10048 42560 10100 42566
rect 10046 42528 10048 42537
rect 10100 42528 10102 42537
rect 10046 42463 10102 42472
rect 10048 42016 10100 42022
rect 10048 41958 10100 41964
rect 10060 41857 10088 41958
rect 10046 41848 10102 41857
rect 9680 41812 9732 41818
rect 9680 41754 9732 41760
rect 9956 41812 10008 41818
rect 10046 41783 10102 41792
rect 9956 41754 10008 41760
rect 10244 41698 10272 54198
rect 9692 41670 10272 41698
rect 9496 40724 9548 40730
rect 9496 40666 9548 40672
rect 9110 39740 9418 39760
rect 9110 39738 9116 39740
rect 9172 39738 9196 39740
rect 9252 39738 9276 39740
rect 9332 39738 9356 39740
rect 9412 39738 9418 39740
rect 9172 39686 9174 39738
rect 9354 39686 9356 39738
rect 9110 39684 9116 39686
rect 9172 39684 9196 39686
rect 9252 39684 9276 39686
rect 9332 39684 9356 39686
rect 9412 39684 9418 39686
rect 9110 39664 9418 39684
rect 8760 39432 8812 39438
rect 8760 39374 8812 39380
rect 8772 33658 8800 39374
rect 9110 38652 9418 38672
rect 9110 38650 9116 38652
rect 9172 38650 9196 38652
rect 9252 38650 9276 38652
rect 9332 38650 9356 38652
rect 9412 38650 9418 38652
rect 9172 38598 9174 38650
rect 9354 38598 9356 38650
rect 9110 38596 9116 38598
rect 9172 38596 9196 38598
rect 9252 38596 9276 38598
rect 9332 38596 9356 38598
rect 9412 38596 9418 38598
rect 9110 38576 9418 38596
rect 9110 37564 9418 37584
rect 9110 37562 9116 37564
rect 9172 37562 9196 37564
rect 9252 37562 9276 37564
rect 9332 37562 9356 37564
rect 9412 37562 9418 37564
rect 9172 37510 9174 37562
rect 9354 37510 9356 37562
rect 9110 37508 9116 37510
rect 9172 37508 9196 37510
rect 9252 37508 9276 37510
rect 9332 37508 9356 37510
rect 9412 37508 9418 37510
rect 9110 37488 9418 37508
rect 9110 36476 9418 36496
rect 9110 36474 9116 36476
rect 9172 36474 9196 36476
rect 9252 36474 9276 36476
rect 9332 36474 9356 36476
rect 9412 36474 9418 36476
rect 9172 36422 9174 36474
rect 9354 36422 9356 36474
rect 9110 36420 9116 36422
rect 9172 36420 9196 36422
rect 9252 36420 9276 36422
rect 9332 36420 9356 36422
rect 9412 36420 9418 36422
rect 9110 36400 9418 36420
rect 9110 35388 9418 35408
rect 9110 35386 9116 35388
rect 9172 35386 9196 35388
rect 9252 35386 9276 35388
rect 9332 35386 9356 35388
rect 9412 35386 9418 35388
rect 9172 35334 9174 35386
rect 9354 35334 9356 35386
rect 9110 35332 9116 35334
rect 9172 35332 9196 35334
rect 9252 35332 9276 35334
rect 9332 35332 9356 35334
rect 9412 35332 9418 35334
rect 9110 35312 9418 35332
rect 9588 34740 9640 34746
rect 9588 34682 9640 34688
rect 9110 34300 9418 34320
rect 9110 34298 9116 34300
rect 9172 34298 9196 34300
rect 9252 34298 9276 34300
rect 9332 34298 9356 34300
rect 9412 34298 9418 34300
rect 9172 34246 9174 34298
rect 9354 34246 9356 34298
rect 9110 34244 9116 34246
rect 9172 34244 9196 34246
rect 9252 34244 9276 34246
rect 9332 34244 9356 34246
rect 9412 34244 9418 34246
rect 9110 34224 9418 34244
rect 9600 34105 9628 34682
rect 9586 34096 9642 34105
rect 9586 34031 9642 34040
rect 8760 33652 8812 33658
rect 8760 33594 8812 33600
rect 9110 33212 9418 33232
rect 9110 33210 9116 33212
rect 9172 33210 9196 33212
rect 9252 33210 9276 33212
rect 9332 33210 9356 33212
rect 9412 33210 9418 33212
rect 9172 33158 9174 33210
rect 9354 33158 9356 33210
rect 9110 33156 9116 33158
rect 9172 33156 9196 33158
rect 9252 33156 9276 33158
rect 9332 33156 9356 33158
rect 9412 33156 9418 33158
rect 9110 33136 9418 33156
rect 9692 32978 9720 41670
rect 9772 41608 9824 41614
rect 9772 41550 9824 41556
rect 9784 38010 9812 41550
rect 10046 41032 10102 41041
rect 10046 40967 10048 40976
rect 10100 40967 10102 40976
rect 10048 40938 10100 40944
rect 9864 40520 9916 40526
rect 9864 40462 9916 40468
rect 9876 40186 9904 40462
rect 10048 40384 10100 40390
rect 10046 40352 10048 40361
rect 10100 40352 10102 40361
rect 10046 40287 10102 40296
rect 9864 40180 9916 40186
rect 9864 40122 9916 40128
rect 9864 40044 9916 40050
rect 9864 39986 9916 39992
rect 9876 39642 9904 39986
rect 10048 39840 10100 39846
rect 10048 39782 10100 39788
rect 9864 39636 9916 39642
rect 9864 39578 9916 39584
rect 10060 39545 10088 39782
rect 10046 39536 10102 39545
rect 10046 39471 10102 39480
rect 10048 38752 10100 38758
rect 10046 38720 10048 38729
rect 10100 38720 10102 38729
rect 10046 38655 10102 38664
rect 10048 38208 10100 38214
rect 10048 38150 10100 38156
rect 10060 38049 10088 38150
rect 10046 38040 10102 38049
rect 9772 38004 9824 38010
rect 10046 37975 10102 37984
rect 9772 37946 9824 37952
rect 10046 37224 10102 37233
rect 10046 37159 10102 37168
rect 10060 37126 10088 37159
rect 10048 37120 10100 37126
rect 10048 37062 10100 37068
rect 9864 36780 9916 36786
rect 9864 36722 9916 36728
rect 9876 36378 9904 36722
rect 10048 36576 10100 36582
rect 10048 36518 10100 36524
rect 10060 36417 10088 36518
rect 10046 36408 10102 36417
rect 9864 36372 9916 36378
rect 10046 36343 10102 36352
rect 9864 36314 9916 36320
rect 9864 36168 9916 36174
rect 9864 36110 9916 36116
rect 9876 35290 9904 36110
rect 10048 36032 10100 36038
rect 10048 35974 10100 35980
rect 10060 35737 10088 35974
rect 10046 35728 10102 35737
rect 10046 35663 10102 35672
rect 9864 35284 9916 35290
rect 9864 35226 9916 35232
rect 10048 34944 10100 34950
rect 10046 34912 10048 34921
rect 10100 34912 10102 34921
rect 10046 34847 10102 34856
rect 9864 33516 9916 33522
rect 9864 33458 9916 33464
rect 9680 32972 9732 32978
rect 9680 32914 9732 32920
rect 9110 32124 9418 32144
rect 9110 32122 9116 32124
rect 9172 32122 9196 32124
rect 9252 32122 9276 32124
rect 9332 32122 9356 32124
rect 9412 32122 9418 32124
rect 9172 32070 9174 32122
rect 9354 32070 9356 32122
rect 9110 32068 9116 32070
rect 9172 32068 9196 32070
rect 9252 32068 9276 32070
rect 9332 32068 9356 32070
rect 9412 32068 9418 32070
rect 9110 32048 9418 32068
rect 9110 31036 9418 31056
rect 9110 31034 9116 31036
rect 9172 31034 9196 31036
rect 9252 31034 9276 31036
rect 9332 31034 9356 31036
rect 9412 31034 9418 31036
rect 9172 30982 9174 31034
rect 9354 30982 9356 31034
rect 9110 30980 9116 30982
rect 9172 30980 9196 30982
rect 9252 30980 9276 30982
rect 9332 30980 9356 30982
rect 9412 30980 9418 30982
rect 9110 30960 9418 30980
rect 8668 30184 8720 30190
rect 8668 30126 8720 30132
rect 9110 29948 9418 29968
rect 9110 29946 9116 29948
rect 9172 29946 9196 29948
rect 9252 29946 9276 29948
rect 9332 29946 9356 29948
rect 9412 29946 9418 29948
rect 9172 29894 9174 29946
rect 9354 29894 9356 29946
rect 9110 29892 9116 29894
rect 9172 29892 9196 29894
rect 9252 29892 9276 29894
rect 9332 29892 9356 29894
rect 9412 29892 9418 29894
rect 9110 29872 9418 29892
rect 9110 28860 9418 28880
rect 9110 28858 9116 28860
rect 9172 28858 9196 28860
rect 9252 28858 9276 28860
rect 9332 28858 9356 28860
rect 9412 28858 9418 28860
rect 9172 28806 9174 28858
rect 9354 28806 9356 28858
rect 9110 28804 9116 28806
rect 9172 28804 9196 28806
rect 9252 28804 9276 28806
rect 9332 28804 9356 28806
rect 9412 28804 9418 28806
rect 9110 28784 9418 28804
rect 9876 28762 9904 33458
rect 10046 33416 10102 33425
rect 10046 33351 10048 33360
rect 10100 33351 10102 33360
rect 10048 33322 10100 33328
rect 10048 32768 10100 32774
rect 10048 32710 10100 32716
rect 10060 32609 10088 32710
rect 10046 32600 10102 32609
rect 10046 32535 10102 32544
rect 10048 31952 10100 31958
rect 10048 31894 10100 31900
rect 10060 31793 10088 31894
rect 10046 31784 10102 31793
rect 10046 31719 10102 31728
rect 10048 31136 10100 31142
rect 10046 31104 10048 31113
rect 10100 31104 10102 31113
rect 10046 31039 10102 31048
rect 10048 30592 10100 30598
rect 10048 30534 10100 30540
rect 10060 30297 10088 30534
rect 10046 30288 10102 30297
rect 10046 30223 10102 30232
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 10152 29481 10180 29582
rect 10138 29472 10194 29481
rect 10138 29407 10194 29416
rect 10140 29028 10192 29034
rect 10140 28970 10192 28976
rect 10152 28801 10180 28970
rect 10138 28792 10194 28801
rect 9864 28756 9916 28762
rect 10138 28727 10194 28736
rect 9864 28698 9916 28704
rect 9956 28008 10008 28014
rect 9954 27976 9956 27985
rect 10008 27976 10010 27985
rect 9954 27911 10010 27920
rect 9110 27772 9418 27792
rect 9110 27770 9116 27772
rect 9172 27770 9196 27772
rect 9252 27770 9276 27772
rect 9332 27770 9356 27772
rect 9412 27770 9418 27772
rect 9172 27718 9174 27770
rect 9354 27718 9356 27770
rect 9110 27716 9116 27718
rect 9172 27716 9196 27718
rect 9252 27716 9276 27718
rect 9332 27716 9356 27718
rect 9412 27716 9418 27718
rect 9110 27696 9418 27716
rect 9956 27328 10008 27334
rect 9956 27270 10008 27276
rect 9968 27169 9996 27270
rect 9954 27160 10010 27169
rect 9954 27095 10010 27104
rect 10140 26784 10192 26790
rect 10140 26726 10192 26732
rect 9110 26684 9418 26704
rect 9110 26682 9116 26684
rect 9172 26682 9196 26684
rect 9252 26682 9276 26684
rect 9332 26682 9356 26684
rect 9412 26682 9418 26684
rect 9172 26630 9174 26682
rect 9354 26630 9356 26682
rect 9110 26628 9116 26630
rect 9172 26628 9196 26630
rect 9252 26628 9276 26630
rect 9332 26628 9356 26630
rect 9412 26628 9418 26630
rect 9110 26608 9418 26628
rect 10152 26489 10180 26726
rect 10138 26480 10194 26489
rect 10138 26415 10194 26424
rect 10140 25696 10192 25702
rect 10138 25664 10140 25673
rect 10192 25664 10194 25673
rect 9110 25596 9418 25616
rect 10138 25599 10194 25608
rect 9110 25594 9116 25596
rect 9172 25594 9196 25596
rect 9252 25594 9276 25596
rect 9332 25594 9356 25596
rect 9412 25594 9418 25596
rect 9172 25542 9174 25594
rect 9354 25542 9356 25594
rect 9110 25540 9116 25542
rect 9172 25540 9196 25542
rect 9252 25540 9276 25542
rect 9332 25540 9356 25542
rect 9412 25540 9418 25542
rect 9110 25520 9418 25540
rect 10140 25288 10192 25294
rect 10140 25230 10192 25236
rect 10152 24857 10180 25230
rect 10138 24848 10194 24857
rect 10138 24783 10194 24792
rect 9110 24508 9418 24528
rect 9110 24506 9116 24508
rect 9172 24506 9196 24508
rect 9252 24506 9276 24508
rect 9332 24506 9356 24508
rect 9412 24506 9418 24508
rect 9172 24454 9174 24506
rect 9354 24454 9356 24506
rect 9110 24452 9116 24454
rect 9172 24452 9196 24454
rect 9252 24452 9276 24454
rect 9332 24452 9356 24454
rect 9412 24452 9418 24454
rect 9110 24432 9418 24452
rect 10140 24200 10192 24206
rect 10138 24168 10140 24177
rect 10192 24168 10194 24177
rect 10138 24103 10194 24112
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 9110 23420 9418 23440
rect 9110 23418 9116 23420
rect 9172 23418 9196 23420
rect 9252 23418 9276 23420
rect 9332 23418 9356 23420
rect 9412 23418 9418 23420
rect 9172 23366 9174 23418
rect 9354 23366 9356 23418
rect 9110 23364 9116 23366
rect 9172 23364 9196 23366
rect 9252 23364 9276 23366
rect 9332 23364 9356 23366
rect 9412 23364 9418 23366
rect 9110 23344 9418 23364
rect 10152 23361 10180 23462
rect 10138 23352 10194 23361
rect 10138 23287 10194 23296
rect 10138 22536 10194 22545
rect 10138 22471 10140 22480
rect 10192 22471 10194 22480
rect 10140 22442 10192 22448
rect 9110 22332 9418 22352
rect 9110 22330 9116 22332
rect 9172 22330 9196 22332
rect 9252 22330 9276 22332
rect 9332 22330 9356 22332
rect 9412 22330 9418 22332
rect 9172 22278 9174 22330
rect 9354 22278 9356 22330
rect 9110 22276 9116 22278
rect 9172 22276 9196 22278
rect 9252 22276 9276 22278
rect 9332 22276 9356 22278
rect 9412 22276 9418 22278
rect 9110 22256 9418 22276
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 10152 21865 10180 22102
rect 10138 21856 10194 21865
rect 10138 21791 10194 21800
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 9110 21244 9418 21264
rect 9110 21242 9116 21244
rect 9172 21242 9196 21244
rect 9252 21242 9276 21244
rect 9332 21242 9356 21244
rect 9412 21242 9418 21244
rect 9172 21190 9174 21242
rect 9354 21190 9356 21242
rect 9110 21188 9116 21190
rect 9172 21188 9196 21190
rect 9252 21188 9276 21190
rect 9332 21188 9356 21190
rect 9412 21188 9418 21190
rect 9110 21168 9418 21188
rect 10152 21049 10180 21286
rect 10138 21040 10194 21049
rect 10138 20975 10194 20984
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10046 20360 10102 20369
rect 10046 20295 10048 20304
rect 10100 20295 10102 20304
rect 10048 20266 10100 20272
rect 9110 20156 9418 20176
rect 9110 20154 9116 20156
rect 9172 20154 9196 20156
rect 9252 20154 9276 20156
rect 9332 20154 9356 20156
rect 9412 20154 9418 20156
rect 9172 20102 9174 20154
rect 9354 20102 9356 20154
rect 9110 20100 9116 20102
rect 9172 20100 9196 20102
rect 9252 20100 9276 20102
rect 9332 20100 9356 20102
rect 9412 20100 9418 20102
rect 9110 20080 9418 20100
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9232 19514 9260 19790
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10060 19553 10088 19654
rect 10046 19544 10102 19553
rect 9220 19508 9272 19514
rect 10046 19479 10102 19488
rect 9220 19450 9272 19456
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9110 19068 9418 19088
rect 9110 19066 9116 19068
rect 9172 19066 9196 19068
rect 9252 19066 9276 19068
rect 9332 19066 9356 19068
rect 9412 19066 9418 19068
rect 9172 19014 9174 19066
rect 9354 19014 9356 19066
rect 9110 19012 9116 19014
rect 9172 19012 9196 19014
rect 9252 19012 9276 19014
rect 9332 19012 9356 19014
rect 9412 19012 9418 19014
rect 9110 18992 9418 19012
rect 9876 18766 9904 19110
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 10046 18728 10102 18737
rect 10046 18663 10102 18672
rect 10060 18630 10088 18663
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9110 17980 9418 18000
rect 9110 17978 9116 17980
rect 9172 17978 9196 17980
rect 9252 17978 9276 17980
rect 9332 17978 9356 17980
rect 9412 17978 9418 17980
rect 9172 17926 9174 17978
rect 9354 17926 9356 17978
rect 9110 17924 9116 17926
rect 9172 17924 9196 17926
rect 9252 17924 9276 17926
rect 9332 17924 9356 17926
rect 9412 17924 9418 17926
rect 9110 17904 9418 17924
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 9048 13530 9076 17614
rect 9876 17338 9904 18226
rect 10048 18080 10100 18086
rect 10046 18048 10048 18057
rect 10100 18048 10102 18057
rect 10046 17983 10102 17992
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 10060 17241 10088 17478
rect 10046 17232 10102 17241
rect 10046 17167 10102 17176
rect 9110 16892 9418 16912
rect 9110 16890 9116 16892
rect 9172 16890 9196 16892
rect 9252 16890 9276 16892
rect 9332 16890 9356 16892
rect 9412 16890 9418 16892
rect 9172 16838 9174 16890
rect 9354 16838 9356 16890
rect 9110 16836 9116 16838
rect 9172 16836 9196 16838
rect 9252 16836 9276 16838
rect 9332 16836 9356 16838
rect 9412 16836 9418 16838
rect 9110 16816 9418 16836
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 9232 16250 9260 16526
rect 10048 16448 10100 16454
rect 10046 16416 10048 16425
rect 10100 16416 10102 16425
rect 10046 16351 10102 16360
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9110 15804 9418 15824
rect 9110 15802 9116 15804
rect 9172 15802 9196 15804
rect 9252 15802 9276 15804
rect 9332 15802 9356 15804
rect 9412 15802 9418 15804
rect 9172 15750 9174 15802
rect 9354 15750 9356 15802
rect 9110 15748 9116 15750
rect 9172 15748 9196 15750
rect 9252 15748 9276 15750
rect 9332 15748 9356 15750
rect 9412 15748 9418 15750
rect 9110 15728 9418 15748
rect 9968 15706 9996 16050
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10060 15745 10088 15846
rect 10046 15736 10102 15745
rect 9956 15700 10008 15706
rect 10046 15671 10102 15680
rect 9956 15642 10008 15648
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9110 14716 9418 14736
rect 9110 14714 9116 14716
rect 9172 14714 9196 14716
rect 9252 14714 9276 14716
rect 9332 14714 9356 14716
rect 9412 14714 9418 14716
rect 9172 14662 9174 14714
rect 9354 14662 9356 14714
rect 9110 14660 9116 14662
rect 9172 14660 9196 14662
rect 9252 14660 9276 14662
rect 9332 14660 9356 14662
rect 9412 14660 9418 14662
rect 9110 14640 9418 14660
rect 9508 14074 9536 14962
rect 10046 14920 10102 14929
rect 10046 14855 10048 14864
rect 10100 14855 10102 14864
rect 10048 14826 10100 14832
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9110 13628 9418 13648
rect 9110 13626 9116 13628
rect 9172 13626 9196 13628
rect 9252 13626 9276 13628
rect 9332 13626 9356 13628
rect 9412 13626 9418 13628
rect 9172 13574 9174 13626
rect 9354 13574 9356 13626
rect 9110 13572 9116 13574
rect 9172 13572 9196 13574
rect 9252 13572 9276 13574
rect 9332 13572 9356 13574
rect 9412 13572 9418 13574
rect 9110 13552 9418 13572
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9600 13433 9628 14010
rect 9876 13530 9904 14350
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 14113 10088 14214
rect 10046 14104 10102 14113
rect 10046 14039 10102 14048
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9586 13424 9642 13433
rect 9586 13359 9642 13368
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9508 12782 9536 13262
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 10048 12640 10100 12646
rect 10046 12608 10048 12617
rect 10100 12608 10102 12617
rect 9110 12540 9418 12560
rect 10046 12543 10102 12552
rect 9110 12538 9116 12540
rect 9172 12538 9196 12540
rect 9252 12538 9276 12540
rect 9332 12538 9356 12540
rect 9412 12538 9418 12540
rect 9172 12486 9174 12538
rect 9354 12486 9356 12538
rect 9110 12484 9116 12486
rect 9172 12484 9196 12486
rect 9252 12484 9276 12486
rect 9332 12484 9356 12486
rect 9412 12484 9418 12486
rect 9110 12464 9418 12484
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10060 11801 10088 12038
rect 10152 11898 10180 20402
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10046 11792 10102 11801
rect 10046 11727 10102 11736
rect 9110 11452 9418 11472
rect 9110 11450 9116 11452
rect 9172 11450 9196 11452
rect 9252 11450 9276 11452
rect 9332 11450 9356 11452
rect 9412 11450 9418 11452
rect 9172 11398 9174 11450
rect 9354 11398 9356 11450
rect 9110 11396 9116 11398
rect 9172 11396 9196 11398
rect 9252 11396 9276 11398
rect 9332 11396 9356 11398
rect 9412 11396 9418 11398
rect 9110 11376 9418 11396
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9864 11144 9916 11150
rect 10060 11121 10088 11222
rect 9864 11086 9916 11092
rect 10046 11112 10102 11121
rect 9876 10810 9904 11086
rect 10046 11047 10102 11056
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9110 10364 9418 10384
rect 9110 10362 9116 10364
rect 9172 10362 9196 10364
rect 9252 10362 9276 10364
rect 9332 10362 9356 10364
rect 9412 10362 9418 10364
rect 9172 10310 9174 10362
rect 9354 10310 9356 10362
rect 9110 10308 9116 10310
rect 9172 10308 9196 10310
rect 9252 10308 9276 10310
rect 9332 10308 9356 10310
rect 9412 10308 9418 10310
rect 9110 10288 9418 10308
rect 9876 9450 9904 10610
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 10305 10088 10406
rect 10046 10296 10102 10305
rect 10046 10231 10102 10240
rect 10046 9480 10102 9489
rect 9864 9444 9916 9450
rect 10046 9415 10048 9424
rect 9864 9386 9916 9392
rect 10100 9415 10102 9424
rect 10048 9386 10100 9392
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 5846 9276 6154 9296
rect 5846 9274 5852 9276
rect 5908 9274 5932 9276
rect 5988 9274 6012 9276
rect 6068 9274 6092 9276
rect 6148 9274 6154 9276
rect 5908 9222 5910 9274
rect 6090 9222 6092 9274
rect 5846 9220 5852 9222
rect 5908 9220 5932 9222
rect 5988 9220 6012 9222
rect 6068 9220 6092 9222
rect 6148 9220 6154 9222
rect 5846 9200 6154 9220
rect 9110 9276 9418 9296
rect 9110 9274 9116 9276
rect 9172 9274 9196 9276
rect 9252 9274 9276 9276
rect 9332 9274 9356 9276
rect 9412 9274 9418 9276
rect 9172 9222 9174 9274
rect 9354 9222 9356 9274
rect 9110 9220 9116 9222
rect 9172 9220 9196 9222
rect 9252 9220 9276 9222
rect 9332 9220 9356 9222
rect 9412 9220 9418 9222
rect 9110 9200 9418 9220
rect 10048 8832 10100 8838
rect 10046 8800 10048 8809
rect 10100 8800 10102 8809
rect 7478 8732 7786 8752
rect 10046 8735 10102 8744
rect 7478 8730 7484 8732
rect 7540 8730 7564 8732
rect 7620 8730 7644 8732
rect 7700 8730 7724 8732
rect 7780 8730 7786 8732
rect 7540 8678 7542 8730
rect 7722 8678 7724 8730
rect 7478 8676 7484 8678
rect 7540 8676 7564 8678
rect 7620 8676 7644 8678
rect 7700 8676 7724 8678
rect 7780 8676 7786 8678
rect 7478 8656 7786 8676
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 5846 8188 6154 8208
rect 5846 8186 5852 8188
rect 5908 8186 5932 8188
rect 5988 8186 6012 8188
rect 6068 8186 6092 8188
rect 6148 8186 6154 8188
rect 5908 8134 5910 8186
rect 6090 8134 6092 8186
rect 5846 8132 5852 8134
rect 5908 8132 5932 8134
rect 5988 8132 6012 8134
rect 6068 8132 6092 8134
rect 6148 8132 6154 8134
rect 5846 8112 6154 8132
rect 9110 8188 9418 8208
rect 9110 8186 9116 8188
rect 9172 8186 9196 8188
rect 9252 8186 9276 8188
rect 9332 8186 9356 8188
rect 9412 8186 9418 8188
rect 9172 8134 9174 8186
rect 9354 8134 9356 8186
rect 9110 8132 9116 8134
rect 9172 8132 9196 8134
rect 9252 8132 9276 8134
rect 9332 8132 9356 8134
rect 9412 8132 9418 8134
rect 9110 8112 9418 8132
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 10060 7993 10088 8298
rect 10046 7984 10102 7993
rect 10046 7919 10102 7928
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 7478 7644 7786 7664
rect 7478 7642 7484 7644
rect 7540 7642 7564 7644
rect 7620 7642 7644 7644
rect 7700 7642 7724 7644
rect 7780 7642 7786 7644
rect 7540 7590 7542 7642
rect 7722 7590 7724 7642
rect 7478 7588 7484 7590
rect 7540 7588 7564 7590
rect 7620 7588 7644 7590
rect 7700 7588 7724 7590
rect 7780 7588 7786 7590
rect 7478 7568 7786 7588
rect 9876 7410 9904 7686
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9864 7200 9916 7206
rect 10048 7200 10100 7206
rect 9864 7142 9916 7148
rect 10046 7168 10048 7177
rect 10100 7168 10102 7177
rect 5846 7100 6154 7120
rect 5846 7098 5852 7100
rect 5908 7098 5932 7100
rect 5988 7098 6012 7100
rect 6068 7098 6092 7100
rect 6148 7098 6154 7100
rect 5908 7046 5910 7098
rect 6090 7046 6092 7098
rect 5846 7044 5852 7046
rect 5908 7044 5932 7046
rect 5988 7044 6012 7046
rect 6068 7044 6092 7046
rect 6148 7044 6154 7046
rect 5846 7024 6154 7044
rect 9110 7100 9418 7120
rect 9110 7098 9116 7100
rect 9172 7098 9196 7100
rect 9252 7098 9276 7100
rect 9332 7098 9356 7100
rect 9412 7098 9418 7100
rect 9172 7046 9174 7098
rect 9354 7046 9356 7098
rect 9110 7044 9116 7046
rect 9172 7044 9196 7046
rect 9252 7044 9276 7046
rect 9332 7044 9356 7046
rect 9412 7044 9418 7046
rect 9110 7024 9418 7044
rect 9876 6798 9904 7142
rect 10046 7103 10102 7112
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 7478 6556 7786 6576
rect 7478 6554 7484 6556
rect 7540 6554 7564 6556
rect 7620 6554 7644 6556
rect 7700 6554 7724 6556
rect 7780 6554 7786 6556
rect 7540 6502 7542 6554
rect 7722 6502 7724 6554
rect 7478 6500 7484 6502
rect 7540 6500 7564 6502
rect 7620 6500 7644 6502
rect 7700 6500 7724 6502
rect 7780 6500 7786 6502
rect 7478 6480 7786 6500
rect 10060 6497 10088 6598
rect 10046 6488 10102 6497
rect 10046 6423 10102 6432
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 5846 6012 6154 6032
rect 5846 6010 5852 6012
rect 5908 6010 5932 6012
rect 5988 6010 6012 6012
rect 6068 6010 6092 6012
rect 6148 6010 6154 6012
rect 5908 5958 5910 6010
rect 6090 5958 6092 6010
rect 5846 5956 5852 5958
rect 5908 5956 5932 5958
rect 5988 5956 6012 5958
rect 6068 5956 6092 5958
rect 6148 5956 6154 5958
rect 5846 5936 6154 5956
rect 7478 5468 7786 5488
rect 7478 5466 7484 5468
rect 7540 5466 7564 5468
rect 7620 5466 7644 5468
rect 7700 5466 7724 5468
rect 7780 5466 7786 5468
rect 7540 5414 7542 5466
rect 7722 5414 7724 5466
rect 7478 5412 7484 5414
rect 7540 5412 7564 5414
rect 7620 5412 7644 5414
rect 7700 5412 7724 5414
rect 7780 5412 7786 5414
rect 7478 5392 7786 5412
rect 9048 5234 9076 6054
rect 9110 6012 9418 6032
rect 9110 6010 9116 6012
rect 9172 6010 9196 6012
rect 9252 6010 9276 6012
rect 9332 6010 9356 6012
rect 9412 6010 9418 6012
rect 9172 5958 9174 6010
rect 9354 5958 9356 6010
rect 9110 5956 9116 5958
rect 9172 5956 9196 5958
rect 9252 5956 9276 5958
rect 9332 5956 9356 5958
rect 9412 5956 9418 5958
rect 9110 5936 9418 5956
rect 10046 5672 10102 5681
rect 10046 5607 10102 5616
rect 10060 5574 10088 5607
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 5846 4924 6154 4944
rect 5846 4922 5852 4924
rect 5908 4922 5932 4924
rect 5988 4922 6012 4924
rect 6068 4922 6092 4924
rect 6148 4922 6154 4924
rect 5908 4870 5910 4922
rect 6090 4870 6092 4922
rect 5846 4868 5852 4870
rect 5908 4868 5932 4870
rect 5988 4868 6012 4870
rect 6068 4868 6092 4870
rect 6148 4868 6154 4870
rect 5846 4848 6154 4868
rect 9110 4924 9418 4944
rect 9110 4922 9116 4924
rect 9172 4922 9196 4924
rect 9252 4922 9276 4924
rect 9332 4922 9356 4924
rect 9412 4922 9418 4924
rect 9172 4870 9174 4922
rect 9354 4870 9356 4922
rect 9110 4868 9116 4870
rect 9172 4868 9196 4870
rect 9252 4868 9276 4870
rect 9332 4868 9356 4870
rect 9412 4868 9418 4870
rect 9110 4848 9418 4868
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4066 4720 4122 4729
rect 4066 4655 4122 4664
rect 9876 4622 9904 4966
rect 10060 4865 10088 4966
rect 10046 4856 10102 4865
rect 10046 4791 10102 4800
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 4160 4548 4212 4554
rect 4080 4508 4160 4536
rect 4080 4162 4108 4508
rect 4160 4490 4212 4496
rect 4214 4380 4522 4400
rect 4214 4378 4220 4380
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4516 4378 4522 4380
rect 4276 4326 4278 4378
rect 4458 4326 4460 4378
rect 4214 4324 4220 4326
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4516 4324 4522 4326
rect 4214 4304 4522 4324
rect 4816 4282 4844 4558
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 7478 4380 7786 4400
rect 7478 4378 7484 4380
rect 7540 4378 7564 4380
rect 7620 4378 7644 4380
rect 7700 4378 7724 4380
rect 7780 4378 7786 4380
rect 7540 4326 7542 4378
rect 7722 4326 7724 4378
rect 7478 4324 7484 4326
rect 7540 4324 7564 4326
rect 7620 4324 7644 4326
rect 7700 4324 7724 4326
rect 7780 4324 7786 4326
rect 7478 4304 7786 4324
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4080 4134 4200 4162
rect 4172 3534 4200 4134
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4632 3534 4660 3878
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4214 3292 4522 3312
rect 4214 3290 4220 3292
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4516 3290 4522 3292
rect 4276 3238 4278 3290
rect 4458 3238 4460 3290
rect 4214 3236 4220 3238
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4516 3236 4522 3238
rect 4214 3216 4522 3236
rect 5092 3058 5120 3878
rect 5846 3836 6154 3856
rect 5846 3834 5852 3836
rect 5908 3834 5932 3836
rect 5988 3834 6012 3836
rect 6068 3834 6092 3836
rect 6148 3834 6154 3836
rect 5908 3782 5910 3834
rect 6090 3782 6092 3834
rect 5846 3780 5852 3782
rect 5908 3780 5932 3782
rect 5988 3780 6012 3782
rect 6068 3780 6092 3782
rect 6148 3780 6154 3782
rect 5846 3760 6154 3780
rect 9110 3836 9418 3856
rect 9110 3834 9116 3836
rect 9172 3834 9196 3836
rect 9252 3834 9276 3836
rect 9332 3834 9356 3836
rect 9412 3834 9418 3836
rect 9172 3782 9174 3834
rect 9354 3782 9356 3834
rect 9110 3780 9116 3782
rect 9172 3780 9196 3782
rect 9252 3780 9276 3782
rect 9332 3780 9356 3782
rect 9412 3780 9418 3782
rect 9110 3760 9418 3780
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 3976 2576 4028 2582
rect 3514 2544 3570 2553
rect 3976 2518 4028 2524
rect 3514 2479 3570 2488
rect 5552 2446 5580 3606
rect 9876 3534 9904 4422
rect 10060 4185 10088 4422
rect 10046 4176 10102 4185
rect 10046 4111 10102 4120
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 7478 3292 7786 3312
rect 7478 3290 7484 3292
rect 7540 3290 7564 3292
rect 7620 3290 7644 3292
rect 7700 3290 7724 3292
rect 7780 3290 7786 3292
rect 7540 3238 7542 3290
rect 7722 3238 7724 3290
rect 7478 3236 7484 3238
rect 7540 3236 7564 3238
rect 7620 3236 7644 3238
rect 7700 3236 7724 3238
rect 7780 3236 7786 3238
rect 7478 3216 7786 3236
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 5846 2748 6154 2768
rect 5846 2746 5852 2748
rect 5908 2746 5932 2748
rect 5988 2746 6012 2748
rect 6068 2746 6092 2748
rect 6148 2746 6154 2748
rect 5908 2694 5910 2746
rect 6090 2694 6092 2746
rect 5846 2692 5852 2694
rect 5908 2692 5932 2694
rect 5988 2692 6012 2694
rect 6068 2692 6092 2694
rect 6148 2692 6154 2694
rect 5846 2672 6154 2692
rect 9110 2748 9418 2768
rect 9110 2746 9116 2748
rect 9172 2746 9196 2748
rect 9252 2746 9276 2748
rect 9332 2746 9356 2748
rect 9412 2746 9418 2748
rect 9172 2694 9174 2746
rect 9354 2694 9356 2746
rect 9110 2692 9116 2694
rect 9172 2692 9196 2694
rect 9252 2692 9276 2694
rect 9332 2692 9356 2694
rect 9412 2692 9418 2694
rect 9110 2672 9418 2692
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 2962 2272 3018 2281
rect 2962 2207 3018 2216
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 2872 1080 2924 1086
rect 2870 1048 2872 1057
rect 2924 1048 2926 1057
rect 2870 983 2926 992
rect 2778 640 2834 649
rect 2778 575 2834 584
rect 3988 241 4016 2382
rect 4214 2204 4522 2224
rect 4214 2202 4220 2204
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4516 2202 4522 2204
rect 4276 2150 4278 2202
rect 4458 2150 4460 2202
rect 4214 2148 4220 2150
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4516 2148 4522 2150
rect 4214 2128 4522 2148
rect 4632 1086 4660 2382
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 7478 2204 7786 2224
rect 7478 2202 7484 2204
rect 7540 2202 7564 2204
rect 7620 2202 7644 2204
rect 7700 2202 7724 2204
rect 7780 2202 7786 2204
rect 7540 2150 7542 2202
rect 7722 2150 7724 2202
rect 7478 2148 7484 2150
rect 7540 2148 7564 2150
rect 7620 2148 7644 2150
rect 7700 2148 7724 2150
rect 7780 2148 7786 2150
rect 7478 2128 7786 2148
rect 4620 1080 4672 1086
rect 4620 1022 4672 1028
rect 9324 377 9352 2246
rect 9508 1873 9536 2790
rect 9692 2446 9720 3402
rect 9864 3392 9916 3398
rect 10048 3392 10100 3398
rect 9864 3334 9916 3340
rect 10046 3360 10048 3369
rect 10100 3360 10102 3369
rect 9876 3058 9904 3334
rect 10046 3295 10102 3304
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10060 2553 10088 2790
rect 10046 2544 10102 2553
rect 10046 2479 10102 2488
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9494 1864 9550 1873
rect 9494 1799 9550 1808
rect 9600 1057 9628 2246
rect 9586 1048 9642 1057
rect 9586 983 9642 992
rect 9310 368 9366 377
rect 9310 303 9366 312
rect 3974 232 4030 241
rect 3974 167 4030 176
<< via2 >>
rect 1398 79192 1454 79248
rect 9954 79464 10010 79520
rect 1306 78784 1362 78840
rect 9586 78648 9642 78704
rect 3882 78376 3938 78432
rect 2588 77818 2644 77820
rect 2668 77818 2724 77820
rect 2748 77818 2804 77820
rect 2828 77818 2884 77820
rect 2588 77766 2634 77818
rect 2634 77766 2644 77818
rect 2668 77766 2698 77818
rect 2698 77766 2710 77818
rect 2710 77766 2724 77818
rect 2748 77766 2762 77818
rect 2762 77766 2774 77818
rect 2774 77766 2804 77818
rect 2828 77766 2838 77818
rect 2838 77766 2884 77818
rect 2588 77764 2644 77766
rect 2668 77764 2724 77766
rect 2748 77764 2804 77766
rect 2828 77764 2884 77766
rect 3606 77560 3662 77616
rect 1490 75792 1546 75848
rect 1582 74568 1638 74624
rect 1582 72800 1638 72856
rect 1398 71576 1454 71632
rect 938 70352 994 70408
rect 1582 72120 1638 72176
rect 1582 71168 1638 71224
rect 478 59880 534 59936
rect 18 45770 74 45826
rect 110 39888 166 39944
rect 662 56888 718 56944
rect 846 56092 902 56094
rect 846 56040 848 56092
rect 848 56040 900 56092
rect 900 56040 902 56092
rect 846 56038 902 56040
rect 1490 70352 1546 70408
rect 1398 69944 1454 70000
rect 2870 76880 2926 76936
rect 1950 74704 2006 74760
rect 1858 70624 1914 70680
rect 1766 70080 1822 70136
rect 1582 69844 1584 69864
rect 1584 69844 1636 69864
rect 1636 69844 1638 69864
rect 1582 69808 1638 69844
rect 1674 69400 1730 69456
rect 1582 68176 1638 68232
rect 1582 67360 1638 67416
rect 1398 66952 1454 67008
rect 1398 66408 1454 66464
rect 1306 66000 1362 66056
rect 1398 65592 1454 65648
rect 1398 65048 1454 65104
rect 1674 66272 1730 66328
rect 1582 65048 1638 65104
rect 1674 64912 1730 64968
rect 1582 63552 1638 63608
rect 1674 62600 1730 62656
rect 1950 70216 2006 70272
rect 1582 61376 1638 61432
rect 1582 60152 1638 60208
rect 1582 59200 1638 59256
rect 1398 57976 1454 58032
rect 1214 56752 1270 56808
rect 1030 46824 1086 46880
rect 662 39888 718 39944
rect 1030 37884 1032 37904
rect 1032 37884 1084 37904
rect 1084 37884 1086 37904
rect 1030 37848 1086 37884
rect 938 28736 994 28792
rect 1582 57568 1638 57624
rect 1582 57432 1638 57488
rect 2226 73208 2282 73264
rect 2588 76730 2644 76732
rect 2668 76730 2724 76732
rect 2748 76730 2804 76732
rect 2828 76730 2884 76732
rect 2588 76678 2634 76730
rect 2634 76678 2644 76730
rect 2668 76678 2698 76730
rect 2698 76678 2710 76730
rect 2710 76678 2724 76730
rect 2748 76678 2762 76730
rect 2762 76678 2774 76730
rect 2774 76678 2804 76730
rect 2828 76678 2838 76730
rect 2838 76678 2884 76730
rect 2588 76676 2644 76678
rect 2668 76676 2724 76678
rect 2748 76676 2804 76678
rect 2828 76676 2884 76678
rect 2962 76200 3018 76256
rect 2588 75642 2644 75644
rect 2668 75642 2724 75644
rect 2748 75642 2804 75644
rect 2828 75642 2884 75644
rect 2588 75590 2634 75642
rect 2634 75590 2644 75642
rect 2668 75590 2698 75642
rect 2698 75590 2710 75642
rect 2710 75590 2724 75642
rect 2748 75590 2762 75642
rect 2762 75590 2774 75642
rect 2774 75590 2804 75642
rect 2828 75590 2838 75642
rect 2838 75590 2884 75642
rect 2588 75588 2644 75590
rect 2668 75588 2724 75590
rect 2748 75588 2804 75590
rect 2828 75588 2884 75590
rect 2226 71984 2282 72040
rect 2226 70760 2282 70816
rect 2318 70216 2374 70272
rect 2226 68992 2282 69048
rect 2588 74554 2644 74556
rect 2668 74554 2724 74556
rect 2748 74554 2804 74556
rect 2828 74554 2884 74556
rect 2588 74502 2634 74554
rect 2634 74502 2644 74554
rect 2668 74502 2698 74554
rect 2698 74502 2710 74554
rect 2710 74502 2724 74554
rect 2748 74502 2762 74554
rect 2762 74502 2774 74554
rect 2774 74502 2804 74554
rect 2828 74502 2838 74554
rect 2838 74502 2884 74554
rect 2588 74500 2644 74502
rect 2668 74500 2724 74502
rect 2748 74500 2804 74502
rect 2828 74500 2884 74502
rect 4066 77968 4122 78024
rect 9494 77968 9550 78024
rect 5852 77818 5908 77820
rect 5932 77818 5988 77820
rect 6012 77818 6068 77820
rect 6092 77818 6148 77820
rect 5852 77766 5898 77818
rect 5898 77766 5908 77818
rect 5932 77766 5962 77818
rect 5962 77766 5974 77818
rect 5974 77766 5988 77818
rect 6012 77766 6026 77818
rect 6026 77766 6038 77818
rect 6038 77766 6068 77818
rect 6092 77766 6102 77818
rect 6102 77766 6148 77818
rect 5852 77764 5908 77766
rect 5932 77764 5988 77766
rect 6012 77764 6068 77766
rect 6092 77764 6148 77766
rect 9116 77818 9172 77820
rect 9196 77818 9252 77820
rect 9276 77818 9332 77820
rect 9356 77818 9412 77820
rect 9116 77766 9162 77818
rect 9162 77766 9172 77818
rect 9196 77766 9226 77818
rect 9226 77766 9238 77818
rect 9238 77766 9252 77818
rect 9276 77766 9290 77818
rect 9290 77766 9302 77818
rect 9302 77766 9332 77818
rect 9356 77766 9366 77818
rect 9366 77766 9412 77818
rect 9116 77764 9172 77766
rect 9196 77764 9252 77766
rect 9276 77764 9332 77766
rect 9356 77764 9412 77766
rect 3974 77152 4030 77208
rect 4220 77274 4276 77276
rect 4300 77274 4356 77276
rect 4380 77274 4436 77276
rect 4460 77274 4516 77276
rect 4220 77222 4266 77274
rect 4266 77222 4276 77274
rect 4300 77222 4330 77274
rect 4330 77222 4342 77274
rect 4342 77222 4356 77274
rect 4380 77222 4394 77274
rect 4394 77222 4406 77274
rect 4406 77222 4436 77274
rect 4460 77222 4470 77274
rect 4470 77222 4516 77274
rect 4220 77220 4276 77222
rect 4300 77220 4356 77222
rect 4380 77220 4436 77222
rect 4460 77220 4516 77222
rect 7484 77274 7540 77276
rect 7564 77274 7620 77276
rect 7644 77274 7700 77276
rect 7724 77274 7780 77276
rect 7484 77222 7530 77274
rect 7530 77222 7540 77274
rect 7564 77222 7594 77274
rect 7594 77222 7606 77274
rect 7606 77222 7620 77274
rect 7644 77222 7658 77274
rect 7658 77222 7670 77274
rect 7670 77222 7700 77274
rect 7724 77222 7734 77274
rect 7734 77222 7780 77274
rect 7484 77220 7540 77222
rect 7564 77220 7620 77222
rect 7644 77220 7700 77222
rect 7724 77220 7780 77222
rect 3238 74976 3294 75032
rect 3238 74196 3240 74216
rect 3240 74196 3292 74216
rect 3292 74196 3294 74216
rect 3238 74160 3294 74196
rect 2962 73752 3018 73808
rect 2588 73466 2644 73468
rect 2668 73466 2724 73468
rect 2748 73466 2804 73468
rect 2828 73466 2884 73468
rect 2588 73414 2634 73466
rect 2634 73414 2644 73466
rect 2668 73414 2698 73466
rect 2698 73414 2710 73466
rect 2710 73414 2724 73466
rect 2748 73414 2762 73466
rect 2762 73414 2774 73466
rect 2774 73414 2804 73466
rect 2828 73414 2838 73466
rect 2838 73414 2884 73466
rect 2588 73412 2644 73414
rect 2668 73412 2724 73414
rect 2748 73412 2804 73414
rect 2828 73412 2884 73414
rect 2502 72664 2558 72720
rect 2870 72528 2926 72584
rect 1950 60424 2006 60480
rect 1858 57840 1914 57896
rect 1490 57296 1546 57352
rect 1582 56616 1638 56672
rect 1766 57024 1822 57080
rect 1490 54848 1546 54904
rect 1398 53216 1454 53272
rect 1582 52808 1638 52864
rect 1490 52536 1546 52592
rect 1398 51992 1454 52048
rect 1582 51584 1638 51640
rect 1490 51176 1546 51232
rect 1306 50904 1362 50960
rect 1122 23604 1124 23624
rect 1124 23604 1176 23624
rect 1176 23604 1178 23624
rect 1122 23568 1178 23604
rect 1582 50904 1638 50960
rect 1490 50496 1546 50552
rect 1398 49408 1454 49464
rect 1306 47912 1362 47968
rect 1398 47504 1454 47560
rect 1214 21392 1270 21448
rect 1214 19216 1270 19272
rect 1214 15000 1270 15056
rect 1214 11192 1270 11248
rect 1766 51312 1822 51368
rect 1674 50496 1730 50552
rect 1674 50360 1730 50416
rect 1674 49544 1730 49600
rect 1674 48864 1730 48920
rect 1766 48456 1822 48512
rect 1582 47776 1638 47832
rect 1582 47404 1584 47424
rect 1584 47404 1636 47424
rect 1636 47404 1638 47424
rect 1582 47368 1638 47404
rect 1582 45464 1638 45520
rect 1582 44784 1638 44840
rect 1766 47096 1822 47152
rect 1674 42472 1730 42528
rect 1490 41112 1546 41168
rect 1766 42336 1822 42392
rect 1674 40840 1730 40896
rect 1582 40568 1638 40624
rect 1582 38800 1638 38856
rect 1398 37576 1454 37632
rect 1582 35436 1584 35456
rect 1584 35436 1636 35456
rect 1636 35436 1638 35456
rect 1582 35400 1638 35436
rect 1766 40704 1822 40760
rect 1490 34992 1546 35048
rect 1674 34856 1730 34912
rect 1582 34584 1638 34640
rect 1398 32272 1454 32328
rect 1950 51176 2006 51232
rect 1950 50788 2006 50824
rect 1950 50768 1952 50788
rect 1952 50768 2004 50788
rect 2004 50768 2006 50788
rect 1950 50496 2006 50552
rect 1950 49680 2006 49736
rect 2134 61104 2190 61160
rect 2588 72378 2644 72380
rect 2668 72378 2724 72380
rect 2748 72378 2804 72380
rect 2828 72378 2884 72380
rect 2588 72326 2634 72378
rect 2634 72326 2644 72378
rect 2668 72326 2698 72378
rect 2698 72326 2710 72378
rect 2710 72326 2724 72378
rect 2748 72326 2762 72378
rect 2762 72326 2774 72378
rect 2774 72326 2804 72378
rect 2828 72326 2838 72378
rect 2838 72326 2884 72378
rect 2588 72324 2644 72326
rect 2668 72324 2724 72326
rect 2748 72324 2804 72326
rect 2828 72324 2884 72326
rect 2588 71290 2644 71292
rect 2668 71290 2724 71292
rect 2748 71290 2804 71292
rect 2828 71290 2884 71292
rect 2588 71238 2634 71290
rect 2634 71238 2644 71290
rect 2668 71238 2698 71290
rect 2698 71238 2710 71290
rect 2710 71238 2724 71290
rect 2748 71238 2762 71290
rect 2762 71238 2774 71290
rect 2774 71238 2804 71290
rect 2828 71238 2838 71290
rect 2838 71238 2884 71290
rect 2588 71236 2644 71238
rect 2668 71236 2724 71238
rect 2748 71236 2804 71238
rect 2828 71236 2884 71238
rect 2588 70202 2644 70204
rect 2668 70202 2724 70204
rect 2748 70202 2804 70204
rect 2828 70202 2884 70204
rect 2588 70150 2634 70202
rect 2634 70150 2644 70202
rect 2668 70150 2698 70202
rect 2698 70150 2710 70202
rect 2710 70150 2724 70202
rect 2748 70150 2762 70202
rect 2762 70150 2774 70202
rect 2774 70150 2804 70202
rect 2828 70150 2838 70202
rect 2838 70150 2884 70202
rect 2588 70148 2644 70150
rect 2668 70148 2724 70150
rect 2748 70148 2804 70150
rect 2828 70148 2884 70150
rect 2588 69114 2644 69116
rect 2668 69114 2724 69116
rect 2748 69114 2804 69116
rect 2828 69114 2884 69116
rect 2588 69062 2634 69114
rect 2634 69062 2644 69114
rect 2668 69062 2698 69114
rect 2698 69062 2710 69114
rect 2710 69062 2724 69114
rect 2748 69062 2762 69114
rect 2762 69062 2774 69114
rect 2774 69062 2804 69114
rect 2828 69062 2838 69114
rect 2838 69062 2884 69114
rect 2588 69060 2644 69062
rect 2668 69060 2724 69062
rect 2748 69060 2804 69062
rect 2828 69060 2884 69062
rect 2778 68584 2834 68640
rect 2588 68026 2644 68028
rect 2668 68026 2724 68028
rect 2748 68026 2804 68028
rect 2828 68026 2884 68028
rect 2588 67974 2634 68026
rect 2634 67974 2644 68026
rect 2668 67974 2698 68026
rect 2698 67974 2710 68026
rect 2710 67974 2724 68026
rect 2748 67974 2762 68026
rect 2762 67974 2774 68026
rect 2774 67974 2804 68026
rect 2828 67974 2838 68026
rect 2838 67974 2884 68026
rect 2588 67972 2644 67974
rect 2668 67972 2724 67974
rect 2748 67972 2804 67974
rect 2828 67972 2884 67974
rect 2962 67768 3018 67824
rect 2778 67632 2834 67688
rect 2588 66938 2644 66940
rect 2668 66938 2724 66940
rect 2748 66938 2804 66940
rect 2828 66938 2884 66940
rect 2588 66886 2634 66938
rect 2634 66886 2644 66938
rect 2668 66886 2698 66938
rect 2698 66886 2710 66938
rect 2710 66886 2724 66938
rect 2748 66886 2762 66938
rect 2762 66886 2774 66938
rect 2774 66886 2804 66938
rect 2828 66886 2838 66938
rect 2838 66886 2884 66938
rect 2588 66884 2644 66886
rect 2668 66884 2724 66886
rect 2748 66884 2804 66886
rect 2828 66884 2884 66886
rect 2778 66000 2834 66056
rect 2588 65850 2644 65852
rect 2668 65850 2724 65852
rect 2748 65850 2804 65852
rect 2828 65850 2884 65852
rect 2588 65798 2634 65850
rect 2634 65798 2644 65850
rect 2668 65798 2698 65850
rect 2698 65798 2710 65850
rect 2710 65798 2724 65850
rect 2748 65798 2762 65850
rect 2762 65798 2774 65850
rect 2774 65798 2804 65850
rect 2828 65798 2838 65850
rect 2838 65798 2884 65850
rect 2588 65796 2644 65798
rect 2668 65796 2724 65798
rect 2748 65796 2804 65798
rect 2828 65796 2884 65798
rect 3330 67632 3386 67688
rect 3054 65048 3110 65104
rect 2588 64762 2644 64764
rect 2668 64762 2724 64764
rect 2748 64762 2804 64764
rect 2828 64762 2884 64764
rect 2588 64710 2634 64762
rect 2634 64710 2644 64762
rect 2668 64710 2698 64762
rect 2698 64710 2710 64762
rect 2710 64710 2724 64762
rect 2748 64710 2762 64762
rect 2762 64710 2774 64762
rect 2774 64710 2804 64762
rect 2828 64710 2838 64762
rect 2838 64710 2884 64762
rect 2588 64708 2644 64710
rect 2668 64708 2724 64710
rect 2748 64708 2804 64710
rect 2828 64708 2884 64710
rect 3054 64368 3110 64424
rect 2502 63824 2558 63880
rect 2588 63674 2644 63676
rect 2668 63674 2724 63676
rect 2748 63674 2804 63676
rect 2828 63674 2884 63676
rect 2588 63622 2634 63674
rect 2634 63622 2644 63674
rect 2668 63622 2698 63674
rect 2698 63622 2710 63674
rect 2710 63622 2724 63674
rect 2748 63622 2762 63674
rect 2762 63622 2774 63674
rect 2774 63622 2804 63674
rect 2828 63622 2838 63674
rect 2838 63622 2884 63674
rect 2588 63620 2644 63622
rect 2668 63620 2724 63622
rect 2748 63620 2804 63622
rect 2828 63620 2884 63622
rect 2318 61784 2374 61840
rect 2318 61004 2320 61024
rect 2320 61004 2372 61024
rect 2372 61004 2374 61024
rect 2318 60968 2374 61004
rect 2318 60832 2374 60888
rect 2318 59608 2374 59664
rect 2318 58384 2374 58440
rect 2318 58248 2374 58304
rect 2870 63416 2926 63472
rect 2594 62908 2596 62928
rect 2596 62908 2648 62928
rect 2648 62908 2650 62928
rect 2594 62872 2650 62908
rect 3146 63960 3202 64016
rect 3054 63552 3110 63608
rect 2588 62586 2644 62588
rect 2668 62586 2724 62588
rect 2748 62586 2804 62588
rect 2828 62586 2884 62588
rect 2588 62534 2634 62586
rect 2634 62534 2644 62586
rect 2668 62534 2698 62586
rect 2698 62534 2710 62586
rect 2710 62534 2724 62586
rect 2748 62534 2762 62586
rect 2762 62534 2774 62586
rect 2774 62534 2804 62586
rect 2828 62534 2838 62586
rect 2838 62534 2884 62586
rect 2588 62532 2644 62534
rect 2668 62532 2724 62534
rect 2748 62532 2804 62534
rect 2828 62532 2884 62534
rect 2778 62192 2834 62248
rect 2594 61648 2650 61704
rect 2588 61498 2644 61500
rect 2668 61498 2724 61500
rect 2748 61498 2804 61500
rect 2828 61498 2884 61500
rect 2588 61446 2634 61498
rect 2634 61446 2644 61498
rect 2668 61446 2698 61498
rect 2698 61446 2710 61498
rect 2710 61446 2724 61498
rect 2748 61446 2762 61498
rect 2762 61446 2774 61498
rect 2774 61446 2804 61498
rect 2828 61446 2838 61498
rect 2838 61446 2884 61498
rect 2588 61444 2644 61446
rect 2668 61444 2724 61446
rect 2748 61444 2804 61446
rect 2828 61444 2884 61446
rect 3054 60716 3110 60752
rect 3054 60696 3056 60716
rect 3056 60696 3108 60716
rect 3108 60696 3110 60716
rect 2778 60580 2834 60616
rect 2778 60560 2780 60580
rect 2780 60560 2832 60580
rect 2832 60560 2834 60580
rect 2588 60410 2644 60412
rect 2668 60410 2724 60412
rect 2748 60410 2804 60412
rect 2828 60410 2884 60412
rect 2588 60358 2634 60410
rect 2634 60358 2644 60410
rect 2668 60358 2698 60410
rect 2698 60358 2710 60410
rect 2710 60358 2724 60410
rect 2748 60358 2762 60410
rect 2762 60358 2774 60410
rect 2774 60358 2804 60410
rect 2828 60358 2838 60410
rect 2838 60358 2884 60410
rect 2588 60356 2644 60358
rect 2668 60356 2724 60358
rect 2748 60356 2804 60358
rect 2828 60356 2884 60358
rect 2502 60152 2558 60208
rect 2410 57704 2466 57760
rect 2594 60016 2650 60072
rect 2588 59322 2644 59324
rect 2668 59322 2724 59324
rect 2748 59322 2804 59324
rect 2828 59322 2884 59324
rect 2588 59270 2634 59322
rect 2634 59270 2644 59322
rect 2668 59270 2698 59322
rect 2698 59270 2710 59322
rect 2710 59270 2724 59322
rect 2748 59270 2762 59322
rect 2762 59270 2774 59322
rect 2774 59270 2804 59322
rect 2828 59270 2838 59322
rect 2838 59270 2884 59322
rect 2588 59268 2644 59270
rect 2668 59268 2724 59270
rect 2748 59268 2804 59270
rect 2828 59268 2884 59270
rect 2686 59064 2742 59120
rect 2686 58384 2742 58440
rect 2588 58234 2644 58236
rect 2668 58234 2724 58236
rect 2748 58234 2804 58236
rect 2828 58234 2884 58236
rect 2588 58182 2634 58234
rect 2634 58182 2644 58234
rect 2668 58182 2698 58234
rect 2698 58182 2710 58234
rect 2710 58182 2724 58234
rect 2748 58182 2762 58234
rect 2762 58182 2774 58234
rect 2774 58182 2804 58234
rect 2828 58182 2838 58234
rect 2838 58182 2884 58234
rect 2588 58180 2644 58182
rect 2668 58180 2724 58182
rect 2748 58180 2804 58182
rect 2828 58180 2884 58182
rect 2594 57976 2650 58032
rect 2778 57976 2834 58032
rect 2686 57568 2742 57624
rect 2594 57296 2650 57352
rect 2318 56752 2374 56808
rect 2318 55256 2374 55312
rect 2318 54848 2374 54904
rect 2318 53760 2374 53816
rect 2318 53100 2374 53136
rect 2318 53080 2320 53100
rect 2320 53080 2372 53100
rect 2372 53080 2374 53100
rect 2318 52400 2374 52456
rect 2588 57146 2644 57148
rect 2668 57146 2724 57148
rect 2748 57146 2804 57148
rect 2828 57146 2884 57148
rect 2588 57094 2634 57146
rect 2634 57094 2644 57146
rect 2668 57094 2698 57146
rect 2698 57094 2710 57146
rect 2710 57094 2724 57146
rect 2748 57094 2762 57146
rect 2762 57094 2774 57146
rect 2774 57094 2804 57146
rect 2828 57094 2838 57146
rect 2838 57094 2884 57146
rect 2588 57092 2644 57094
rect 2668 57092 2724 57094
rect 2748 57092 2804 57094
rect 2828 57092 2884 57094
rect 3146 59064 3202 59120
rect 3054 58828 3056 58848
rect 3056 58828 3108 58848
rect 3108 58828 3110 58848
rect 3054 58792 3110 58828
rect 3054 57704 3110 57760
rect 3146 57568 3202 57624
rect 3054 57296 3110 57352
rect 2502 56888 2558 56944
rect 2502 56616 2558 56672
rect 2594 56480 2650 56536
rect 2778 56480 2834 56536
rect 2962 56364 3018 56400
rect 2962 56344 2964 56364
rect 2964 56344 3016 56364
rect 3016 56344 3018 56364
rect 2588 56058 2644 56060
rect 2668 56058 2724 56060
rect 2748 56058 2804 56060
rect 2828 56058 2884 56060
rect 2588 56006 2634 56058
rect 2634 56006 2644 56058
rect 2668 56006 2698 56058
rect 2698 56006 2710 56058
rect 2710 56006 2724 56058
rect 2748 56006 2762 56058
rect 2762 56006 2774 56058
rect 2774 56006 2804 56058
rect 2828 56006 2838 56058
rect 2838 56006 2884 56058
rect 2588 56004 2644 56006
rect 2668 56004 2724 56006
rect 2748 56004 2804 56006
rect 2828 56004 2884 56006
rect 2502 55664 2558 55720
rect 3054 55800 3110 55856
rect 3054 55528 3110 55584
rect 2588 54970 2644 54972
rect 2668 54970 2724 54972
rect 2748 54970 2804 54972
rect 2828 54970 2884 54972
rect 2588 54918 2634 54970
rect 2634 54918 2644 54970
rect 2668 54918 2698 54970
rect 2698 54918 2710 54970
rect 2710 54918 2724 54970
rect 2748 54918 2762 54970
rect 2762 54918 2774 54970
rect 2774 54918 2804 54970
rect 2828 54918 2838 54970
rect 2838 54918 2884 54970
rect 2588 54916 2644 54918
rect 2668 54916 2724 54918
rect 2748 54916 2804 54918
rect 2828 54916 2884 54918
rect 2502 54576 2558 54632
rect 2962 54304 3018 54360
rect 2778 54168 2834 54224
rect 2686 54032 2742 54088
rect 2588 53882 2644 53884
rect 2668 53882 2724 53884
rect 2748 53882 2804 53884
rect 2828 53882 2884 53884
rect 2588 53830 2634 53882
rect 2634 53830 2644 53882
rect 2668 53830 2698 53882
rect 2698 53830 2710 53882
rect 2710 53830 2724 53882
rect 2748 53830 2762 53882
rect 2762 53830 2774 53882
rect 2774 53830 2804 53882
rect 2828 53830 2838 53882
rect 2838 53830 2884 53882
rect 2588 53828 2644 53830
rect 2668 53828 2724 53830
rect 2748 53828 2804 53830
rect 2828 53828 2884 53830
rect 2410 52128 2466 52184
rect 2318 51992 2374 52048
rect 2588 52794 2644 52796
rect 2668 52794 2724 52796
rect 2748 52794 2804 52796
rect 2828 52794 2884 52796
rect 2588 52742 2634 52794
rect 2634 52742 2644 52794
rect 2668 52742 2698 52794
rect 2698 52742 2710 52794
rect 2710 52742 2724 52794
rect 2748 52742 2762 52794
rect 2762 52742 2774 52794
rect 2774 52742 2804 52794
rect 2828 52742 2838 52794
rect 2838 52742 2884 52794
rect 2588 52740 2644 52742
rect 2668 52740 2724 52742
rect 2748 52740 2804 52742
rect 2828 52740 2884 52742
rect 2502 51892 2504 51912
rect 2504 51892 2556 51912
rect 2556 51892 2558 51912
rect 2502 51856 2558 51892
rect 2318 51312 2374 51368
rect 2318 49952 2374 50008
rect 2226 48592 2282 48648
rect 2588 51706 2644 51708
rect 2668 51706 2724 51708
rect 2748 51706 2804 51708
rect 2828 51706 2884 51708
rect 2588 51654 2634 51706
rect 2634 51654 2644 51706
rect 2668 51654 2698 51706
rect 2698 51654 2710 51706
rect 2710 51654 2724 51706
rect 2748 51654 2762 51706
rect 2762 51654 2774 51706
rect 2774 51654 2804 51706
rect 2828 51654 2838 51706
rect 2838 51654 2884 51706
rect 2588 51652 2644 51654
rect 2668 51652 2724 51654
rect 2748 51652 2804 51654
rect 2828 51652 2884 51654
rect 3054 51448 3110 51504
rect 3330 64812 3332 64832
rect 3332 64812 3384 64832
rect 3384 64812 3386 64832
rect 3330 64776 3386 64812
rect 3330 63008 3386 63064
rect 3238 53624 3294 53680
rect 3422 55120 3478 55176
rect 2588 50618 2644 50620
rect 2668 50618 2724 50620
rect 2748 50618 2804 50620
rect 2828 50618 2884 50620
rect 2588 50566 2634 50618
rect 2634 50566 2644 50618
rect 2668 50566 2698 50618
rect 2698 50566 2710 50618
rect 2710 50566 2724 50618
rect 2748 50566 2762 50618
rect 2762 50566 2774 50618
rect 2774 50566 2804 50618
rect 2828 50566 2838 50618
rect 2838 50566 2884 50618
rect 2588 50564 2644 50566
rect 2668 50564 2724 50566
rect 2748 50564 2804 50566
rect 2828 50564 2884 50566
rect 2778 49816 2834 49872
rect 2588 49530 2644 49532
rect 2668 49530 2724 49532
rect 2748 49530 2804 49532
rect 2828 49530 2884 49532
rect 2588 49478 2634 49530
rect 2634 49478 2644 49530
rect 2668 49478 2698 49530
rect 2698 49478 2710 49530
rect 2710 49478 2724 49530
rect 2748 49478 2762 49530
rect 2762 49478 2774 49530
rect 2774 49478 2804 49530
rect 2828 49478 2838 49530
rect 2838 49478 2884 49530
rect 2588 49476 2644 49478
rect 2668 49476 2724 49478
rect 2748 49476 2804 49478
rect 2828 49476 2884 49478
rect 2686 48864 2742 48920
rect 3146 51312 3202 51368
rect 3606 75384 3662 75440
rect 3054 48884 3110 48920
rect 3054 48864 3056 48884
rect 3056 48864 3108 48884
rect 3108 48864 3110 48884
rect 3238 50768 3294 50824
rect 2778 48592 2834 48648
rect 2588 48442 2644 48444
rect 2668 48442 2724 48444
rect 2748 48442 2804 48444
rect 2828 48442 2884 48444
rect 2588 48390 2634 48442
rect 2634 48390 2644 48442
rect 2668 48390 2698 48442
rect 2698 48390 2710 48442
rect 2710 48390 2724 48442
rect 2748 48390 2762 48442
rect 2762 48390 2774 48442
rect 2774 48390 2804 48442
rect 2828 48390 2838 48442
rect 2838 48390 2884 48442
rect 2588 48388 2644 48390
rect 2668 48388 2724 48390
rect 2748 48388 2804 48390
rect 2828 48388 2884 48390
rect 2318 48320 2374 48376
rect 2962 48320 3018 48376
rect 2588 47354 2644 47356
rect 2668 47354 2724 47356
rect 2748 47354 2804 47356
rect 2828 47354 2884 47356
rect 2588 47302 2634 47354
rect 2634 47302 2644 47354
rect 2668 47302 2698 47354
rect 2698 47302 2710 47354
rect 2710 47302 2724 47354
rect 2748 47302 2762 47354
rect 2762 47302 2774 47354
rect 2774 47302 2804 47354
rect 2828 47302 2838 47354
rect 2838 47302 2884 47354
rect 2588 47300 2644 47302
rect 2668 47300 2724 47302
rect 2748 47300 2804 47302
rect 2828 47300 2884 47302
rect 2318 46552 2374 46608
rect 2318 46416 2374 46472
rect 2318 45464 2374 45520
rect 2318 44784 2374 44840
rect 2502 46416 2558 46472
rect 2588 46266 2644 46268
rect 2668 46266 2724 46268
rect 2748 46266 2804 46268
rect 2828 46266 2884 46268
rect 2588 46214 2634 46266
rect 2634 46214 2644 46266
rect 2668 46214 2698 46266
rect 2698 46214 2710 46266
rect 2710 46214 2724 46266
rect 2748 46214 2762 46266
rect 2762 46214 2774 46266
rect 2774 46214 2804 46266
rect 2828 46214 2838 46266
rect 2838 46214 2884 46266
rect 2588 46212 2644 46214
rect 2668 46212 2724 46214
rect 2748 46212 2804 46214
rect 2828 46212 2884 46214
rect 2502 46008 2558 46064
rect 2502 45872 2558 45928
rect 2870 45908 2872 45928
rect 2872 45908 2924 45928
rect 2924 45908 2926 45928
rect 2870 45872 2926 45908
rect 2870 45484 2926 45520
rect 2870 45464 2872 45484
rect 2872 45464 2924 45484
rect 2924 45464 2926 45484
rect 2594 45348 2650 45384
rect 2594 45328 2596 45348
rect 2596 45328 2648 45348
rect 2648 45328 2650 45348
rect 3054 45772 3056 45792
rect 3056 45772 3108 45792
rect 3108 45772 3110 45792
rect 3054 45736 3110 45772
rect 2588 45178 2644 45180
rect 2668 45178 2724 45180
rect 2748 45178 2804 45180
rect 2828 45178 2884 45180
rect 2588 45126 2634 45178
rect 2634 45126 2644 45178
rect 2668 45126 2698 45178
rect 2698 45126 2710 45178
rect 2710 45126 2724 45178
rect 2748 45126 2762 45178
rect 2762 45126 2774 45178
rect 2774 45126 2804 45178
rect 2828 45126 2838 45178
rect 2838 45126 2884 45178
rect 2588 45124 2644 45126
rect 2668 45124 2724 45126
rect 2748 45124 2804 45126
rect 2828 45124 2884 45126
rect 2962 44684 2964 44704
rect 2964 44684 3016 44704
rect 3016 44684 3018 44704
rect 2962 44648 3018 44684
rect 2588 44090 2644 44092
rect 2668 44090 2724 44092
rect 2748 44090 2804 44092
rect 2828 44090 2884 44092
rect 2588 44038 2634 44090
rect 2634 44038 2644 44090
rect 2668 44038 2698 44090
rect 2698 44038 2710 44090
rect 2710 44038 2724 44090
rect 2748 44038 2762 44090
rect 2762 44038 2774 44090
rect 2774 44038 2804 44090
rect 2828 44038 2838 44090
rect 2838 44038 2884 44090
rect 2588 44036 2644 44038
rect 2668 44036 2724 44038
rect 2748 44036 2804 44038
rect 2828 44036 2884 44038
rect 3146 44240 3202 44296
rect 3146 43832 3202 43888
rect 3054 43424 3110 43480
rect 2588 43002 2644 43004
rect 2668 43002 2724 43004
rect 2748 43002 2804 43004
rect 2828 43002 2884 43004
rect 2588 42950 2634 43002
rect 2634 42950 2644 43002
rect 2668 42950 2698 43002
rect 2698 42950 2710 43002
rect 2710 42950 2724 43002
rect 2748 42950 2762 43002
rect 2762 42950 2774 43002
rect 2774 42950 2804 43002
rect 2828 42950 2838 43002
rect 2838 42950 2884 43002
rect 2588 42948 2644 42950
rect 2668 42948 2724 42950
rect 2748 42948 2804 42950
rect 2828 42948 2884 42950
rect 2962 42880 3018 42936
rect 2870 42744 2926 42800
rect 2778 42200 2834 42256
rect 2502 42064 2558 42120
rect 2588 41914 2644 41916
rect 2668 41914 2724 41916
rect 2748 41914 2804 41916
rect 2828 41914 2884 41916
rect 2588 41862 2634 41914
rect 2634 41862 2644 41914
rect 2668 41862 2698 41914
rect 2698 41862 2710 41914
rect 2710 41862 2724 41914
rect 2748 41862 2762 41914
rect 2762 41862 2774 41914
rect 2774 41862 2804 41914
rect 2828 41862 2838 41914
rect 2838 41862 2884 41914
rect 2588 41860 2644 41862
rect 2668 41860 2724 41862
rect 2748 41860 2804 41862
rect 2828 41860 2884 41862
rect 2410 41520 2466 41576
rect 2318 41420 2320 41440
rect 2320 41420 2372 41440
rect 2372 41420 2374 41440
rect 2318 41384 2374 41420
rect 2226 41248 2282 41304
rect 2226 41112 2282 41168
rect 2134 40024 2190 40080
rect 2778 40996 2834 41032
rect 2778 40976 2780 40996
rect 2780 40976 2832 40996
rect 2832 40976 2834 40996
rect 2588 40826 2644 40828
rect 2668 40826 2724 40828
rect 2748 40826 2804 40828
rect 2828 40826 2884 40828
rect 2588 40774 2634 40826
rect 2634 40774 2644 40826
rect 2668 40774 2698 40826
rect 2698 40774 2710 40826
rect 2710 40774 2724 40826
rect 2748 40774 2762 40826
rect 2762 40774 2774 40826
rect 2774 40774 2804 40826
rect 2828 40774 2838 40826
rect 2838 40774 2884 40826
rect 2588 40772 2644 40774
rect 2668 40772 2724 40774
rect 2748 40772 2804 40774
rect 2828 40772 2884 40774
rect 2778 40044 2834 40080
rect 2778 40024 2780 40044
rect 2780 40024 2832 40044
rect 2832 40024 2834 40044
rect 3054 41656 3110 41712
rect 3054 41012 3056 41032
rect 3056 41012 3108 41032
rect 3108 41012 3110 41032
rect 3054 40976 3110 41012
rect 2870 39908 2926 39944
rect 2870 39888 2872 39908
rect 2872 39888 2924 39908
rect 2924 39888 2926 39908
rect 2588 39738 2644 39740
rect 2668 39738 2724 39740
rect 2748 39738 2804 39740
rect 2828 39738 2884 39740
rect 2588 39686 2634 39738
rect 2634 39686 2644 39738
rect 2668 39686 2698 39738
rect 2698 39686 2710 39738
rect 2710 39686 2724 39738
rect 2748 39686 2762 39738
rect 2762 39686 2774 39738
rect 2774 39686 2804 39738
rect 2828 39686 2838 39738
rect 2838 39686 2884 39738
rect 2588 39684 2644 39686
rect 2668 39684 2724 39686
rect 2748 39684 2804 39686
rect 2828 39684 2884 39686
rect 1582 32000 1638 32056
rect 1490 29824 1546 29880
rect 1490 28192 1546 28248
rect 1490 28056 1546 28112
rect 1398 27784 1454 27840
rect 1398 27412 1400 27432
rect 1400 27412 1452 27432
rect 1452 27412 1454 27432
rect 1398 27376 1454 27412
rect 1950 32136 2006 32192
rect 2318 34176 2374 34232
rect 2226 33224 2282 33280
rect 2410 33532 2412 33552
rect 2412 33532 2464 33552
rect 2464 33532 2466 33552
rect 2410 33496 2466 33532
rect 2134 31320 2190 31376
rect 2042 29960 2098 30016
rect 2042 29824 2098 29880
rect 1858 29416 1914 29472
rect 1858 29280 1914 29336
rect 1950 28872 2006 28928
rect 2134 28872 2190 28928
rect 2318 31048 2374 31104
rect 2318 28872 2374 28928
rect 1766 28636 1768 28656
rect 1768 28636 1820 28656
rect 1820 28636 1822 28656
rect 1766 28600 1822 28636
rect 1674 26852 1730 26888
rect 1674 26832 1676 26852
rect 1676 26832 1728 26852
rect 1728 26832 1730 26852
rect 1398 23060 1400 23080
rect 1400 23060 1452 23080
rect 1452 23060 1454 23080
rect 1398 23024 1454 23060
rect 1398 21800 1454 21856
rect 1398 20984 1454 21040
rect 1398 20168 1454 20224
rect 1398 19624 1454 19680
rect 2318 28736 2374 28792
rect 3054 38936 3110 38992
rect 2870 38800 2926 38856
rect 2588 38650 2644 38652
rect 2668 38650 2724 38652
rect 2748 38650 2804 38652
rect 2828 38650 2884 38652
rect 2588 38598 2634 38650
rect 2634 38598 2644 38650
rect 2668 38598 2698 38650
rect 2698 38598 2710 38650
rect 2710 38598 2724 38650
rect 2748 38598 2762 38650
rect 2762 38598 2774 38650
rect 2774 38598 2804 38650
rect 2828 38598 2838 38650
rect 2838 38598 2884 38650
rect 2588 38596 2644 38598
rect 2668 38596 2724 38598
rect 2748 38596 2804 38598
rect 2828 38596 2884 38598
rect 2778 38256 2834 38312
rect 2594 38120 2650 38176
rect 2962 37984 3018 38040
rect 2588 37562 2644 37564
rect 2668 37562 2724 37564
rect 2748 37562 2804 37564
rect 2828 37562 2884 37564
rect 2588 37510 2634 37562
rect 2634 37510 2644 37562
rect 2668 37510 2698 37562
rect 2698 37510 2710 37562
rect 2710 37510 2724 37562
rect 2748 37510 2762 37562
rect 2762 37510 2774 37562
rect 2774 37510 2804 37562
rect 2828 37510 2838 37562
rect 2838 37510 2884 37562
rect 2588 37508 2644 37510
rect 2668 37508 2724 37510
rect 2748 37508 2804 37510
rect 2828 37508 2884 37510
rect 2686 37304 2742 37360
rect 2588 36474 2644 36476
rect 2668 36474 2724 36476
rect 2748 36474 2804 36476
rect 2828 36474 2884 36476
rect 2588 36422 2634 36474
rect 2634 36422 2644 36474
rect 2668 36422 2698 36474
rect 2698 36422 2710 36474
rect 2710 36422 2724 36474
rect 2748 36422 2762 36474
rect 2762 36422 2774 36474
rect 2774 36422 2804 36474
rect 2828 36422 2838 36474
rect 2838 36422 2884 36474
rect 2588 36420 2644 36422
rect 2668 36420 2724 36422
rect 2748 36420 2804 36422
rect 2828 36420 2884 36422
rect 2778 35808 2834 35864
rect 2588 35386 2644 35388
rect 2668 35386 2724 35388
rect 2748 35386 2804 35388
rect 2828 35386 2884 35388
rect 2588 35334 2634 35386
rect 2634 35334 2644 35386
rect 2668 35334 2698 35386
rect 2698 35334 2710 35386
rect 2710 35334 2724 35386
rect 2748 35334 2762 35386
rect 2762 35334 2774 35386
rect 2774 35334 2804 35386
rect 2828 35334 2838 35386
rect 2838 35334 2884 35386
rect 2588 35332 2644 35334
rect 2668 35332 2724 35334
rect 2748 35332 2804 35334
rect 2828 35332 2884 35334
rect 2588 34298 2644 34300
rect 2668 34298 2724 34300
rect 2748 34298 2804 34300
rect 2828 34298 2884 34300
rect 2588 34246 2634 34298
rect 2634 34246 2644 34298
rect 2668 34246 2698 34298
rect 2698 34246 2710 34298
rect 2710 34246 2724 34298
rect 2748 34246 2762 34298
rect 2762 34246 2774 34298
rect 2774 34246 2804 34298
rect 2828 34246 2838 34298
rect 2838 34246 2884 34298
rect 2588 34244 2644 34246
rect 2668 34244 2724 34246
rect 2748 34244 2804 34246
rect 2828 34244 2884 34246
rect 3054 33768 3110 33824
rect 3054 33496 3110 33552
rect 2588 33210 2644 33212
rect 2668 33210 2724 33212
rect 2748 33210 2804 33212
rect 2828 33210 2884 33212
rect 2588 33158 2634 33210
rect 2634 33158 2644 33210
rect 2668 33158 2698 33210
rect 2698 33158 2710 33210
rect 2710 33158 2724 33210
rect 2748 33158 2762 33210
rect 2762 33158 2774 33210
rect 2774 33158 2804 33210
rect 2828 33158 2838 33210
rect 2838 33158 2884 33210
rect 2588 33156 2644 33158
rect 2668 33156 2724 33158
rect 2748 33156 2804 33158
rect 2828 33156 2884 33158
rect 2588 32122 2644 32124
rect 2668 32122 2724 32124
rect 2748 32122 2804 32124
rect 2828 32122 2884 32124
rect 2588 32070 2634 32122
rect 2634 32070 2644 32122
rect 2668 32070 2698 32122
rect 2698 32070 2710 32122
rect 2710 32070 2724 32122
rect 2748 32070 2762 32122
rect 2762 32070 2774 32122
rect 2774 32070 2804 32122
rect 2828 32070 2838 32122
rect 2838 32070 2884 32122
rect 2588 32068 2644 32070
rect 2668 32068 2724 32070
rect 2748 32068 2804 32070
rect 2828 32068 2884 32070
rect 3330 49272 3386 49328
rect 3698 62756 3754 62792
rect 3698 62736 3700 62756
rect 3700 62736 3752 62756
rect 3752 62736 3754 62756
rect 3698 62600 3754 62656
rect 5852 76730 5908 76732
rect 5932 76730 5988 76732
rect 6012 76730 6068 76732
rect 6092 76730 6148 76732
rect 5852 76678 5898 76730
rect 5898 76678 5908 76730
rect 5932 76678 5962 76730
rect 5962 76678 5974 76730
rect 5974 76678 5988 76730
rect 6012 76678 6026 76730
rect 6026 76678 6038 76730
rect 6038 76678 6068 76730
rect 6092 76678 6102 76730
rect 6102 76678 6148 76730
rect 5852 76676 5908 76678
rect 5932 76676 5988 76678
rect 6012 76676 6068 76678
rect 6092 76676 6148 76678
rect 4220 76186 4276 76188
rect 4300 76186 4356 76188
rect 4380 76186 4436 76188
rect 4460 76186 4516 76188
rect 4220 76134 4266 76186
rect 4266 76134 4276 76186
rect 4300 76134 4330 76186
rect 4330 76134 4342 76186
rect 4342 76134 4356 76186
rect 4380 76134 4394 76186
rect 4394 76134 4406 76186
rect 4406 76134 4436 76186
rect 4460 76134 4470 76186
rect 4470 76134 4516 76186
rect 4220 76132 4276 76134
rect 4300 76132 4356 76134
rect 4380 76132 4436 76134
rect 4460 76132 4516 76134
rect 7484 76186 7540 76188
rect 7564 76186 7620 76188
rect 7644 76186 7700 76188
rect 7724 76186 7780 76188
rect 7484 76134 7530 76186
rect 7530 76134 7540 76186
rect 7564 76134 7594 76186
rect 7594 76134 7606 76186
rect 7606 76134 7620 76186
rect 7644 76134 7658 76186
rect 7658 76134 7670 76186
rect 7670 76134 7700 76186
rect 7724 76134 7734 76186
rect 7734 76134 7780 76186
rect 7484 76132 7540 76134
rect 7564 76132 7620 76134
rect 7644 76132 7700 76134
rect 7724 76132 7780 76134
rect 5852 75642 5908 75644
rect 5932 75642 5988 75644
rect 6012 75642 6068 75644
rect 6092 75642 6148 75644
rect 5852 75590 5898 75642
rect 5898 75590 5908 75642
rect 5932 75590 5962 75642
rect 5962 75590 5974 75642
rect 5974 75590 5988 75642
rect 6012 75590 6026 75642
rect 6026 75590 6038 75642
rect 6038 75590 6068 75642
rect 6092 75590 6102 75642
rect 6102 75590 6148 75642
rect 5852 75588 5908 75590
rect 5932 75588 5988 75590
rect 6012 75588 6068 75590
rect 6092 75588 6148 75590
rect 4220 75098 4276 75100
rect 4300 75098 4356 75100
rect 4380 75098 4436 75100
rect 4460 75098 4516 75100
rect 4220 75046 4266 75098
rect 4266 75046 4276 75098
rect 4300 75046 4330 75098
rect 4330 75046 4342 75098
rect 4342 75046 4356 75098
rect 4380 75046 4394 75098
rect 4394 75046 4406 75098
rect 4406 75046 4436 75098
rect 4460 75046 4470 75098
rect 4470 75046 4516 75098
rect 4220 75044 4276 75046
rect 4300 75044 4356 75046
rect 4380 75044 4436 75046
rect 4460 75044 4516 75046
rect 7484 75098 7540 75100
rect 7564 75098 7620 75100
rect 7644 75098 7700 75100
rect 7724 75098 7780 75100
rect 7484 75046 7530 75098
rect 7530 75046 7540 75098
rect 7564 75046 7594 75098
rect 7594 75046 7606 75098
rect 7606 75046 7620 75098
rect 7644 75046 7658 75098
rect 7658 75046 7670 75098
rect 7670 75046 7700 75098
rect 7724 75046 7734 75098
rect 7734 75046 7780 75098
rect 7484 75044 7540 75046
rect 7564 75044 7620 75046
rect 7644 75044 7700 75046
rect 7724 75044 7780 75046
rect 9402 77152 9458 77208
rect 9116 76730 9172 76732
rect 9196 76730 9252 76732
rect 9276 76730 9332 76732
rect 9356 76730 9412 76732
rect 9116 76678 9162 76730
rect 9162 76678 9172 76730
rect 9196 76678 9226 76730
rect 9226 76678 9238 76730
rect 9238 76678 9252 76730
rect 9276 76678 9290 76730
rect 9290 76678 9302 76730
rect 9302 76678 9332 76730
rect 9356 76678 9366 76730
rect 9366 76678 9412 76730
rect 9116 76676 9172 76678
rect 9196 76676 9252 76678
rect 9276 76676 9332 76678
rect 9356 76676 9412 76678
rect 9116 75642 9172 75644
rect 9196 75642 9252 75644
rect 9276 75642 9332 75644
rect 9356 75642 9412 75644
rect 9116 75590 9162 75642
rect 9162 75590 9172 75642
rect 9196 75590 9226 75642
rect 9226 75590 9238 75642
rect 9238 75590 9252 75642
rect 9276 75590 9290 75642
rect 9290 75590 9302 75642
rect 9302 75590 9332 75642
rect 9356 75590 9366 75642
rect 9366 75590 9412 75642
rect 9116 75588 9172 75590
rect 9196 75588 9252 75590
rect 9276 75588 9332 75590
rect 9356 75588 9412 75590
rect 5852 74554 5908 74556
rect 5932 74554 5988 74556
rect 6012 74554 6068 74556
rect 6092 74554 6148 74556
rect 5852 74502 5898 74554
rect 5898 74502 5908 74554
rect 5932 74502 5962 74554
rect 5962 74502 5974 74554
rect 5974 74502 5988 74554
rect 6012 74502 6026 74554
rect 6026 74502 6038 74554
rect 6038 74502 6068 74554
rect 6092 74502 6102 74554
rect 6102 74502 6148 74554
rect 5852 74500 5908 74502
rect 5932 74500 5988 74502
rect 6012 74500 6068 74502
rect 6092 74500 6148 74502
rect 9116 74554 9172 74556
rect 9196 74554 9252 74556
rect 9276 74554 9332 74556
rect 9356 74554 9412 74556
rect 9116 74502 9162 74554
rect 9162 74502 9172 74554
rect 9196 74502 9226 74554
rect 9226 74502 9238 74554
rect 9238 74502 9252 74554
rect 9276 74502 9290 74554
rect 9290 74502 9302 74554
rect 9302 74502 9332 74554
rect 9356 74502 9366 74554
rect 9366 74502 9412 74554
rect 9116 74500 9172 74502
rect 9196 74500 9252 74502
rect 9276 74500 9332 74502
rect 9356 74500 9412 74502
rect 4220 74010 4276 74012
rect 4300 74010 4356 74012
rect 4380 74010 4436 74012
rect 4460 74010 4516 74012
rect 4220 73958 4266 74010
rect 4266 73958 4276 74010
rect 4300 73958 4330 74010
rect 4330 73958 4342 74010
rect 4342 73958 4356 74010
rect 4380 73958 4394 74010
rect 4394 73958 4406 74010
rect 4406 73958 4436 74010
rect 4460 73958 4470 74010
rect 4470 73958 4516 74010
rect 4220 73956 4276 73958
rect 4300 73956 4356 73958
rect 4380 73956 4436 73958
rect 4460 73956 4516 73958
rect 7484 74010 7540 74012
rect 7564 74010 7620 74012
rect 7644 74010 7700 74012
rect 7724 74010 7780 74012
rect 7484 73958 7530 74010
rect 7530 73958 7540 74010
rect 7564 73958 7594 74010
rect 7594 73958 7606 74010
rect 7606 73958 7620 74010
rect 7644 73958 7658 74010
rect 7658 73958 7670 74010
rect 7670 73958 7700 74010
rect 7724 73958 7734 74010
rect 7734 73958 7780 74010
rect 7484 73956 7540 73958
rect 7564 73956 7620 73958
rect 7644 73956 7700 73958
rect 7724 73956 7780 73958
rect 5852 73466 5908 73468
rect 5932 73466 5988 73468
rect 6012 73466 6068 73468
rect 6092 73466 6148 73468
rect 5852 73414 5898 73466
rect 5898 73414 5908 73466
rect 5932 73414 5962 73466
rect 5962 73414 5974 73466
rect 5974 73414 5988 73466
rect 6012 73414 6026 73466
rect 6026 73414 6038 73466
rect 6038 73414 6068 73466
rect 6092 73414 6102 73466
rect 6102 73414 6148 73466
rect 5852 73412 5908 73414
rect 5932 73412 5988 73414
rect 6012 73412 6068 73414
rect 6092 73412 6148 73414
rect 9116 73466 9172 73468
rect 9196 73466 9252 73468
rect 9276 73466 9332 73468
rect 9356 73466 9412 73468
rect 9116 73414 9162 73466
rect 9162 73414 9172 73466
rect 9196 73414 9226 73466
rect 9226 73414 9238 73466
rect 9238 73414 9252 73466
rect 9276 73414 9290 73466
rect 9290 73414 9302 73466
rect 9302 73414 9332 73466
rect 9356 73414 9366 73466
rect 9366 73414 9412 73466
rect 9116 73412 9172 73414
rect 9196 73412 9252 73414
rect 9276 73412 9332 73414
rect 9356 73412 9412 73414
rect 4220 72922 4276 72924
rect 4300 72922 4356 72924
rect 4380 72922 4436 72924
rect 4460 72922 4516 72924
rect 4220 72870 4266 72922
rect 4266 72870 4276 72922
rect 4300 72870 4330 72922
rect 4330 72870 4342 72922
rect 4342 72870 4356 72922
rect 4380 72870 4394 72922
rect 4394 72870 4406 72922
rect 4406 72870 4436 72922
rect 4460 72870 4470 72922
rect 4470 72870 4516 72922
rect 4220 72868 4276 72870
rect 4300 72868 4356 72870
rect 4380 72868 4436 72870
rect 4460 72868 4516 72870
rect 4220 71834 4276 71836
rect 4300 71834 4356 71836
rect 4380 71834 4436 71836
rect 4460 71834 4516 71836
rect 4220 71782 4266 71834
rect 4266 71782 4276 71834
rect 4300 71782 4330 71834
rect 4330 71782 4342 71834
rect 4342 71782 4356 71834
rect 4380 71782 4394 71834
rect 4394 71782 4406 71834
rect 4406 71782 4436 71834
rect 4460 71782 4470 71834
rect 4470 71782 4516 71834
rect 4220 71780 4276 71782
rect 4300 71780 4356 71782
rect 4380 71780 4436 71782
rect 4460 71780 4516 71782
rect 4220 70746 4276 70748
rect 4300 70746 4356 70748
rect 4380 70746 4436 70748
rect 4460 70746 4516 70748
rect 4220 70694 4266 70746
rect 4266 70694 4276 70746
rect 4300 70694 4330 70746
rect 4330 70694 4342 70746
rect 4342 70694 4356 70746
rect 4380 70694 4394 70746
rect 4394 70694 4406 70746
rect 4406 70694 4436 70746
rect 4460 70694 4470 70746
rect 4470 70694 4516 70746
rect 4220 70692 4276 70694
rect 4300 70692 4356 70694
rect 4380 70692 4436 70694
rect 4460 70692 4516 70694
rect 4220 69658 4276 69660
rect 4300 69658 4356 69660
rect 4380 69658 4436 69660
rect 4460 69658 4516 69660
rect 4220 69606 4266 69658
rect 4266 69606 4276 69658
rect 4300 69606 4330 69658
rect 4330 69606 4342 69658
rect 4342 69606 4356 69658
rect 4380 69606 4394 69658
rect 4394 69606 4406 69658
rect 4406 69606 4436 69658
rect 4460 69606 4470 69658
rect 4470 69606 4516 69658
rect 4220 69604 4276 69606
rect 4300 69604 4356 69606
rect 4380 69604 4436 69606
rect 4460 69604 4516 69606
rect 4220 68570 4276 68572
rect 4300 68570 4356 68572
rect 4380 68570 4436 68572
rect 4460 68570 4516 68572
rect 4220 68518 4266 68570
rect 4266 68518 4276 68570
rect 4300 68518 4330 68570
rect 4330 68518 4342 68570
rect 4342 68518 4356 68570
rect 4380 68518 4394 68570
rect 4394 68518 4406 68570
rect 4406 68518 4436 68570
rect 4460 68518 4470 68570
rect 4470 68518 4516 68570
rect 4220 68516 4276 68518
rect 4300 68516 4356 68518
rect 4380 68516 4436 68518
rect 4460 68516 4516 68518
rect 4220 67482 4276 67484
rect 4300 67482 4356 67484
rect 4380 67482 4436 67484
rect 4460 67482 4516 67484
rect 4220 67430 4266 67482
rect 4266 67430 4276 67482
rect 4300 67430 4330 67482
rect 4330 67430 4342 67482
rect 4342 67430 4356 67482
rect 4380 67430 4394 67482
rect 4394 67430 4406 67482
rect 4406 67430 4436 67482
rect 4460 67430 4470 67482
rect 4470 67430 4516 67482
rect 4220 67428 4276 67430
rect 4300 67428 4356 67430
rect 4380 67428 4436 67430
rect 4460 67428 4516 67430
rect 4220 66394 4276 66396
rect 4300 66394 4356 66396
rect 4380 66394 4436 66396
rect 4460 66394 4516 66396
rect 4220 66342 4266 66394
rect 4266 66342 4276 66394
rect 4300 66342 4330 66394
rect 4330 66342 4342 66394
rect 4342 66342 4356 66394
rect 4380 66342 4394 66394
rect 4394 66342 4406 66394
rect 4406 66342 4436 66394
rect 4460 66342 4470 66394
rect 4470 66342 4516 66394
rect 4220 66340 4276 66342
rect 4300 66340 4356 66342
rect 4380 66340 4436 66342
rect 4460 66340 4516 66342
rect 3974 65184 4030 65240
rect 3974 62600 4030 62656
rect 3974 60832 4030 60888
rect 3974 60716 4030 60752
rect 3974 60696 3976 60716
rect 3976 60696 4028 60716
rect 4028 60696 4030 60716
rect 3974 60560 4030 60616
rect 4220 65306 4276 65308
rect 4300 65306 4356 65308
rect 4380 65306 4436 65308
rect 4460 65306 4516 65308
rect 4220 65254 4266 65306
rect 4266 65254 4276 65306
rect 4300 65254 4330 65306
rect 4330 65254 4342 65306
rect 4342 65254 4356 65306
rect 4380 65254 4394 65306
rect 4394 65254 4406 65306
rect 4406 65254 4436 65306
rect 4460 65254 4470 65306
rect 4470 65254 4516 65306
rect 4220 65252 4276 65254
rect 4300 65252 4356 65254
rect 4380 65252 4436 65254
rect 4460 65252 4516 65254
rect 4220 64218 4276 64220
rect 4300 64218 4356 64220
rect 4380 64218 4436 64220
rect 4460 64218 4516 64220
rect 4220 64166 4266 64218
rect 4266 64166 4276 64218
rect 4300 64166 4330 64218
rect 4330 64166 4342 64218
rect 4342 64166 4356 64218
rect 4380 64166 4394 64218
rect 4394 64166 4406 64218
rect 4406 64166 4436 64218
rect 4460 64166 4470 64218
rect 4470 64166 4516 64218
rect 4220 64164 4276 64166
rect 4300 64164 4356 64166
rect 4380 64164 4436 64166
rect 4460 64164 4516 64166
rect 4220 63130 4276 63132
rect 4300 63130 4356 63132
rect 4380 63130 4436 63132
rect 4460 63130 4516 63132
rect 4220 63078 4266 63130
rect 4266 63078 4276 63130
rect 4300 63078 4330 63130
rect 4330 63078 4342 63130
rect 4342 63078 4356 63130
rect 4380 63078 4394 63130
rect 4394 63078 4406 63130
rect 4406 63078 4436 63130
rect 4460 63078 4470 63130
rect 4470 63078 4516 63130
rect 4220 63076 4276 63078
rect 4300 63076 4356 63078
rect 4380 63076 4436 63078
rect 4460 63076 4516 63078
rect 4220 62042 4276 62044
rect 4300 62042 4356 62044
rect 4380 62042 4436 62044
rect 4460 62042 4516 62044
rect 4220 61990 4266 62042
rect 4266 61990 4276 62042
rect 4300 61990 4330 62042
rect 4330 61990 4342 62042
rect 4342 61990 4356 62042
rect 4380 61990 4394 62042
rect 4394 61990 4406 62042
rect 4406 61990 4436 62042
rect 4460 61990 4470 62042
rect 4470 61990 4516 62042
rect 4220 61988 4276 61990
rect 4300 61988 4356 61990
rect 4380 61988 4436 61990
rect 4460 61988 4516 61990
rect 4220 60954 4276 60956
rect 4300 60954 4356 60956
rect 4380 60954 4436 60956
rect 4460 60954 4516 60956
rect 4220 60902 4266 60954
rect 4266 60902 4276 60954
rect 4300 60902 4330 60954
rect 4330 60902 4342 60954
rect 4342 60902 4356 60954
rect 4380 60902 4394 60954
rect 4394 60902 4406 60954
rect 4406 60902 4436 60954
rect 4460 60902 4470 60954
rect 4470 60902 4516 60954
rect 4220 60900 4276 60902
rect 4300 60900 4356 60902
rect 4380 60900 4436 60902
rect 4460 60900 4516 60902
rect 4220 59866 4276 59868
rect 4300 59866 4356 59868
rect 4380 59866 4436 59868
rect 4460 59866 4516 59868
rect 4220 59814 4266 59866
rect 4266 59814 4276 59866
rect 4300 59814 4330 59866
rect 4330 59814 4342 59866
rect 4342 59814 4356 59866
rect 4380 59814 4394 59866
rect 4394 59814 4406 59866
rect 4406 59814 4436 59866
rect 4460 59814 4470 59866
rect 4470 59814 4516 59866
rect 4220 59812 4276 59814
rect 4300 59812 4356 59814
rect 4380 59812 4436 59814
rect 4460 59812 4516 59814
rect 4220 58778 4276 58780
rect 4300 58778 4356 58780
rect 4380 58778 4436 58780
rect 4460 58778 4516 58780
rect 4220 58726 4266 58778
rect 4266 58726 4276 58778
rect 4300 58726 4330 58778
rect 4330 58726 4342 58778
rect 4342 58726 4356 58778
rect 4380 58726 4394 58778
rect 4394 58726 4406 58778
rect 4406 58726 4436 58778
rect 4460 58726 4470 58778
rect 4470 58726 4516 58778
rect 4220 58724 4276 58726
rect 4300 58724 4356 58726
rect 4380 58724 4436 58726
rect 4460 58724 4516 58726
rect 4220 57690 4276 57692
rect 4300 57690 4356 57692
rect 4380 57690 4436 57692
rect 4460 57690 4516 57692
rect 4220 57638 4266 57690
rect 4266 57638 4276 57690
rect 4300 57638 4330 57690
rect 4330 57638 4342 57690
rect 4342 57638 4356 57690
rect 4380 57638 4394 57690
rect 4394 57638 4406 57690
rect 4406 57638 4436 57690
rect 4460 57638 4470 57690
rect 4470 57638 4516 57690
rect 4220 57636 4276 57638
rect 4300 57636 4356 57638
rect 4380 57636 4436 57638
rect 4460 57636 4516 57638
rect 3974 55392 4030 55448
rect 4220 56602 4276 56604
rect 4300 56602 4356 56604
rect 4380 56602 4436 56604
rect 4460 56602 4516 56604
rect 4220 56550 4266 56602
rect 4266 56550 4276 56602
rect 4300 56550 4330 56602
rect 4330 56550 4342 56602
rect 4342 56550 4356 56602
rect 4380 56550 4394 56602
rect 4394 56550 4406 56602
rect 4406 56550 4436 56602
rect 4460 56550 4470 56602
rect 4470 56550 4516 56602
rect 4220 56548 4276 56550
rect 4300 56548 4356 56550
rect 4380 56548 4436 56550
rect 4460 56548 4516 56550
rect 7484 72922 7540 72924
rect 7564 72922 7620 72924
rect 7644 72922 7700 72924
rect 7724 72922 7780 72924
rect 7484 72870 7530 72922
rect 7530 72870 7540 72922
rect 7564 72870 7594 72922
rect 7594 72870 7606 72922
rect 7606 72870 7620 72922
rect 7644 72870 7658 72922
rect 7658 72870 7670 72922
rect 7670 72870 7700 72922
rect 7724 72870 7734 72922
rect 7734 72870 7780 72922
rect 7484 72868 7540 72870
rect 7564 72868 7620 72870
rect 7644 72868 7700 72870
rect 7724 72868 7780 72870
rect 5852 72378 5908 72380
rect 5932 72378 5988 72380
rect 6012 72378 6068 72380
rect 6092 72378 6148 72380
rect 5852 72326 5898 72378
rect 5898 72326 5908 72378
rect 5932 72326 5962 72378
rect 5962 72326 5974 72378
rect 5974 72326 5988 72378
rect 6012 72326 6026 72378
rect 6026 72326 6038 72378
rect 6038 72326 6068 72378
rect 6092 72326 6102 72378
rect 6102 72326 6148 72378
rect 5852 72324 5908 72326
rect 5932 72324 5988 72326
rect 6012 72324 6068 72326
rect 6092 72324 6148 72326
rect 7484 71834 7540 71836
rect 7564 71834 7620 71836
rect 7644 71834 7700 71836
rect 7724 71834 7780 71836
rect 7484 71782 7530 71834
rect 7530 71782 7540 71834
rect 7564 71782 7594 71834
rect 7594 71782 7606 71834
rect 7606 71782 7620 71834
rect 7644 71782 7658 71834
rect 7658 71782 7670 71834
rect 7670 71782 7700 71834
rect 7724 71782 7734 71834
rect 7734 71782 7780 71834
rect 7484 71780 7540 71782
rect 7564 71780 7620 71782
rect 7644 71780 7700 71782
rect 7724 71780 7780 71782
rect 9116 72378 9172 72380
rect 9196 72378 9252 72380
rect 9276 72378 9332 72380
rect 9356 72378 9412 72380
rect 9116 72326 9162 72378
rect 9162 72326 9172 72378
rect 9196 72326 9226 72378
rect 9226 72326 9238 72378
rect 9238 72326 9252 72378
rect 9276 72326 9290 72378
rect 9290 72326 9302 72378
rect 9302 72326 9332 72378
rect 9356 72326 9366 72378
rect 9366 72326 9412 72378
rect 9116 72324 9172 72326
rect 9196 72324 9252 72326
rect 9276 72324 9332 72326
rect 9356 72324 9412 72326
rect 5852 71290 5908 71292
rect 5932 71290 5988 71292
rect 6012 71290 6068 71292
rect 6092 71290 6148 71292
rect 5852 71238 5898 71290
rect 5898 71238 5908 71290
rect 5932 71238 5962 71290
rect 5962 71238 5974 71290
rect 5974 71238 5988 71290
rect 6012 71238 6026 71290
rect 6026 71238 6038 71290
rect 6038 71238 6068 71290
rect 6092 71238 6102 71290
rect 6102 71238 6148 71290
rect 5852 71236 5908 71238
rect 5932 71236 5988 71238
rect 6012 71236 6068 71238
rect 6092 71236 6148 71238
rect 9116 71290 9172 71292
rect 9196 71290 9252 71292
rect 9276 71290 9332 71292
rect 9356 71290 9412 71292
rect 9116 71238 9162 71290
rect 9162 71238 9172 71290
rect 9196 71238 9226 71290
rect 9226 71238 9238 71290
rect 9238 71238 9252 71290
rect 9276 71238 9290 71290
rect 9290 71238 9302 71290
rect 9302 71238 9332 71290
rect 9356 71238 9366 71290
rect 9366 71238 9412 71290
rect 9116 71236 9172 71238
rect 9196 71236 9252 71238
rect 9276 71236 9332 71238
rect 9356 71236 9412 71238
rect 7484 70746 7540 70748
rect 7564 70746 7620 70748
rect 7644 70746 7700 70748
rect 7724 70746 7780 70748
rect 7484 70694 7530 70746
rect 7530 70694 7540 70746
rect 7564 70694 7594 70746
rect 7594 70694 7606 70746
rect 7606 70694 7620 70746
rect 7644 70694 7658 70746
rect 7658 70694 7670 70746
rect 7670 70694 7700 70746
rect 7724 70694 7734 70746
rect 7734 70694 7780 70746
rect 7484 70692 7540 70694
rect 7564 70692 7620 70694
rect 7644 70692 7700 70694
rect 7724 70692 7780 70694
rect 5852 70202 5908 70204
rect 5932 70202 5988 70204
rect 6012 70202 6068 70204
rect 6092 70202 6148 70204
rect 5852 70150 5898 70202
rect 5898 70150 5908 70202
rect 5932 70150 5962 70202
rect 5962 70150 5974 70202
rect 5974 70150 5988 70202
rect 6012 70150 6026 70202
rect 6026 70150 6038 70202
rect 6038 70150 6068 70202
rect 6092 70150 6102 70202
rect 6102 70150 6148 70202
rect 5852 70148 5908 70150
rect 5932 70148 5988 70150
rect 6012 70148 6068 70150
rect 6092 70148 6148 70150
rect 9116 70202 9172 70204
rect 9196 70202 9252 70204
rect 9276 70202 9332 70204
rect 9356 70202 9412 70204
rect 9116 70150 9162 70202
rect 9162 70150 9172 70202
rect 9196 70150 9226 70202
rect 9226 70150 9238 70202
rect 9238 70150 9252 70202
rect 9276 70150 9290 70202
rect 9290 70150 9302 70202
rect 9302 70150 9332 70202
rect 9356 70150 9366 70202
rect 9366 70150 9412 70202
rect 9116 70148 9172 70150
rect 9196 70148 9252 70150
rect 9276 70148 9332 70150
rect 9356 70148 9412 70150
rect 7484 69658 7540 69660
rect 7564 69658 7620 69660
rect 7644 69658 7700 69660
rect 7724 69658 7780 69660
rect 7484 69606 7530 69658
rect 7530 69606 7540 69658
rect 7564 69606 7594 69658
rect 7594 69606 7606 69658
rect 7606 69606 7620 69658
rect 7644 69606 7658 69658
rect 7658 69606 7670 69658
rect 7670 69606 7700 69658
rect 7724 69606 7734 69658
rect 7734 69606 7780 69658
rect 7484 69604 7540 69606
rect 7564 69604 7620 69606
rect 7644 69604 7700 69606
rect 7724 69604 7780 69606
rect 5852 69114 5908 69116
rect 5932 69114 5988 69116
rect 6012 69114 6068 69116
rect 6092 69114 6148 69116
rect 5852 69062 5898 69114
rect 5898 69062 5908 69114
rect 5932 69062 5962 69114
rect 5962 69062 5974 69114
rect 5974 69062 5988 69114
rect 6012 69062 6026 69114
rect 6026 69062 6038 69114
rect 6038 69062 6068 69114
rect 6092 69062 6102 69114
rect 6102 69062 6148 69114
rect 5852 69060 5908 69062
rect 5932 69060 5988 69062
rect 6012 69060 6068 69062
rect 6092 69060 6148 69062
rect 9116 69114 9172 69116
rect 9196 69114 9252 69116
rect 9276 69114 9332 69116
rect 9356 69114 9412 69116
rect 9116 69062 9162 69114
rect 9162 69062 9172 69114
rect 9196 69062 9226 69114
rect 9226 69062 9238 69114
rect 9238 69062 9252 69114
rect 9276 69062 9290 69114
rect 9290 69062 9302 69114
rect 9302 69062 9332 69114
rect 9356 69062 9366 69114
rect 9366 69062 9412 69114
rect 9116 69060 9172 69062
rect 9196 69060 9252 69062
rect 9276 69060 9332 69062
rect 9356 69060 9412 69062
rect 4158 55800 4214 55856
rect 4618 55800 4674 55856
rect 4220 55514 4276 55516
rect 4300 55514 4356 55516
rect 4380 55514 4436 55516
rect 4460 55514 4516 55516
rect 4220 55462 4266 55514
rect 4266 55462 4276 55514
rect 4300 55462 4330 55514
rect 4330 55462 4342 55514
rect 4342 55462 4356 55514
rect 4380 55462 4394 55514
rect 4394 55462 4406 55514
rect 4406 55462 4436 55514
rect 4460 55462 4470 55514
rect 4470 55462 4516 55514
rect 4220 55460 4276 55462
rect 4300 55460 4356 55462
rect 4380 55460 4436 55462
rect 4460 55460 4516 55462
rect 4158 55276 4214 55312
rect 4158 55256 4160 55276
rect 4160 55256 4212 55276
rect 4212 55256 4214 55276
rect 4220 54426 4276 54428
rect 4300 54426 4356 54428
rect 4380 54426 4436 54428
rect 4460 54426 4516 54428
rect 4220 54374 4266 54426
rect 4266 54374 4276 54426
rect 4300 54374 4330 54426
rect 4330 54374 4342 54426
rect 4342 54374 4356 54426
rect 4380 54374 4394 54426
rect 4394 54374 4406 54426
rect 4406 54374 4436 54426
rect 4460 54374 4470 54426
rect 4470 54374 4516 54426
rect 4220 54372 4276 54374
rect 4300 54372 4356 54374
rect 4380 54372 4436 54374
rect 4460 54372 4516 54374
rect 4434 53624 4490 53680
rect 4526 53488 4582 53544
rect 4220 53338 4276 53340
rect 4300 53338 4356 53340
rect 4380 53338 4436 53340
rect 4460 53338 4516 53340
rect 4220 53286 4266 53338
rect 4266 53286 4276 53338
rect 4300 53286 4330 53338
rect 4330 53286 4342 53338
rect 4342 53286 4356 53338
rect 4380 53286 4394 53338
rect 4394 53286 4406 53338
rect 4406 53286 4436 53338
rect 4460 53286 4470 53338
rect 4470 53286 4516 53338
rect 4220 53284 4276 53286
rect 4300 53284 4356 53286
rect 4380 53284 4436 53286
rect 4460 53284 4516 53286
rect 4220 52250 4276 52252
rect 4300 52250 4356 52252
rect 4380 52250 4436 52252
rect 4460 52250 4516 52252
rect 4220 52198 4266 52250
rect 4266 52198 4276 52250
rect 4300 52198 4330 52250
rect 4330 52198 4342 52250
rect 4342 52198 4356 52250
rect 4380 52198 4394 52250
rect 4394 52198 4406 52250
rect 4406 52198 4436 52250
rect 4460 52198 4470 52250
rect 4470 52198 4516 52250
rect 4220 52196 4276 52198
rect 4300 52196 4356 52198
rect 4380 52196 4436 52198
rect 4460 52196 4516 52198
rect 4220 51162 4276 51164
rect 4300 51162 4356 51164
rect 4380 51162 4436 51164
rect 4460 51162 4516 51164
rect 4220 51110 4266 51162
rect 4266 51110 4276 51162
rect 4300 51110 4330 51162
rect 4330 51110 4342 51162
rect 4342 51110 4356 51162
rect 4380 51110 4394 51162
rect 4394 51110 4406 51162
rect 4406 51110 4436 51162
rect 4460 51110 4470 51162
rect 4470 51110 4516 51162
rect 4220 51108 4276 51110
rect 4300 51108 4356 51110
rect 4380 51108 4436 51110
rect 4460 51108 4516 51110
rect 3882 49408 3938 49464
rect 3422 46416 3478 46472
rect 3330 42200 3386 42256
rect 3054 32000 3110 32056
rect 3974 49172 3976 49192
rect 3976 49172 4028 49192
rect 4028 49172 4030 49192
rect 3974 49136 4030 49172
rect 3974 49036 3976 49056
rect 3976 49036 4028 49056
rect 4028 49036 4030 49056
rect 3974 49000 4030 49036
rect 3974 48864 4030 48920
rect 4250 50360 4306 50416
rect 4220 50074 4276 50076
rect 4300 50074 4356 50076
rect 4380 50074 4436 50076
rect 4460 50074 4516 50076
rect 4220 50022 4266 50074
rect 4266 50022 4276 50074
rect 4300 50022 4330 50074
rect 4330 50022 4342 50074
rect 4342 50022 4356 50074
rect 4380 50022 4394 50074
rect 4394 50022 4406 50074
rect 4406 50022 4436 50074
rect 4460 50022 4470 50074
rect 4470 50022 4516 50074
rect 4220 50020 4276 50022
rect 4300 50020 4356 50022
rect 4380 50020 4436 50022
rect 4460 50020 4516 50022
rect 4526 49136 4582 49192
rect 4220 48986 4276 48988
rect 4300 48986 4356 48988
rect 4380 48986 4436 48988
rect 4460 48986 4516 48988
rect 4220 48934 4266 48986
rect 4266 48934 4276 48986
rect 4300 48934 4330 48986
rect 4330 48934 4342 48986
rect 4342 48934 4356 48986
rect 4380 48934 4394 48986
rect 4394 48934 4406 48986
rect 4406 48934 4436 48986
rect 4460 48934 4470 48986
rect 4470 48934 4516 48986
rect 4220 48932 4276 48934
rect 4300 48932 4356 48934
rect 4380 48932 4436 48934
rect 4460 48932 4516 48934
rect 3974 48592 4030 48648
rect 3882 48320 3938 48376
rect 3790 48184 3846 48240
rect 3790 48048 3846 48104
rect 3790 45600 3846 45656
rect 3606 43016 3662 43072
rect 3606 41656 3662 41712
rect 3606 41112 3662 41168
rect 3514 32272 3570 32328
rect 3422 32136 3478 32192
rect 3330 31628 3332 31648
rect 3332 31628 3384 31648
rect 3384 31628 3386 31648
rect 3330 31592 3386 31628
rect 3330 31456 3386 31512
rect 2778 31320 2834 31376
rect 2588 31034 2644 31036
rect 2668 31034 2724 31036
rect 2748 31034 2804 31036
rect 2828 31034 2884 31036
rect 2588 30982 2634 31034
rect 2634 30982 2644 31034
rect 2668 30982 2698 31034
rect 2698 30982 2710 31034
rect 2710 30982 2724 31034
rect 2748 30982 2762 31034
rect 2762 30982 2774 31034
rect 2774 30982 2804 31034
rect 2828 30982 2838 31034
rect 2838 30982 2884 31034
rect 2588 30980 2644 30982
rect 2668 30980 2724 30982
rect 2748 30980 2804 30982
rect 2828 30980 2884 30982
rect 2962 30776 3018 30832
rect 2778 30368 2834 30424
rect 2594 30252 2650 30288
rect 2594 30232 2596 30252
rect 2596 30232 2648 30252
rect 2648 30232 2650 30252
rect 2588 29946 2644 29948
rect 2668 29946 2724 29948
rect 2748 29946 2804 29948
rect 2828 29946 2884 29948
rect 2588 29894 2634 29946
rect 2634 29894 2644 29946
rect 2668 29894 2698 29946
rect 2698 29894 2710 29946
rect 2710 29894 2724 29946
rect 2748 29894 2762 29946
rect 2762 29894 2774 29946
rect 2774 29894 2804 29946
rect 2828 29894 2838 29946
rect 2838 29894 2884 29946
rect 2588 29892 2644 29894
rect 2668 29892 2724 29894
rect 2748 29892 2804 29894
rect 2828 29892 2884 29894
rect 3146 30504 3202 30560
rect 3054 30368 3110 30424
rect 2588 28858 2644 28860
rect 2668 28858 2724 28860
rect 2748 28858 2804 28860
rect 2828 28858 2884 28860
rect 2588 28806 2634 28858
rect 2634 28806 2644 28858
rect 2668 28806 2698 28858
rect 2698 28806 2710 28858
rect 2710 28806 2724 28858
rect 2748 28806 2762 28858
rect 2762 28806 2774 28858
rect 2774 28806 2804 28858
rect 2828 28806 2838 28858
rect 2838 28806 2884 28858
rect 2588 28804 2644 28806
rect 2668 28804 2724 28806
rect 2748 28804 2804 28806
rect 2828 28804 2884 28806
rect 2134 28464 2190 28520
rect 2226 28328 2282 28384
rect 2134 28192 2190 28248
rect 1950 28056 2006 28112
rect 1950 27920 2006 27976
rect 1858 23976 1914 24032
rect 1398 18808 1454 18864
rect 1582 16632 1638 16688
rect 1398 14592 1454 14648
rect 1490 12416 1546 12472
rect 1582 12008 1638 12064
rect 1398 10784 1454 10840
rect 1490 10376 1546 10432
rect 1398 9832 1454 9888
rect 1490 9424 1546 9480
rect 1398 9016 1454 9072
rect 1398 8608 1454 8664
rect 1398 8200 1454 8256
rect 1398 7828 1400 7848
rect 1400 7828 1452 7848
rect 1452 7828 1454 7848
rect 1398 7792 1454 7828
rect 1306 5616 1362 5672
rect 1398 5208 1454 5264
rect 1490 3984 1546 4040
rect 1398 3576 1454 3632
rect 2410 24112 2466 24168
rect 2594 28600 2650 28656
rect 2588 27770 2644 27772
rect 2668 27770 2724 27772
rect 2748 27770 2804 27772
rect 2828 27770 2884 27772
rect 2588 27718 2634 27770
rect 2634 27718 2644 27770
rect 2668 27718 2698 27770
rect 2698 27718 2710 27770
rect 2710 27718 2724 27770
rect 2748 27718 2762 27770
rect 2762 27718 2774 27770
rect 2774 27718 2804 27770
rect 2828 27718 2838 27770
rect 2838 27718 2884 27770
rect 2588 27716 2644 27718
rect 2668 27716 2724 27718
rect 2748 27716 2804 27718
rect 2828 27716 2884 27718
rect 3054 27956 3056 27976
rect 3056 27956 3108 27976
rect 3108 27956 3110 27976
rect 3054 27920 3110 27956
rect 2870 26968 2926 27024
rect 2588 26682 2644 26684
rect 2668 26682 2724 26684
rect 2748 26682 2804 26684
rect 2828 26682 2884 26684
rect 2588 26630 2634 26682
rect 2634 26630 2644 26682
rect 2668 26630 2698 26682
rect 2698 26630 2710 26682
rect 2710 26630 2724 26682
rect 2748 26630 2762 26682
rect 2762 26630 2774 26682
rect 2774 26630 2804 26682
rect 2828 26630 2838 26682
rect 2838 26630 2884 26682
rect 2588 26628 2644 26630
rect 2668 26628 2724 26630
rect 2748 26628 2804 26630
rect 2828 26628 2884 26630
rect 3054 26424 3110 26480
rect 3146 26288 3202 26344
rect 2594 26016 2650 26072
rect 2588 25594 2644 25596
rect 2668 25594 2724 25596
rect 2748 25594 2804 25596
rect 2828 25594 2884 25596
rect 2588 25542 2634 25594
rect 2634 25542 2644 25594
rect 2668 25542 2698 25594
rect 2698 25542 2710 25594
rect 2710 25542 2724 25594
rect 2748 25542 2762 25594
rect 2762 25542 2774 25594
rect 2774 25542 2804 25594
rect 2828 25542 2838 25594
rect 2838 25542 2884 25594
rect 2588 25540 2644 25542
rect 2668 25540 2724 25542
rect 2748 25540 2804 25542
rect 2828 25540 2884 25542
rect 2962 25200 3018 25256
rect 2870 24656 2926 24712
rect 2588 24506 2644 24508
rect 2668 24506 2724 24508
rect 2748 24506 2804 24508
rect 2828 24506 2884 24508
rect 2588 24454 2634 24506
rect 2634 24454 2644 24506
rect 2668 24454 2698 24506
rect 2698 24454 2710 24506
rect 2710 24454 2724 24506
rect 2748 24454 2762 24506
rect 2762 24454 2774 24506
rect 2774 24454 2804 24506
rect 2828 24454 2838 24506
rect 2838 24454 2884 24506
rect 2588 24452 2644 24454
rect 2668 24452 2724 24454
rect 2748 24452 2804 24454
rect 2828 24452 2884 24454
rect 2588 23418 2644 23420
rect 2668 23418 2724 23420
rect 2748 23418 2804 23420
rect 2828 23418 2884 23420
rect 2588 23366 2634 23418
rect 2634 23366 2644 23418
rect 2668 23366 2698 23418
rect 2698 23366 2710 23418
rect 2710 23366 2724 23418
rect 2748 23366 2762 23418
rect 2762 23366 2774 23418
rect 2774 23366 2804 23418
rect 2828 23366 2838 23418
rect 2838 23366 2884 23418
rect 2588 23364 2644 23366
rect 2668 23364 2724 23366
rect 2748 23364 2804 23366
rect 2828 23364 2884 23366
rect 2588 22330 2644 22332
rect 2668 22330 2724 22332
rect 2748 22330 2804 22332
rect 2828 22330 2884 22332
rect 2588 22278 2634 22330
rect 2634 22278 2644 22330
rect 2668 22278 2698 22330
rect 2698 22278 2710 22330
rect 2710 22278 2724 22330
rect 2748 22278 2762 22330
rect 2762 22278 2774 22330
rect 2774 22278 2804 22330
rect 2828 22278 2838 22330
rect 2838 22278 2884 22330
rect 2588 22276 2644 22278
rect 2668 22276 2724 22278
rect 2748 22276 2804 22278
rect 2828 22276 2884 22278
rect 2588 21242 2644 21244
rect 2668 21242 2724 21244
rect 2748 21242 2804 21244
rect 2828 21242 2884 21244
rect 2588 21190 2634 21242
rect 2634 21190 2644 21242
rect 2668 21190 2698 21242
rect 2698 21190 2710 21242
rect 2710 21190 2724 21242
rect 2748 21190 2762 21242
rect 2762 21190 2774 21242
rect 2774 21190 2804 21242
rect 2828 21190 2838 21242
rect 2838 21190 2884 21242
rect 2588 21188 2644 21190
rect 2668 21188 2724 21190
rect 2748 21188 2804 21190
rect 2828 21188 2884 21190
rect 3330 27376 3386 27432
rect 3330 25744 3386 25800
rect 2778 20576 2834 20632
rect 2588 20154 2644 20156
rect 2668 20154 2724 20156
rect 2748 20154 2804 20156
rect 2828 20154 2884 20156
rect 2588 20102 2634 20154
rect 2634 20102 2644 20154
rect 2668 20102 2698 20154
rect 2698 20102 2710 20154
rect 2710 20102 2724 20154
rect 2748 20102 2762 20154
rect 2762 20102 2774 20154
rect 2774 20102 2804 20154
rect 2828 20102 2838 20154
rect 2838 20102 2884 20154
rect 2588 20100 2644 20102
rect 2668 20100 2724 20102
rect 2748 20100 2804 20102
rect 2828 20100 2884 20102
rect 2588 19066 2644 19068
rect 2668 19066 2724 19068
rect 2748 19066 2804 19068
rect 2828 19066 2884 19068
rect 2588 19014 2634 19066
rect 2634 19014 2644 19066
rect 2668 19014 2698 19066
rect 2698 19014 2710 19066
rect 2710 19014 2724 19066
rect 2748 19014 2762 19066
rect 2762 19014 2774 19066
rect 2774 19014 2804 19066
rect 2828 19014 2838 19066
rect 2838 19014 2884 19066
rect 2588 19012 2644 19014
rect 2668 19012 2724 19014
rect 2748 19012 2804 19014
rect 2828 19012 2884 19014
rect 2226 15408 2282 15464
rect 2588 17978 2644 17980
rect 2668 17978 2724 17980
rect 2748 17978 2804 17980
rect 2828 17978 2884 17980
rect 2588 17926 2634 17978
rect 2634 17926 2644 17978
rect 2668 17926 2698 17978
rect 2698 17926 2710 17978
rect 2710 17926 2724 17978
rect 2748 17926 2762 17978
rect 2762 17926 2774 17978
rect 2774 17926 2804 17978
rect 2828 17926 2838 17978
rect 2838 17926 2884 17978
rect 2588 17924 2644 17926
rect 2668 17924 2724 17926
rect 2748 17924 2804 17926
rect 2828 17924 2884 17926
rect 2410 17176 2466 17232
rect 3054 17584 3110 17640
rect 2588 16890 2644 16892
rect 2668 16890 2724 16892
rect 2748 16890 2804 16892
rect 2828 16890 2884 16892
rect 2588 16838 2634 16890
rect 2634 16838 2644 16890
rect 2668 16838 2698 16890
rect 2698 16838 2710 16890
rect 2710 16838 2724 16890
rect 2748 16838 2762 16890
rect 2762 16838 2774 16890
rect 2774 16838 2804 16890
rect 2828 16838 2838 16890
rect 2838 16838 2884 16890
rect 2588 16836 2644 16838
rect 2668 16836 2724 16838
rect 2748 16836 2804 16838
rect 2828 16836 2884 16838
rect 2870 15952 2926 16008
rect 2588 15802 2644 15804
rect 2668 15802 2724 15804
rect 2748 15802 2804 15804
rect 2828 15802 2884 15804
rect 2588 15750 2634 15802
rect 2634 15750 2644 15802
rect 2668 15750 2698 15802
rect 2698 15750 2710 15802
rect 2710 15750 2724 15802
rect 2748 15750 2762 15802
rect 2762 15750 2774 15802
rect 2774 15750 2804 15802
rect 2828 15750 2838 15802
rect 2838 15750 2884 15802
rect 2588 15748 2644 15750
rect 2668 15748 2724 15750
rect 2748 15748 2804 15750
rect 2828 15748 2884 15750
rect 2588 14714 2644 14716
rect 2668 14714 2724 14716
rect 2748 14714 2804 14716
rect 2828 14714 2884 14716
rect 2588 14662 2634 14714
rect 2634 14662 2644 14714
rect 2668 14662 2698 14714
rect 2698 14662 2710 14714
rect 2710 14662 2724 14714
rect 2748 14662 2762 14714
rect 2762 14662 2774 14714
rect 2774 14662 2804 14714
rect 2828 14662 2838 14714
rect 2838 14662 2884 14714
rect 2588 14660 2644 14662
rect 2668 14660 2724 14662
rect 2748 14660 2804 14662
rect 2828 14660 2884 14662
rect 2962 13776 3018 13832
rect 2588 13626 2644 13628
rect 2668 13626 2724 13628
rect 2748 13626 2804 13628
rect 2828 13626 2884 13628
rect 2588 13574 2634 13626
rect 2634 13574 2644 13626
rect 2668 13574 2698 13626
rect 2698 13574 2710 13626
rect 2710 13574 2724 13626
rect 2748 13574 2762 13626
rect 2762 13574 2774 13626
rect 2774 13574 2804 13626
rect 2828 13574 2838 13626
rect 2838 13574 2884 13626
rect 2588 13572 2644 13574
rect 2668 13572 2724 13574
rect 2748 13572 2804 13574
rect 2828 13572 2884 13574
rect 2588 12538 2644 12540
rect 2668 12538 2724 12540
rect 2748 12538 2804 12540
rect 2828 12538 2884 12540
rect 2588 12486 2634 12538
rect 2634 12486 2644 12538
rect 2668 12486 2698 12538
rect 2698 12486 2710 12538
rect 2710 12486 2724 12538
rect 2748 12486 2762 12538
rect 2762 12486 2774 12538
rect 2774 12486 2804 12538
rect 2828 12486 2838 12538
rect 2838 12486 2884 12538
rect 2588 12484 2644 12486
rect 2668 12484 2724 12486
rect 2748 12484 2804 12486
rect 2828 12484 2884 12486
rect 3238 17076 3240 17096
rect 3240 17076 3292 17096
rect 3292 17076 3294 17096
rect 3238 17040 3294 17076
rect 3698 40976 3754 41032
rect 3698 38392 3754 38448
rect 3974 46960 4030 47016
rect 4220 47898 4276 47900
rect 4300 47898 4356 47900
rect 4380 47898 4436 47900
rect 4460 47898 4516 47900
rect 4220 47846 4266 47898
rect 4266 47846 4276 47898
rect 4300 47846 4330 47898
rect 4330 47846 4342 47898
rect 4342 47846 4356 47898
rect 4380 47846 4394 47898
rect 4394 47846 4406 47898
rect 4406 47846 4436 47898
rect 4460 47846 4470 47898
rect 4470 47846 4516 47898
rect 4220 47844 4276 47846
rect 4300 47844 4356 47846
rect 4380 47844 4436 47846
rect 4460 47844 4516 47846
rect 4250 46980 4306 47016
rect 4250 46960 4252 46980
rect 4252 46960 4304 46980
rect 4304 46960 4306 46980
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4266 46810
rect 4266 46758 4276 46810
rect 4300 46758 4330 46810
rect 4330 46758 4342 46810
rect 4342 46758 4356 46810
rect 4380 46758 4394 46810
rect 4394 46758 4406 46810
rect 4406 46758 4436 46810
rect 4460 46758 4470 46810
rect 4470 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 3974 45600 4030 45656
rect 3974 43596 3976 43616
rect 3976 43596 4028 43616
rect 4028 43596 4030 43616
rect 3974 43560 4030 43596
rect 3974 43172 4030 43208
rect 3974 43152 3976 43172
rect 3976 43152 4028 43172
rect 4028 43152 4030 43172
rect 3974 42608 4030 42664
rect 3790 36216 3846 36272
rect 3974 40160 4030 40216
rect 3974 39480 4030 39536
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4266 45722
rect 4266 45670 4276 45722
rect 4300 45670 4330 45722
rect 4330 45670 4342 45722
rect 4342 45670 4356 45722
rect 4380 45670 4394 45722
rect 4394 45670 4406 45722
rect 4406 45670 4436 45722
rect 4460 45670 4470 45722
rect 4470 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4158 44784 4214 44840
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4266 44634
rect 4266 44582 4276 44634
rect 4300 44582 4330 44634
rect 4330 44582 4342 44634
rect 4342 44582 4356 44634
rect 4380 44582 4394 44634
rect 4394 44582 4406 44634
rect 4406 44582 4436 44634
rect 4460 44582 4470 44634
rect 4470 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4266 43546
rect 4266 43494 4276 43546
rect 4300 43494 4330 43546
rect 4330 43494 4342 43546
rect 4342 43494 4356 43546
rect 4380 43494 4394 43546
rect 4394 43494 4406 43546
rect 4406 43494 4436 43546
rect 4460 43494 4470 43546
rect 4470 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4158 43288 4214 43344
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4266 42458
rect 4266 42406 4276 42458
rect 4300 42406 4330 42458
rect 4330 42406 4342 42458
rect 4342 42406 4356 42458
rect 4380 42406 4394 42458
rect 4394 42406 4406 42458
rect 4406 42406 4436 42458
rect 4460 42406 4470 42458
rect 4470 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4434 41520 4490 41576
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4266 41370
rect 4266 41318 4276 41370
rect 4300 41318 4330 41370
rect 4330 41318 4342 41370
rect 4342 41318 4356 41370
rect 4380 41318 4394 41370
rect 4394 41318 4406 41370
rect 4406 41318 4436 41370
rect 4460 41318 4470 41370
rect 4470 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4266 40282
rect 4266 40230 4276 40282
rect 4300 40230 4330 40282
rect 4330 40230 4342 40282
rect 4342 40230 4356 40282
rect 4380 40230 4394 40282
rect 4394 40230 4406 40282
rect 4406 40230 4436 40282
rect 4460 40230 4470 40282
rect 4470 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 3974 39244 3976 39264
rect 3976 39244 4028 39264
rect 4028 39244 4030 39264
rect 3974 39208 4030 39244
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4266 39194
rect 4266 39142 4276 39194
rect 4300 39142 4330 39194
rect 4330 39142 4342 39194
rect 4342 39142 4356 39194
rect 4380 39142 4394 39194
rect 4394 39142 4406 39194
rect 4406 39142 4436 39194
rect 4460 39142 4470 39194
rect 4470 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4802 55800 4858 55856
rect 4158 38936 4214 38992
rect 3974 38800 4030 38856
rect 3974 37712 4030 37768
rect 3974 37168 4030 37224
rect 7484 68570 7540 68572
rect 7564 68570 7620 68572
rect 7644 68570 7700 68572
rect 7724 68570 7780 68572
rect 7484 68518 7530 68570
rect 7530 68518 7540 68570
rect 7564 68518 7594 68570
rect 7594 68518 7606 68570
rect 7606 68518 7620 68570
rect 7644 68518 7658 68570
rect 7658 68518 7670 68570
rect 7670 68518 7700 68570
rect 7724 68518 7734 68570
rect 7734 68518 7780 68570
rect 7484 68516 7540 68518
rect 7564 68516 7620 68518
rect 7644 68516 7700 68518
rect 7724 68516 7780 68518
rect 5852 68026 5908 68028
rect 5932 68026 5988 68028
rect 6012 68026 6068 68028
rect 6092 68026 6148 68028
rect 5852 67974 5898 68026
rect 5898 67974 5908 68026
rect 5932 67974 5962 68026
rect 5962 67974 5974 68026
rect 5974 67974 5988 68026
rect 6012 67974 6026 68026
rect 6026 67974 6038 68026
rect 6038 67974 6068 68026
rect 6092 67974 6102 68026
rect 6102 67974 6148 68026
rect 5852 67972 5908 67974
rect 5932 67972 5988 67974
rect 6012 67972 6068 67974
rect 6092 67972 6148 67974
rect 9116 68026 9172 68028
rect 9196 68026 9252 68028
rect 9276 68026 9332 68028
rect 9356 68026 9412 68028
rect 9116 67974 9162 68026
rect 9162 67974 9172 68026
rect 9196 67974 9226 68026
rect 9226 67974 9238 68026
rect 9238 67974 9252 68026
rect 9276 67974 9290 68026
rect 9290 67974 9302 68026
rect 9302 67974 9332 68026
rect 9356 67974 9366 68026
rect 9366 67974 9412 68026
rect 9116 67972 9172 67974
rect 9196 67972 9252 67974
rect 9276 67972 9332 67974
rect 9356 67972 9412 67974
rect 7484 67482 7540 67484
rect 7564 67482 7620 67484
rect 7644 67482 7700 67484
rect 7724 67482 7780 67484
rect 7484 67430 7530 67482
rect 7530 67430 7540 67482
rect 7564 67430 7594 67482
rect 7594 67430 7606 67482
rect 7606 67430 7620 67482
rect 7644 67430 7658 67482
rect 7658 67430 7670 67482
rect 7670 67430 7700 67482
rect 7724 67430 7734 67482
rect 7734 67430 7780 67482
rect 7484 67428 7540 67430
rect 7564 67428 7620 67430
rect 7644 67428 7700 67430
rect 7724 67428 7780 67430
rect 5852 66938 5908 66940
rect 5932 66938 5988 66940
rect 6012 66938 6068 66940
rect 6092 66938 6148 66940
rect 5852 66886 5898 66938
rect 5898 66886 5908 66938
rect 5932 66886 5962 66938
rect 5962 66886 5974 66938
rect 5974 66886 5988 66938
rect 6012 66886 6026 66938
rect 6026 66886 6038 66938
rect 6038 66886 6068 66938
rect 6092 66886 6102 66938
rect 6102 66886 6148 66938
rect 5852 66884 5908 66886
rect 5932 66884 5988 66886
rect 6012 66884 6068 66886
rect 6092 66884 6148 66886
rect 7484 66394 7540 66396
rect 7564 66394 7620 66396
rect 7644 66394 7700 66396
rect 7724 66394 7780 66396
rect 7484 66342 7530 66394
rect 7530 66342 7540 66394
rect 7564 66342 7594 66394
rect 7594 66342 7606 66394
rect 7606 66342 7620 66394
rect 7644 66342 7658 66394
rect 7658 66342 7670 66394
rect 7670 66342 7700 66394
rect 7724 66342 7734 66394
rect 7734 66342 7780 66394
rect 7484 66340 7540 66342
rect 7564 66340 7620 66342
rect 7644 66340 7700 66342
rect 7724 66340 7780 66342
rect 5852 65850 5908 65852
rect 5932 65850 5988 65852
rect 6012 65850 6068 65852
rect 6092 65850 6148 65852
rect 5852 65798 5898 65850
rect 5898 65798 5908 65850
rect 5932 65798 5962 65850
rect 5962 65798 5974 65850
rect 5974 65798 5988 65850
rect 6012 65798 6026 65850
rect 6026 65798 6038 65850
rect 6038 65798 6068 65850
rect 6092 65798 6102 65850
rect 6102 65798 6148 65850
rect 5852 65796 5908 65798
rect 5932 65796 5988 65798
rect 6012 65796 6068 65798
rect 6092 65796 6148 65798
rect 7484 65306 7540 65308
rect 7564 65306 7620 65308
rect 7644 65306 7700 65308
rect 7724 65306 7780 65308
rect 7484 65254 7530 65306
rect 7530 65254 7540 65306
rect 7564 65254 7594 65306
rect 7594 65254 7606 65306
rect 7606 65254 7620 65306
rect 7644 65254 7658 65306
rect 7658 65254 7670 65306
rect 7670 65254 7700 65306
rect 7724 65254 7734 65306
rect 7734 65254 7780 65306
rect 7484 65252 7540 65254
rect 7564 65252 7620 65254
rect 7644 65252 7700 65254
rect 7724 65252 7780 65254
rect 5852 64762 5908 64764
rect 5932 64762 5988 64764
rect 6012 64762 6068 64764
rect 6092 64762 6148 64764
rect 5852 64710 5898 64762
rect 5898 64710 5908 64762
rect 5932 64710 5962 64762
rect 5962 64710 5974 64762
rect 5974 64710 5988 64762
rect 6012 64710 6026 64762
rect 6026 64710 6038 64762
rect 6038 64710 6068 64762
rect 6092 64710 6102 64762
rect 6102 64710 6148 64762
rect 5852 64708 5908 64710
rect 5932 64708 5988 64710
rect 6012 64708 6068 64710
rect 6092 64708 6148 64710
rect 7484 64218 7540 64220
rect 7564 64218 7620 64220
rect 7644 64218 7700 64220
rect 7724 64218 7780 64220
rect 7484 64166 7530 64218
rect 7530 64166 7540 64218
rect 7564 64166 7594 64218
rect 7594 64166 7606 64218
rect 7606 64166 7620 64218
rect 7644 64166 7658 64218
rect 7658 64166 7670 64218
rect 7670 64166 7700 64218
rect 7724 64166 7734 64218
rect 7734 64166 7780 64218
rect 7484 64164 7540 64166
rect 7564 64164 7620 64166
rect 7644 64164 7700 64166
rect 7724 64164 7780 64166
rect 5078 53080 5134 53136
rect 5078 51176 5134 51232
rect 5078 51040 5134 51096
rect 5852 63674 5908 63676
rect 5932 63674 5988 63676
rect 6012 63674 6068 63676
rect 6092 63674 6148 63676
rect 5852 63622 5898 63674
rect 5898 63622 5908 63674
rect 5932 63622 5962 63674
rect 5962 63622 5974 63674
rect 5974 63622 5988 63674
rect 6012 63622 6026 63674
rect 6026 63622 6038 63674
rect 6038 63622 6068 63674
rect 6092 63622 6102 63674
rect 6102 63622 6148 63674
rect 5852 63620 5908 63622
rect 5932 63620 5988 63622
rect 6012 63620 6068 63622
rect 6092 63620 6148 63622
rect 7484 63130 7540 63132
rect 7564 63130 7620 63132
rect 7644 63130 7700 63132
rect 7724 63130 7780 63132
rect 7484 63078 7530 63130
rect 7530 63078 7540 63130
rect 7564 63078 7594 63130
rect 7594 63078 7606 63130
rect 7606 63078 7620 63130
rect 7644 63078 7658 63130
rect 7658 63078 7670 63130
rect 7670 63078 7700 63130
rect 7724 63078 7734 63130
rect 7734 63078 7780 63130
rect 7484 63076 7540 63078
rect 7564 63076 7620 63078
rect 7644 63076 7700 63078
rect 7724 63076 7780 63078
rect 4986 50224 5042 50280
rect 4802 42064 4858 42120
rect 4342 38256 4398 38312
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4266 38106
rect 4266 38054 4276 38106
rect 4300 38054 4330 38106
rect 4330 38054 4342 38106
rect 4342 38054 4356 38106
rect 4380 38054 4394 38106
rect 4394 38054 4406 38106
rect 4406 38054 4436 38106
rect 4460 38054 4470 38106
rect 4470 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4266 37018
rect 4266 36966 4276 37018
rect 4300 36966 4330 37018
rect 4330 36966 4342 37018
rect 4342 36966 4356 37018
rect 4380 36966 4394 37018
rect 4394 36966 4406 37018
rect 4406 36966 4436 37018
rect 4460 36966 4470 37018
rect 4470 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 3974 36624 4030 36680
rect 3698 35808 3754 35864
rect 3698 32816 3754 32872
rect 3606 31204 3662 31240
rect 3606 31184 3608 31204
rect 3608 31184 3660 31204
rect 3660 31184 3662 31204
rect 3606 30640 3662 30696
rect 3606 25744 3662 25800
rect 3514 22480 3570 22536
rect 4158 36080 4214 36136
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4266 35930
rect 4266 35878 4276 35930
rect 4300 35878 4330 35930
rect 4330 35878 4342 35930
rect 4342 35878 4356 35930
rect 4380 35878 4394 35930
rect 4394 35878 4406 35930
rect 4406 35878 4436 35930
rect 4460 35878 4470 35930
rect 4470 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 3974 35808 4030 35864
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4266 34842
rect 4266 34790 4276 34842
rect 4300 34790 4330 34842
rect 4330 34790 4342 34842
rect 4342 34790 4356 34842
rect 4380 34790 4394 34842
rect 4394 34790 4406 34842
rect 4406 34790 4436 34842
rect 4460 34790 4470 34842
rect 4470 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 3974 32408 4030 32464
rect 3974 31864 4030 31920
rect 3882 31728 3938 31784
rect 3882 31456 3938 31512
rect 3974 30912 4030 30968
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4266 33754
rect 4266 33702 4276 33754
rect 4300 33702 4330 33754
rect 4330 33702 4342 33754
rect 4342 33702 4356 33754
rect 4380 33702 4394 33754
rect 4394 33702 4406 33754
rect 4406 33702 4436 33754
rect 4460 33702 4470 33754
rect 4470 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4526 32952 4582 33008
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4266 32666
rect 4266 32614 4276 32666
rect 4300 32614 4330 32666
rect 4330 32614 4342 32666
rect 4342 32614 4356 32666
rect 4380 32614 4394 32666
rect 4394 32614 4406 32666
rect 4406 32614 4436 32666
rect 4460 32614 4470 32666
rect 4470 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4526 32408 4582 32464
rect 4710 32000 4766 32056
rect 5852 62586 5908 62588
rect 5932 62586 5988 62588
rect 6012 62586 6068 62588
rect 6092 62586 6148 62588
rect 5852 62534 5898 62586
rect 5898 62534 5908 62586
rect 5932 62534 5962 62586
rect 5962 62534 5974 62586
rect 5974 62534 5988 62586
rect 6012 62534 6026 62586
rect 6026 62534 6038 62586
rect 6038 62534 6068 62586
rect 6092 62534 6102 62586
rect 6102 62534 6148 62586
rect 5852 62532 5908 62534
rect 5932 62532 5988 62534
rect 6012 62532 6068 62534
rect 6092 62532 6148 62534
rect 7484 62042 7540 62044
rect 7564 62042 7620 62044
rect 7644 62042 7700 62044
rect 7724 62042 7780 62044
rect 7484 61990 7530 62042
rect 7530 61990 7540 62042
rect 7564 61990 7594 62042
rect 7594 61990 7606 62042
rect 7606 61990 7620 62042
rect 7644 61990 7658 62042
rect 7658 61990 7670 62042
rect 7670 61990 7700 62042
rect 7724 61990 7734 62042
rect 7734 61990 7780 62042
rect 7484 61988 7540 61990
rect 7564 61988 7620 61990
rect 7644 61988 7700 61990
rect 7724 61988 7780 61990
rect 5852 61498 5908 61500
rect 5932 61498 5988 61500
rect 6012 61498 6068 61500
rect 6092 61498 6148 61500
rect 5852 61446 5898 61498
rect 5898 61446 5908 61498
rect 5932 61446 5962 61498
rect 5962 61446 5974 61498
rect 5974 61446 5988 61498
rect 6012 61446 6026 61498
rect 6026 61446 6038 61498
rect 6038 61446 6068 61498
rect 6092 61446 6102 61498
rect 6102 61446 6148 61498
rect 5852 61444 5908 61446
rect 5932 61444 5988 61446
rect 6012 61444 6068 61446
rect 6092 61444 6148 61446
rect 7484 60954 7540 60956
rect 7564 60954 7620 60956
rect 7644 60954 7700 60956
rect 7724 60954 7780 60956
rect 7484 60902 7530 60954
rect 7530 60902 7540 60954
rect 7564 60902 7594 60954
rect 7594 60902 7606 60954
rect 7606 60902 7620 60954
rect 7644 60902 7658 60954
rect 7658 60902 7670 60954
rect 7670 60902 7700 60954
rect 7724 60902 7734 60954
rect 7734 60902 7780 60954
rect 7484 60900 7540 60902
rect 7564 60900 7620 60902
rect 7644 60900 7700 60902
rect 7724 60900 7780 60902
rect 5852 60410 5908 60412
rect 5932 60410 5988 60412
rect 6012 60410 6068 60412
rect 6092 60410 6148 60412
rect 5852 60358 5898 60410
rect 5898 60358 5908 60410
rect 5932 60358 5962 60410
rect 5962 60358 5974 60410
rect 5974 60358 5988 60410
rect 6012 60358 6026 60410
rect 6026 60358 6038 60410
rect 6038 60358 6068 60410
rect 6092 60358 6102 60410
rect 6102 60358 6148 60410
rect 5852 60356 5908 60358
rect 5932 60356 5988 60358
rect 6012 60356 6068 60358
rect 6092 60356 6148 60358
rect 5852 59322 5908 59324
rect 5932 59322 5988 59324
rect 6012 59322 6068 59324
rect 6092 59322 6148 59324
rect 5852 59270 5898 59322
rect 5898 59270 5908 59322
rect 5932 59270 5962 59322
rect 5962 59270 5974 59322
rect 5974 59270 5988 59322
rect 6012 59270 6026 59322
rect 6026 59270 6038 59322
rect 6038 59270 6068 59322
rect 6092 59270 6102 59322
rect 6102 59270 6148 59322
rect 5852 59268 5908 59270
rect 5932 59268 5988 59270
rect 6012 59268 6068 59270
rect 6092 59268 6148 59270
rect 5852 58234 5908 58236
rect 5932 58234 5988 58236
rect 6012 58234 6068 58236
rect 6092 58234 6148 58236
rect 5852 58182 5898 58234
rect 5898 58182 5908 58234
rect 5932 58182 5962 58234
rect 5962 58182 5974 58234
rect 5974 58182 5988 58234
rect 6012 58182 6026 58234
rect 6026 58182 6038 58234
rect 6038 58182 6068 58234
rect 6092 58182 6102 58234
rect 6102 58182 6148 58234
rect 5852 58180 5908 58182
rect 5932 58180 5988 58182
rect 6012 58180 6068 58182
rect 6092 58180 6148 58182
rect 7484 59866 7540 59868
rect 7564 59866 7620 59868
rect 7644 59866 7700 59868
rect 7724 59866 7780 59868
rect 7484 59814 7530 59866
rect 7530 59814 7540 59866
rect 7564 59814 7594 59866
rect 7594 59814 7606 59866
rect 7606 59814 7620 59866
rect 7644 59814 7658 59866
rect 7658 59814 7670 59866
rect 7670 59814 7700 59866
rect 7724 59814 7734 59866
rect 7734 59814 7780 59866
rect 7484 59812 7540 59814
rect 7564 59812 7620 59814
rect 7644 59812 7700 59814
rect 7724 59812 7780 59814
rect 7484 58778 7540 58780
rect 7564 58778 7620 58780
rect 7644 58778 7700 58780
rect 7724 58778 7780 58780
rect 7484 58726 7530 58778
rect 7530 58726 7540 58778
rect 7564 58726 7594 58778
rect 7594 58726 7606 58778
rect 7606 58726 7620 58778
rect 7644 58726 7658 58778
rect 7658 58726 7670 58778
rect 7670 58726 7700 58778
rect 7724 58726 7734 58778
rect 7734 58726 7780 58778
rect 7484 58724 7540 58726
rect 7564 58724 7620 58726
rect 7644 58724 7700 58726
rect 7724 58724 7780 58726
rect 7484 57690 7540 57692
rect 7564 57690 7620 57692
rect 7644 57690 7700 57692
rect 7724 57690 7780 57692
rect 7484 57638 7530 57690
rect 7530 57638 7540 57690
rect 7564 57638 7594 57690
rect 7594 57638 7606 57690
rect 7606 57638 7620 57690
rect 7644 57638 7658 57690
rect 7658 57638 7670 57690
rect 7670 57638 7700 57690
rect 7724 57638 7734 57690
rect 7734 57638 7780 57690
rect 7484 57636 7540 57638
rect 7564 57636 7620 57638
rect 7644 57636 7700 57638
rect 7724 57636 7780 57638
rect 6918 57432 6974 57488
rect 5852 57146 5908 57148
rect 5932 57146 5988 57148
rect 6012 57146 6068 57148
rect 6092 57146 6148 57148
rect 5852 57094 5898 57146
rect 5898 57094 5908 57146
rect 5932 57094 5962 57146
rect 5962 57094 5974 57146
rect 5974 57094 5988 57146
rect 6012 57094 6026 57146
rect 6026 57094 6038 57146
rect 6038 57094 6068 57146
rect 6092 57094 6102 57146
rect 6102 57094 6148 57146
rect 5852 57092 5908 57094
rect 5932 57092 5988 57094
rect 6012 57092 6068 57094
rect 6092 57092 6148 57094
rect 5852 56058 5908 56060
rect 5932 56058 5988 56060
rect 6012 56058 6068 56060
rect 6092 56058 6148 56060
rect 5852 56006 5898 56058
rect 5898 56006 5908 56058
rect 5932 56006 5962 56058
rect 5962 56006 5974 56058
rect 5974 56006 5988 56058
rect 6012 56006 6026 56058
rect 6026 56006 6038 56058
rect 6038 56006 6068 56058
rect 6092 56006 6102 56058
rect 6102 56006 6148 56058
rect 5852 56004 5908 56006
rect 5932 56004 5988 56006
rect 6012 56004 6068 56006
rect 6092 56004 6148 56006
rect 5722 55664 5778 55720
rect 5446 51040 5502 51096
rect 5170 50904 5226 50960
rect 5078 41520 5134 41576
rect 4986 36216 5042 36272
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4266 31578
rect 4266 31526 4276 31578
rect 4300 31526 4330 31578
rect 4330 31526 4342 31578
rect 4342 31526 4356 31578
rect 4380 31526 4394 31578
rect 4394 31526 4406 31578
rect 4406 31526 4436 31578
rect 4460 31526 4470 31578
rect 4470 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4158 31320 4214 31376
rect 3882 24792 3938 24848
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4266 30490
rect 4266 30438 4276 30490
rect 4300 30438 4330 30490
rect 4330 30438 4342 30490
rect 4342 30438 4356 30490
rect 4380 30438 4394 30490
rect 4394 30438 4406 30490
rect 4406 30438 4436 30490
rect 4460 30438 4470 30490
rect 4470 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4266 29402
rect 4266 29350 4276 29402
rect 4300 29350 4330 29402
rect 4330 29350 4342 29402
rect 4342 29350 4356 29402
rect 4380 29350 4394 29402
rect 4394 29350 4406 29402
rect 4406 29350 4436 29402
rect 4460 29350 4470 29402
rect 4470 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4066 29044 4068 29064
rect 4068 29044 4120 29064
rect 4120 29044 4122 29064
rect 4066 29008 4122 29044
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4266 28314
rect 4266 28262 4276 28314
rect 4300 28262 4330 28314
rect 4330 28262 4342 28314
rect 4342 28262 4356 28314
rect 4380 28262 4394 28314
rect 4394 28262 4406 28314
rect 4406 28262 4436 28314
rect 4460 28262 4470 28314
rect 4470 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4266 27226
rect 4266 27174 4276 27226
rect 4300 27174 4330 27226
rect 4330 27174 4342 27226
rect 4342 27174 4356 27226
rect 4380 27174 4394 27226
rect 4394 27174 4406 27226
rect 4406 27174 4436 27226
rect 4460 27174 4470 27226
rect 4470 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4526 27004 4528 27024
rect 4528 27004 4580 27024
rect 4580 27004 4582 27024
rect 4526 26968 4582 27004
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4266 26138
rect 4266 26086 4276 26138
rect 4300 26086 4330 26138
rect 4330 26086 4342 26138
rect 4342 26086 4356 26138
rect 4380 26086 4394 26138
rect 4394 26086 4406 26138
rect 4406 26086 4436 26138
rect 4460 26086 4470 26138
rect 4470 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4266 25050
rect 4266 24998 4276 25050
rect 4300 24998 4330 25050
rect 4330 24998 4342 25050
rect 4342 24998 4356 25050
rect 4380 24998 4394 25050
rect 4394 24998 4406 25050
rect 4406 24998 4436 25050
rect 4460 24998 4470 25050
rect 4470 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4266 23962
rect 4266 23910 4276 23962
rect 4300 23910 4330 23962
rect 4330 23910 4342 23962
rect 4342 23910 4356 23962
rect 4380 23910 4394 23962
rect 4394 23910 4406 23962
rect 4406 23910 4436 23962
rect 4460 23910 4470 23962
rect 4470 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 3882 22616 3938 22672
rect 3698 18128 3754 18184
rect 3422 15680 3478 15736
rect 3422 13232 3478 13288
rect 3606 14048 3662 14104
rect 3514 12960 3570 13016
rect 3054 11756 3110 11792
rect 3054 11736 3056 11756
rect 3056 11736 3108 11756
rect 3108 11736 3110 11756
rect 2962 11464 3018 11520
rect 2588 11450 2644 11452
rect 2668 11450 2724 11452
rect 2748 11450 2804 11452
rect 2828 11450 2884 11452
rect 2588 11398 2634 11450
rect 2634 11398 2644 11450
rect 2668 11398 2698 11450
rect 2698 11398 2710 11450
rect 2710 11398 2724 11450
rect 2748 11398 2762 11450
rect 2762 11398 2774 11450
rect 2774 11398 2804 11450
rect 2828 11398 2838 11450
rect 2838 11398 2884 11450
rect 2588 11396 2644 11398
rect 2668 11396 2724 11398
rect 2748 11396 2804 11398
rect 2828 11396 2884 11398
rect 2588 10362 2644 10364
rect 2668 10362 2724 10364
rect 2748 10362 2804 10364
rect 2828 10362 2884 10364
rect 2588 10310 2634 10362
rect 2634 10310 2644 10362
rect 2668 10310 2698 10362
rect 2698 10310 2710 10362
rect 2710 10310 2724 10362
rect 2748 10310 2762 10362
rect 2762 10310 2774 10362
rect 2774 10310 2804 10362
rect 2828 10310 2838 10362
rect 2838 10310 2884 10362
rect 2588 10308 2644 10310
rect 2668 10308 2724 10310
rect 2748 10308 2804 10310
rect 2828 10308 2884 10310
rect 2588 9274 2644 9276
rect 2668 9274 2724 9276
rect 2748 9274 2804 9276
rect 2828 9274 2884 9276
rect 2588 9222 2634 9274
rect 2634 9222 2644 9274
rect 2668 9222 2698 9274
rect 2698 9222 2710 9274
rect 2710 9222 2724 9274
rect 2748 9222 2762 9274
rect 2762 9222 2774 9274
rect 2774 9222 2804 9274
rect 2828 9222 2838 9274
rect 2838 9222 2884 9274
rect 2588 9220 2644 9222
rect 2668 9220 2724 9222
rect 2748 9220 2804 9222
rect 2828 9220 2884 9222
rect 3422 12416 3478 12472
rect 2588 8186 2644 8188
rect 2668 8186 2724 8188
rect 2748 8186 2804 8188
rect 2828 8186 2884 8188
rect 2588 8134 2634 8186
rect 2634 8134 2644 8186
rect 2668 8134 2698 8186
rect 2698 8134 2710 8186
rect 2710 8134 2724 8186
rect 2748 8134 2762 8186
rect 2762 8134 2774 8186
rect 2774 8134 2804 8186
rect 2828 8134 2838 8186
rect 2838 8134 2884 8186
rect 2588 8132 2644 8134
rect 2668 8132 2724 8134
rect 2748 8132 2804 8134
rect 2828 8132 2884 8134
rect 2962 7384 3018 7440
rect 1582 3032 1638 3088
rect 2588 7098 2644 7100
rect 2668 7098 2724 7100
rect 2748 7098 2804 7100
rect 2828 7098 2884 7100
rect 2588 7046 2634 7098
rect 2634 7046 2644 7098
rect 2668 7046 2698 7098
rect 2698 7046 2710 7098
rect 2710 7046 2724 7098
rect 2748 7046 2762 7098
rect 2762 7046 2774 7098
rect 2774 7046 2804 7098
rect 2828 7046 2838 7098
rect 2838 7046 2884 7098
rect 2588 7044 2644 7046
rect 2668 7044 2724 7046
rect 2748 7044 2804 7046
rect 2828 7044 2884 7046
rect 2594 6704 2650 6760
rect 3146 6432 3202 6488
rect 2962 6160 3018 6216
rect 2588 6010 2644 6012
rect 2668 6010 2724 6012
rect 2748 6010 2804 6012
rect 2828 6010 2884 6012
rect 2588 5958 2634 6010
rect 2634 5958 2644 6010
rect 2668 5958 2698 6010
rect 2698 5958 2710 6010
rect 2710 5958 2724 6010
rect 2748 5958 2762 6010
rect 2762 5958 2774 6010
rect 2774 5958 2804 6010
rect 2828 5958 2838 6010
rect 2838 5958 2884 6010
rect 2588 5956 2644 5958
rect 2668 5956 2724 5958
rect 2748 5956 2804 5958
rect 2828 5956 2884 5958
rect 2962 5908 3018 5944
rect 2962 5888 2964 5908
rect 2964 5888 3016 5908
rect 3016 5888 3018 5908
rect 2870 5208 2926 5264
rect 2588 4922 2644 4924
rect 2668 4922 2724 4924
rect 2748 4922 2804 4924
rect 2828 4922 2884 4924
rect 2588 4870 2634 4922
rect 2634 4870 2644 4922
rect 2668 4870 2698 4922
rect 2698 4870 2710 4922
rect 2710 4870 2724 4922
rect 2748 4870 2762 4922
rect 2762 4870 2774 4922
rect 2774 4870 2804 4922
rect 2828 4870 2838 4922
rect 2838 4870 2884 4922
rect 2588 4868 2644 4870
rect 2668 4868 2724 4870
rect 2748 4868 2804 4870
rect 2828 4868 2884 4870
rect 2588 3834 2644 3836
rect 2668 3834 2724 3836
rect 2748 3834 2804 3836
rect 2828 3834 2884 3836
rect 2588 3782 2634 3834
rect 2634 3782 2644 3834
rect 2668 3782 2698 3834
rect 2698 3782 2710 3834
rect 2710 3782 2724 3834
rect 2748 3782 2762 3834
rect 2762 3782 2774 3834
rect 2774 3782 2804 3834
rect 2828 3782 2838 3834
rect 2838 3782 2884 3834
rect 2588 3780 2644 3782
rect 2668 3780 2724 3782
rect 2748 3780 2804 3782
rect 2828 3780 2884 3782
rect 3974 18400 4030 18456
rect 3974 16224 4030 16280
rect 3974 14184 4030 14240
rect 3882 13368 3938 13424
rect 3698 11600 3754 11656
rect 3606 7248 3662 7304
rect 3974 12824 4030 12880
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4266 22874
rect 4266 22822 4276 22874
rect 4300 22822 4330 22874
rect 4330 22822 4342 22874
rect 4342 22822 4356 22874
rect 4380 22822 4394 22874
rect 4394 22822 4406 22874
rect 4406 22822 4436 22874
rect 4460 22822 4470 22874
rect 4470 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4266 21786
rect 4266 21734 4276 21786
rect 4300 21734 4330 21786
rect 4330 21734 4342 21786
rect 4342 21734 4356 21786
rect 4380 21734 4394 21786
rect 4394 21734 4406 21786
rect 4406 21734 4436 21786
rect 4460 21734 4470 21786
rect 4470 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4266 20698
rect 4266 20646 4276 20698
rect 4300 20646 4330 20698
rect 4330 20646 4342 20698
rect 4342 20646 4356 20698
rect 4380 20646 4394 20698
rect 4394 20646 4406 20698
rect 4406 20646 4436 20698
rect 4460 20646 4470 20698
rect 4470 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4266 19610
rect 4266 19558 4276 19610
rect 4300 19558 4330 19610
rect 4330 19558 4342 19610
rect 4342 19558 4356 19610
rect 4380 19558 4394 19610
rect 4394 19558 4406 19610
rect 4406 19558 4436 19610
rect 4460 19558 4470 19610
rect 4470 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4266 18522
rect 4266 18470 4276 18522
rect 4300 18470 4330 18522
rect 4330 18470 4342 18522
rect 4342 18470 4356 18522
rect 4380 18470 4394 18522
rect 4394 18470 4406 18522
rect 4406 18470 4436 18522
rect 4460 18470 4470 18522
rect 4470 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4266 17434
rect 4266 17382 4276 17434
rect 4300 17382 4330 17434
rect 4330 17382 4342 17434
rect 4342 17382 4356 17434
rect 4380 17382 4394 17434
rect 4394 17382 4406 17434
rect 4406 17382 4436 17434
rect 4460 17382 4470 17434
rect 4470 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4986 31728 5042 31784
rect 4894 22888 4950 22944
rect 4894 22616 4950 22672
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4266 16346
rect 4266 16294 4276 16346
rect 4300 16294 4330 16346
rect 4330 16294 4342 16346
rect 4342 16294 4356 16346
rect 4380 16294 4394 16346
rect 4394 16294 4406 16346
rect 4406 16294 4436 16346
rect 4460 16294 4470 16346
rect 4470 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4266 15258
rect 4266 15206 4276 15258
rect 4300 15206 4330 15258
rect 4330 15206 4342 15258
rect 4342 15206 4356 15258
rect 4380 15206 4394 15258
rect 4394 15206 4406 15258
rect 4406 15206 4436 15258
rect 4460 15206 4470 15258
rect 4470 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4266 14170
rect 4266 14118 4276 14170
rect 4300 14118 4330 14170
rect 4330 14118 4342 14170
rect 4342 14118 4356 14170
rect 4380 14118 4394 14170
rect 4394 14118 4406 14170
rect 4406 14118 4436 14170
rect 4460 14118 4470 14170
rect 4470 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4266 13082
rect 4266 13030 4276 13082
rect 4300 13030 4330 13082
rect 4330 13030 4342 13082
rect 4342 13030 4356 13082
rect 4380 13030 4394 13082
rect 4394 13030 4406 13082
rect 4406 13030 4436 13082
rect 4460 13030 4470 13082
rect 4470 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4266 11994
rect 4266 11942 4276 11994
rect 4300 11942 4330 11994
rect 4330 11942 4342 11994
rect 4342 11942 4356 11994
rect 4380 11942 4394 11994
rect 4394 11942 4406 11994
rect 4406 11942 4436 11994
rect 4460 11942 4470 11994
rect 4470 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4266 10906
rect 4266 10854 4276 10906
rect 4300 10854 4330 10906
rect 4330 10854 4342 10906
rect 4342 10854 4356 10906
rect 4380 10854 4394 10906
rect 4394 10854 4406 10906
rect 4406 10854 4436 10906
rect 4460 10854 4470 10906
rect 4470 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 3974 10260 4030 10296
rect 3974 10240 3976 10260
rect 3976 10240 4028 10260
rect 4028 10240 4030 10260
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4266 9818
rect 4266 9766 4276 9818
rect 4300 9766 4330 9818
rect 4330 9766 4342 9818
rect 4342 9766 4356 9818
rect 4380 9766 4394 9818
rect 4394 9766 4406 9818
rect 4406 9766 4436 9818
rect 4460 9766 4470 9818
rect 4470 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4266 8730
rect 4266 8678 4276 8730
rect 4300 8678 4330 8730
rect 4330 8678 4342 8730
rect 4342 8678 4356 8730
rect 4380 8678 4394 8730
rect 4394 8678 4406 8730
rect 4406 8678 4436 8730
rect 4460 8678 4470 8730
rect 4470 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4266 7642
rect 4266 7590 4276 7642
rect 4300 7590 4330 7642
rect 4330 7590 4342 7642
rect 4342 7590 4356 7642
rect 4380 7590 4394 7642
rect 4394 7590 4406 7642
rect 4406 7590 4436 7642
rect 4460 7590 4470 7642
rect 4470 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 5630 51040 5686 51096
rect 5538 50904 5594 50960
rect 5354 50768 5410 50824
rect 5262 50632 5318 50688
rect 5354 45600 5410 45656
rect 5354 44920 5410 44976
rect 5630 41928 5686 41984
rect 5354 41384 5410 41440
rect 5852 54970 5908 54972
rect 5932 54970 5988 54972
rect 6012 54970 6068 54972
rect 6092 54970 6148 54972
rect 5852 54918 5898 54970
rect 5898 54918 5908 54970
rect 5932 54918 5962 54970
rect 5962 54918 5974 54970
rect 5974 54918 5988 54970
rect 6012 54918 6026 54970
rect 6026 54918 6038 54970
rect 6038 54918 6068 54970
rect 6092 54918 6102 54970
rect 6102 54918 6148 54970
rect 5852 54916 5908 54918
rect 5932 54916 5988 54918
rect 6012 54916 6068 54918
rect 6092 54916 6148 54918
rect 5852 53882 5908 53884
rect 5932 53882 5988 53884
rect 6012 53882 6068 53884
rect 6092 53882 6148 53884
rect 5852 53830 5898 53882
rect 5898 53830 5908 53882
rect 5932 53830 5962 53882
rect 5962 53830 5974 53882
rect 5974 53830 5988 53882
rect 6012 53830 6026 53882
rect 6026 53830 6038 53882
rect 6038 53830 6068 53882
rect 6092 53830 6102 53882
rect 6102 53830 6148 53882
rect 5852 53828 5908 53830
rect 5932 53828 5988 53830
rect 6012 53828 6068 53830
rect 6092 53828 6148 53830
rect 5852 52794 5908 52796
rect 5932 52794 5988 52796
rect 6012 52794 6068 52796
rect 6092 52794 6148 52796
rect 5852 52742 5898 52794
rect 5898 52742 5908 52794
rect 5932 52742 5962 52794
rect 5962 52742 5974 52794
rect 5974 52742 5988 52794
rect 6012 52742 6026 52794
rect 6026 52742 6038 52794
rect 6038 52742 6068 52794
rect 6092 52742 6102 52794
rect 6102 52742 6148 52794
rect 5852 52740 5908 52742
rect 5932 52740 5988 52742
rect 6012 52740 6068 52742
rect 6092 52740 6148 52742
rect 5852 51706 5908 51708
rect 5932 51706 5988 51708
rect 6012 51706 6068 51708
rect 6092 51706 6148 51708
rect 5852 51654 5898 51706
rect 5898 51654 5908 51706
rect 5932 51654 5962 51706
rect 5962 51654 5974 51706
rect 5974 51654 5988 51706
rect 6012 51654 6026 51706
rect 6026 51654 6038 51706
rect 6038 51654 6068 51706
rect 6092 51654 6102 51706
rect 6102 51654 6148 51706
rect 5852 51652 5908 51654
rect 5932 51652 5988 51654
rect 6012 51652 6068 51654
rect 6092 51652 6148 51654
rect 5852 50618 5908 50620
rect 5932 50618 5988 50620
rect 6012 50618 6068 50620
rect 6092 50618 6148 50620
rect 5852 50566 5898 50618
rect 5898 50566 5908 50618
rect 5932 50566 5962 50618
rect 5962 50566 5974 50618
rect 5974 50566 5988 50618
rect 6012 50566 6026 50618
rect 6026 50566 6038 50618
rect 6038 50566 6068 50618
rect 6092 50566 6102 50618
rect 6102 50566 6148 50618
rect 5852 50564 5908 50566
rect 5932 50564 5988 50566
rect 6012 50564 6068 50566
rect 6092 50564 6148 50566
rect 5852 49530 5908 49532
rect 5932 49530 5988 49532
rect 6012 49530 6068 49532
rect 6092 49530 6148 49532
rect 5852 49478 5898 49530
rect 5898 49478 5908 49530
rect 5932 49478 5962 49530
rect 5962 49478 5974 49530
rect 5974 49478 5988 49530
rect 6012 49478 6026 49530
rect 6026 49478 6038 49530
rect 6038 49478 6068 49530
rect 6092 49478 6102 49530
rect 6102 49478 6148 49530
rect 5852 49476 5908 49478
rect 5932 49476 5988 49478
rect 6012 49476 6068 49478
rect 6092 49476 6148 49478
rect 5852 48442 5908 48444
rect 5932 48442 5988 48444
rect 6012 48442 6068 48444
rect 6092 48442 6148 48444
rect 5852 48390 5898 48442
rect 5898 48390 5908 48442
rect 5932 48390 5962 48442
rect 5962 48390 5974 48442
rect 5974 48390 5988 48442
rect 6012 48390 6026 48442
rect 6026 48390 6038 48442
rect 6038 48390 6068 48442
rect 6092 48390 6102 48442
rect 6102 48390 6148 48442
rect 5852 48388 5908 48390
rect 5932 48388 5988 48390
rect 6012 48388 6068 48390
rect 6092 48388 6148 48390
rect 5852 47354 5908 47356
rect 5932 47354 5988 47356
rect 6012 47354 6068 47356
rect 6092 47354 6148 47356
rect 5852 47302 5898 47354
rect 5898 47302 5908 47354
rect 5932 47302 5962 47354
rect 5962 47302 5974 47354
rect 5974 47302 5988 47354
rect 6012 47302 6026 47354
rect 6026 47302 6038 47354
rect 6038 47302 6068 47354
rect 6092 47302 6102 47354
rect 6102 47302 6148 47354
rect 5852 47300 5908 47302
rect 5932 47300 5988 47302
rect 6012 47300 6068 47302
rect 6092 47300 6148 47302
rect 5852 46266 5908 46268
rect 5932 46266 5988 46268
rect 6012 46266 6068 46268
rect 6092 46266 6148 46268
rect 5852 46214 5898 46266
rect 5898 46214 5908 46266
rect 5932 46214 5962 46266
rect 5962 46214 5974 46266
rect 5974 46214 5988 46266
rect 6012 46214 6026 46266
rect 6026 46214 6038 46266
rect 6038 46214 6068 46266
rect 6092 46214 6102 46266
rect 6102 46214 6148 46266
rect 5852 46212 5908 46214
rect 5932 46212 5988 46214
rect 6012 46212 6068 46214
rect 6092 46212 6148 46214
rect 5852 45178 5908 45180
rect 5932 45178 5988 45180
rect 6012 45178 6068 45180
rect 6092 45178 6148 45180
rect 5852 45126 5898 45178
rect 5898 45126 5908 45178
rect 5932 45126 5962 45178
rect 5962 45126 5974 45178
rect 5974 45126 5988 45178
rect 6012 45126 6026 45178
rect 6026 45126 6038 45178
rect 6038 45126 6068 45178
rect 6092 45126 6102 45178
rect 6102 45126 6148 45178
rect 5852 45124 5908 45126
rect 5932 45124 5988 45126
rect 6012 45124 6068 45126
rect 6092 45124 6148 45126
rect 5852 44090 5908 44092
rect 5932 44090 5988 44092
rect 6012 44090 6068 44092
rect 6092 44090 6148 44092
rect 5852 44038 5898 44090
rect 5898 44038 5908 44090
rect 5932 44038 5962 44090
rect 5962 44038 5974 44090
rect 5974 44038 5988 44090
rect 6012 44038 6026 44090
rect 6026 44038 6038 44090
rect 6038 44038 6068 44090
rect 6092 44038 6102 44090
rect 6102 44038 6148 44090
rect 5852 44036 5908 44038
rect 5932 44036 5988 44038
rect 6012 44036 6068 44038
rect 6092 44036 6148 44038
rect 5852 43002 5908 43004
rect 5932 43002 5988 43004
rect 6012 43002 6068 43004
rect 6092 43002 6148 43004
rect 5852 42950 5898 43002
rect 5898 42950 5908 43002
rect 5932 42950 5962 43002
rect 5962 42950 5974 43002
rect 5974 42950 5988 43002
rect 6012 42950 6026 43002
rect 6026 42950 6038 43002
rect 6038 42950 6068 43002
rect 6092 42950 6102 43002
rect 6102 42950 6148 43002
rect 5852 42948 5908 42950
rect 5932 42948 5988 42950
rect 6012 42948 6068 42950
rect 6092 42948 6148 42950
rect 5852 41914 5908 41916
rect 5932 41914 5988 41916
rect 6012 41914 6068 41916
rect 6092 41914 6148 41916
rect 5852 41862 5898 41914
rect 5898 41862 5908 41914
rect 5932 41862 5962 41914
rect 5962 41862 5974 41914
rect 5974 41862 5988 41914
rect 6012 41862 6026 41914
rect 6026 41862 6038 41914
rect 6038 41862 6068 41914
rect 6092 41862 6102 41914
rect 6102 41862 6148 41914
rect 5852 41860 5908 41862
rect 5932 41860 5988 41862
rect 6012 41860 6068 41862
rect 6092 41860 6148 41862
rect 5354 36896 5410 36952
rect 5354 36624 5410 36680
rect 5262 31592 5318 31648
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4266 6554
rect 4266 6502 4276 6554
rect 4300 6502 4330 6554
rect 4330 6502 4342 6554
rect 4342 6502 4356 6554
rect 4380 6502 4394 6554
rect 4394 6502 4406 6554
rect 4406 6502 4436 6554
rect 4460 6502 4470 6554
rect 4470 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 3606 4392 3662 4448
rect 2588 2746 2644 2748
rect 2668 2746 2724 2748
rect 2748 2746 2804 2748
rect 2828 2746 2884 2748
rect 2588 2694 2634 2746
rect 2634 2694 2644 2746
rect 2668 2694 2698 2746
rect 2698 2694 2710 2746
rect 2710 2694 2724 2746
rect 2748 2694 2762 2746
rect 2762 2694 2774 2746
rect 2774 2694 2804 2746
rect 2828 2694 2838 2746
rect 2838 2694 2884 2746
rect 2588 2692 2644 2694
rect 2668 2692 2724 2694
rect 2748 2692 2804 2694
rect 2828 2692 2884 2694
rect 2226 1808 2282 1864
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4266 5466
rect 4266 5414 4276 5466
rect 4300 5414 4330 5466
rect 4330 5414 4342 5466
rect 4342 5414 4356 5466
rect 4380 5414 4394 5466
rect 4394 5414 4406 5466
rect 4406 5414 4436 5466
rect 4460 5414 4470 5466
rect 4470 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 5852 40826 5908 40828
rect 5932 40826 5988 40828
rect 6012 40826 6068 40828
rect 6092 40826 6148 40828
rect 5852 40774 5898 40826
rect 5898 40774 5908 40826
rect 5932 40774 5962 40826
rect 5962 40774 5974 40826
rect 5974 40774 5988 40826
rect 6012 40774 6026 40826
rect 6026 40774 6038 40826
rect 6038 40774 6068 40826
rect 6092 40774 6102 40826
rect 6102 40774 6148 40826
rect 5852 40772 5908 40774
rect 5932 40772 5988 40774
rect 6012 40772 6068 40774
rect 6092 40772 6148 40774
rect 5852 39738 5908 39740
rect 5932 39738 5988 39740
rect 6012 39738 6068 39740
rect 6092 39738 6148 39740
rect 5852 39686 5898 39738
rect 5898 39686 5908 39738
rect 5932 39686 5962 39738
rect 5962 39686 5974 39738
rect 5974 39686 5988 39738
rect 6012 39686 6026 39738
rect 6026 39686 6038 39738
rect 6038 39686 6068 39738
rect 6092 39686 6102 39738
rect 6102 39686 6148 39738
rect 5852 39684 5908 39686
rect 5932 39684 5988 39686
rect 6012 39684 6068 39686
rect 6092 39684 6148 39686
rect 5852 38650 5908 38652
rect 5932 38650 5988 38652
rect 6012 38650 6068 38652
rect 6092 38650 6148 38652
rect 5852 38598 5898 38650
rect 5898 38598 5908 38650
rect 5932 38598 5962 38650
rect 5962 38598 5974 38650
rect 5974 38598 5988 38650
rect 6012 38598 6026 38650
rect 6026 38598 6038 38650
rect 6038 38598 6068 38650
rect 6092 38598 6102 38650
rect 6102 38598 6148 38650
rect 5852 38596 5908 38598
rect 5932 38596 5988 38598
rect 6012 38596 6068 38598
rect 6092 38596 6148 38598
rect 5538 36352 5594 36408
rect 5852 37562 5908 37564
rect 5932 37562 5988 37564
rect 6012 37562 6068 37564
rect 6092 37562 6148 37564
rect 5852 37510 5898 37562
rect 5898 37510 5908 37562
rect 5932 37510 5962 37562
rect 5962 37510 5974 37562
rect 5974 37510 5988 37562
rect 6012 37510 6026 37562
rect 6026 37510 6038 37562
rect 6038 37510 6068 37562
rect 6092 37510 6102 37562
rect 6102 37510 6148 37562
rect 5852 37508 5908 37510
rect 5932 37508 5988 37510
rect 6012 37508 6068 37510
rect 6092 37508 6148 37510
rect 5852 36474 5908 36476
rect 5932 36474 5988 36476
rect 6012 36474 6068 36476
rect 6092 36474 6148 36476
rect 5852 36422 5898 36474
rect 5898 36422 5908 36474
rect 5932 36422 5962 36474
rect 5962 36422 5974 36474
rect 5974 36422 5988 36474
rect 6012 36422 6026 36474
rect 6026 36422 6038 36474
rect 6038 36422 6068 36474
rect 6092 36422 6102 36474
rect 6102 36422 6148 36474
rect 5852 36420 5908 36422
rect 5932 36420 5988 36422
rect 6012 36420 6068 36422
rect 6092 36420 6148 36422
rect 5852 35386 5908 35388
rect 5932 35386 5988 35388
rect 6012 35386 6068 35388
rect 6092 35386 6148 35388
rect 5852 35334 5898 35386
rect 5898 35334 5908 35386
rect 5932 35334 5962 35386
rect 5962 35334 5974 35386
rect 5974 35334 5988 35386
rect 6012 35334 6026 35386
rect 6026 35334 6038 35386
rect 6038 35334 6068 35386
rect 6092 35334 6102 35386
rect 6102 35334 6148 35386
rect 5852 35332 5908 35334
rect 5932 35332 5988 35334
rect 6012 35332 6068 35334
rect 6092 35332 6148 35334
rect 5852 34298 5908 34300
rect 5932 34298 5988 34300
rect 6012 34298 6068 34300
rect 6092 34298 6148 34300
rect 5852 34246 5898 34298
rect 5898 34246 5908 34298
rect 5932 34246 5962 34298
rect 5962 34246 5974 34298
rect 5974 34246 5988 34298
rect 6012 34246 6026 34298
rect 6026 34246 6038 34298
rect 6038 34246 6068 34298
rect 6092 34246 6102 34298
rect 6102 34246 6148 34298
rect 5852 34244 5908 34246
rect 5932 34244 5988 34246
rect 6012 34244 6068 34246
rect 6092 34244 6148 34246
rect 5852 33210 5908 33212
rect 5932 33210 5988 33212
rect 6012 33210 6068 33212
rect 6092 33210 6148 33212
rect 5852 33158 5898 33210
rect 5898 33158 5908 33210
rect 5932 33158 5962 33210
rect 5962 33158 5974 33210
rect 5974 33158 5988 33210
rect 6012 33158 6026 33210
rect 6026 33158 6038 33210
rect 6038 33158 6068 33210
rect 6092 33158 6102 33210
rect 6102 33158 6148 33210
rect 5852 33156 5908 33158
rect 5932 33156 5988 33158
rect 6012 33156 6068 33158
rect 6092 33156 6148 33158
rect 5852 32122 5908 32124
rect 5932 32122 5988 32124
rect 6012 32122 6068 32124
rect 6092 32122 6148 32124
rect 5852 32070 5898 32122
rect 5898 32070 5908 32122
rect 5932 32070 5962 32122
rect 5962 32070 5974 32122
rect 5974 32070 5988 32122
rect 6012 32070 6026 32122
rect 6026 32070 6038 32122
rect 6038 32070 6068 32122
rect 6092 32070 6102 32122
rect 6102 32070 6148 32122
rect 5852 32068 5908 32070
rect 5932 32068 5988 32070
rect 6012 32068 6068 32070
rect 6092 32068 6148 32070
rect 7484 56602 7540 56604
rect 7564 56602 7620 56604
rect 7644 56602 7700 56604
rect 7724 56602 7780 56604
rect 7484 56550 7530 56602
rect 7530 56550 7540 56602
rect 7564 56550 7594 56602
rect 7594 56550 7606 56602
rect 7606 56550 7620 56602
rect 7644 56550 7658 56602
rect 7658 56550 7670 56602
rect 7670 56550 7700 56602
rect 7724 56550 7734 56602
rect 7734 56550 7780 56602
rect 7484 56548 7540 56550
rect 7564 56548 7620 56550
rect 7644 56548 7700 56550
rect 7724 56548 7780 56550
rect 7484 55514 7540 55516
rect 7564 55514 7620 55516
rect 7644 55514 7700 55516
rect 7724 55514 7780 55516
rect 7484 55462 7530 55514
rect 7530 55462 7540 55514
rect 7564 55462 7594 55514
rect 7594 55462 7606 55514
rect 7606 55462 7620 55514
rect 7644 55462 7658 55514
rect 7658 55462 7670 55514
rect 7670 55462 7700 55514
rect 7724 55462 7734 55514
rect 7734 55462 7780 55514
rect 7484 55460 7540 55462
rect 7564 55460 7620 55462
rect 7644 55460 7700 55462
rect 7724 55460 7780 55462
rect 9116 66938 9172 66940
rect 9196 66938 9252 66940
rect 9276 66938 9332 66940
rect 9356 66938 9412 66940
rect 9116 66886 9162 66938
rect 9162 66886 9172 66938
rect 9196 66886 9226 66938
rect 9226 66886 9238 66938
rect 9238 66886 9252 66938
rect 9276 66886 9290 66938
rect 9290 66886 9302 66938
rect 9302 66886 9332 66938
rect 9356 66886 9366 66938
rect 9366 66886 9412 66938
rect 9116 66884 9172 66886
rect 9196 66884 9252 66886
rect 9276 66884 9332 66886
rect 9356 66884 9412 66886
rect 9116 65850 9172 65852
rect 9196 65850 9252 65852
rect 9276 65850 9332 65852
rect 9356 65850 9412 65852
rect 9116 65798 9162 65850
rect 9162 65798 9172 65850
rect 9196 65798 9226 65850
rect 9226 65798 9238 65850
rect 9238 65798 9252 65850
rect 9276 65798 9290 65850
rect 9290 65798 9302 65850
rect 9302 65798 9332 65850
rect 9356 65798 9366 65850
rect 9366 65798 9412 65850
rect 9116 65796 9172 65798
rect 9196 65796 9252 65798
rect 9276 65796 9332 65798
rect 9356 65796 9412 65798
rect 9116 64762 9172 64764
rect 9196 64762 9252 64764
rect 9276 64762 9332 64764
rect 9356 64762 9412 64764
rect 9116 64710 9162 64762
rect 9162 64710 9172 64762
rect 9196 64710 9226 64762
rect 9226 64710 9238 64762
rect 9238 64710 9252 64762
rect 9276 64710 9290 64762
rect 9290 64710 9302 64762
rect 9302 64710 9332 64762
rect 9356 64710 9366 64762
rect 9366 64710 9412 64762
rect 9116 64708 9172 64710
rect 9196 64708 9252 64710
rect 9276 64708 9332 64710
rect 9356 64708 9412 64710
rect 9116 63674 9172 63676
rect 9196 63674 9252 63676
rect 9276 63674 9332 63676
rect 9356 63674 9412 63676
rect 9116 63622 9162 63674
rect 9162 63622 9172 63674
rect 9196 63622 9226 63674
rect 9226 63622 9238 63674
rect 9238 63622 9252 63674
rect 9276 63622 9290 63674
rect 9290 63622 9302 63674
rect 9302 63622 9332 63674
rect 9356 63622 9366 63674
rect 9366 63622 9412 63674
rect 9116 63620 9172 63622
rect 9196 63620 9252 63622
rect 9276 63620 9332 63622
rect 9356 63620 9412 63622
rect 9310 63316 9312 63336
rect 9312 63316 9364 63336
rect 9364 63316 9366 63336
rect 9310 63280 9366 63316
rect 9116 62586 9172 62588
rect 9196 62586 9252 62588
rect 9276 62586 9332 62588
rect 9356 62586 9412 62588
rect 9116 62534 9162 62586
rect 9162 62534 9172 62586
rect 9196 62534 9226 62586
rect 9226 62534 9238 62586
rect 9238 62534 9252 62586
rect 9276 62534 9290 62586
rect 9290 62534 9302 62586
rect 9302 62534 9332 62586
rect 9356 62534 9366 62586
rect 9366 62534 9412 62586
rect 9116 62532 9172 62534
rect 9196 62532 9252 62534
rect 9276 62532 9332 62534
rect 9356 62532 9412 62534
rect 9116 61498 9172 61500
rect 9196 61498 9252 61500
rect 9276 61498 9332 61500
rect 9356 61498 9412 61500
rect 9116 61446 9162 61498
rect 9162 61446 9172 61498
rect 9196 61446 9226 61498
rect 9226 61446 9238 61498
rect 9238 61446 9252 61498
rect 9276 61446 9290 61498
rect 9290 61446 9302 61498
rect 9302 61446 9332 61498
rect 9356 61446 9366 61498
rect 9366 61446 9412 61498
rect 9116 61444 9172 61446
rect 9196 61444 9252 61446
rect 9276 61444 9332 61446
rect 9356 61444 9412 61446
rect 9116 60410 9172 60412
rect 9196 60410 9252 60412
rect 9276 60410 9332 60412
rect 9356 60410 9412 60412
rect 9116 60358 9162 60410
rect 9162 60358 9172 60410
rect 9196 60358 9226 60410
rect 9226 60358 9238 60410
rect 9238 60358 9252 60410
rect 9276 60358 9290 60410
rect 9290 60358 9302 60410
rect 9302 60358 9332 60410
rect 9356 60358 9366 60410
rect 9366 60358 9412 60410
rect 9116 60356 9172 60358
rect 9196 60356 9252 60358
rect 9276 60356 9332 60358
rect 9356 60356 9412 60358
rect 9310 59508 9312 59528
rect 9312 59508 9364 59528
rect 9364 59508 9366 59528
rect 9310 59472 9366 59508
rect 9116 59322 9172 59324
rect 9196 59322 9252 59324
rect 9276 59322 9332 59324
rect 9356 59322 9412 59324
rect 9116 59270 9162 59322
rect 9162 59270 9172 59322
rect 9196 59270 9226 59322
rect 9226 59270 9238 59322
rect 9238 59270 9252 59322
rect 9276 59270 9290 59322
rect 9290 59270 9302 59322
rect 9302 59270 9332 59322
rect 9356 59270 9366 59322
rect 9366 59270 9412 59322
rect 9116 59268 9172 59270
rect 9196 59268 9252 59270
rect 9276 59268 9332 59270
rect 9356 59268 9412 59270
rect 9116 58234 9172 58236
rect 9196 58234 9252 58236
rect 9276 58234 9332 58236
rect 9356 58234 9412 58236
rect 9116 58182 9162 58234
rect 9162 58182 9172 58234
rect 9196 58182 9226 58234
rect 9226 58182 9238 58234
rect 9238 58182 9252 58234
rect 9276 58182 9290 58234
rect 9290 58182 9302 58234
rect 9302 58182 9332 58234
rect 9356 58182 9366 58234
rect 9366 58182 9412 58234
rect 9116 58180 9172 58182
rect 9196 58180 9252 58182
rect 9276 58180 9332 58182
rect 9356 58180 9412 58182
rect 9494 57160 9550 57216
rect 9116 57146 9172 57148
rect 9196 57146 9252 57148
rect 9276 57146 9332 57148
rect 9356 57146 9412 57148
rect 9116 57094 9162 57146
rect 9162 57094 9172 57146
rect 9196 57094 9226 57146
rect 9226 57094 9238 57146
rect 9238 57094 9252 57146
rect 9276 57094 9290 57146
rect 9290 57094 9302 57146
rect 9302 57094 9332 57146
rect 9356 57094 9366 57146
rect 9366 57094 9412 57146
rect 9116 57092 9172 57094
rect 9196 57092 9252 57094
rect 9276 57092 9332 57094
rect 9356 57092 9412 57094
rect 9310 56344 9366 56400
rect 7484 54426 7540 54428
rect 7564 54426 7620 54428
rect 7644 54426 7700 54428
rect 7724 54426 7780 54428
rect 7484 54374 7530 54426
rect 7530 54374 7540 54426
rect 7564 54374 7594 54426
rect 7594 54374 7606 54426
rect 7606 54374 7620 54426
rect 7644 54374 7658 54426
rect 7658 54374 7670 54426
rect 7670 54374 7700 54426
rect 7724 54374 7734 54426
rect 7734 54374 7780 54426
rect 7484 54372 7540 54374
rect 7564 54372 7620 54374
rect 7644 54372 7700 54374
rect 7724 54372 7780 54374
rect 7484 53338 7540 53340
rect 7564 53338 7620 53340
rect 7644 53338 7700 53340
rect 7724 53338 7780 53340
rect 7484 53286 7530 53338
rect 7530 53286 7540 53338
rect 7564 53286 7594 53338
rect 7594 53286 7606 53338
rect 7606 53286 7620 53338
rect 7644 53286 7658 53338
rect 7658 53286 7670 53338
rect 7670 53286 7700 53338
rect 7724 53286 7734 53338
rect 7734 53286 7780 53338
rect 7484 53284 7540 53286
rect 7564 53284 7620 53286
rect 7644 53284 7700 53286
rect 7724 53284 7780 53286
rect 7484 52250 7540 52252
rect 7564 52250 7620 52252
rect 7644 52250 7700 52252
rect 7724 52250 7780 52252
rect 7484 52198 7530 52250
rect 7530 52198 7540 52250
rect 7564 52198 7594 52250
rect 7594 52198 7606 52250
rect 7606 52198 7620 52250
rect 7644 52198 7658 52250
rect 7658 52198 7670 52250
rect 7670 52198 7700 52250
rect 7724 52198 7734 52250
rect 7734 52198 7780 52250
rect 7484 52196 7540 52198
rect 7564 52196 7620 52198
rect 7644 52196 7700 52198
rect 7724 52196 7780 52198
rect 7484 51162 7540 51164
rect 7564 51162 7620 51164
rect 7644 51162 7700 51164
rect 7724 51162 7780 51164
rect 7484 51110 7530 51162
rect 7530 51110 7540 51162
rect 7564 51110 7594 51162
rect 7594 51110 7606 51162
rect 7606 51110 7620 51162
rect 7644 51110 7658 51162
rect 7658 51110 7670 51162
rect 7670 51110 7700 51162
rect 7724 51110 7734 51162
rect 7734 51110 7780 51162
rect 7484 51108 7540 51110
rect 7564 51108 7620 51110
rect 7644 51108 7700 51110
rect 7724 51108 7780 51110
rect 6550 41384 6606 41440
rect 5852 31034 5908 31036
rect 5932 31034 5988 31036
rect 6012 31034 6068 31036
rect 6092 31034 6148 31036
rect 5852 30982 5898 31034
rect 5898 30982 5908 31034
rect 5932 30982 5962 31034
rect 5962 30982 5974 31034
rect 5974 30982 5988 31034
rect 6012 30982 6026 31034
rect 6026 30982 6038 31034
rect 6038 30982 6068 31034
rect 6092 30982 6102 31034
rect 6102 30982 6148 31034
rect 5852 30980 5908 30982
rect 5932 30980 5988 30982
rect 6012 30980 6068 30982
rect 6092 30980 6148 30982
rect 7484 50074 7540 50076
rect 7564 50074 7620 50076
rect 7644 50074 7700 50076
rect 7724 50074 7780 50076
rect 7484 50022 7530 50074
rect 7530 50022 7540 50074
rect 7564 50022 7594 50074
rect 7594 50022 7606 50074
rect 7606 50022 7620 50074
rect 7644 50022 7658 50074
rect 7658 50022 7670 50074
rect 7670 50022 7700 50074
rect 7724 50022 7734 50074
rect 7734 50022 7780 50074
rect 7484 50020 7540 50022
rect 7564 50020 7620 50022
rect 7644 50020 7700 50022
rect 7724 50020 7780 50022
rect 7484 48986 7540 48988
rect 7564 48986 7620 48988
rect 7644 48986 7700 48988
rect 7724 48986 7780 48988
rect 7484 48934 7530 48986
rect 7530 48934 7540 48986
rect 7564 48934 7594 48986
rect 7594 48934 7606 48986
rect 7606 48934 7620 48986
rect 7644 48934 7658 48986
rect 7658 48934 7670 48986
rect 7670 48934 7700 48986
rect 7724 48934 7734 48986
rect 7734 48934 7780 48986
rect 7484 48932 7540 48934
rect 7564 48932 7620 48934
rect 7644 48932 7700 48934
rect 7724 48932 7780 48934
rect 7484 47898 7540 47900
rect 7564 47898 7620 47900
rect 7644 47898 7700 47900
rect 7724 47898 7780 47900
rect 7484 47846 7530 47898
rect 7530 47846 7540 47898
rect 7564 47846 7594 47898
rect 7594 47846 7606 47898
rect 7606 47846 7620 47898
rect 7644 47846 7658 47898
rect 7658 47846 7670 47898
rect 7670 47846 7700 47898
rect 7724 47846 7734 47898
rect 7734 47846 7780 47898
rect 7484 47844 7540 47846
rect 7564 47844 7620 47846
rect 7644 47844 7700 47846
rect 7724 47844 7780 47846
rect 7484 46810 7540 46812
rect 7564 46810 7620 46812
rect 7644 46810 7700 46812
rect 7724 46810 7780 46812
rect 7484 46758 7530 46810
rect 7530 46758 7540 46810
rect 7564 46758 7594 46810
rect 7594 46758 7606 46810
rect 7606 46758 7620 46810
rect 7644 46758 7658 46810
rect 7658 46758 7670 46810
rect 7670 46758 7700 46810
rect 7724 46758 7734 46810
rect 7734 46758 7780 46810
rect 7484 46756 7540 46758
rect 7564 46756 7620 46758
rect 7644 46756 7700 46758
rect 7724 46756 7780 46758
rect 7484 45722 7540 45724
rect 7564 45722 7620 45724
rect 7644 45722 7700 45724
rect 7724 45722 7780 45724
rect 7484 45670 7530 45722
rect 7530 45670 7540 45722
rect 7564 45670 7594 45722
rect 7594 45670 7606 45722
rect 7606 45670 7620 45722
rect 7644 45670 7658 45722
rect 7658 45670 7670 45722
rect 7670 45670 7700 45722
rect 7724 45670 7734 45722
rect 7734 45670 7780 45722
rect 7484 45668 7540 45670
rect 7564 45668 7620 45670
rect 7644 45668 7700 45670
rect 7724 45668 7780 45670
rect 7484 44634 7540 44636
rect 7564 44634 7620 44636
rect 7644 44634 7700 44636
rect 7724 44634 7780 44636
rect 7484 44582 7530 44634
rect 7530 44582 7540 44634
rect 7564 44582 7594 44634
rect 7594 44582 7606 44634
rect 7606 44582 7620 44634
rect 7644 44582 7658 44634
rect 7658 44582 7670 44634
rect 7670 44582 7700 44634
rect 7724 44582 7734 44634
rect 7734 44582 7780 44634
rect 7484 44580 7540 44582
rect 7564 44580 7620 44582
rect 7644 44580 7700 44582
rect 7724 44580 7780 44582
rect 7484 43546 7540 43548
rect 7564 43546 7620 43548
rect 7644 43546 7700 43548
rect 7724 43546 7780 43548
rect 7484 43494 7530 43546
rect 7530 43494 7540 43546
rect 7564 43494 7594 43546
rect 7594 43494 7606 43546
rect 7606 43494 7620 43546
rect 7644 43494 7658 43546
rect 7658 43494 7670 43546
rect 7670 43494 7700 43546
rect 7724 43494 7734 43546
rect 7734 43494 7780 43546
rect 7484 43492 7540 43494
rect 7564 43492 7620 43494
rect 7644 43492 7700 43494
rect 7724 43492 7780 43494
rect 9116 56058 9172 56060
rect 9196 56058 9252 56060
rect 9276 56058 9332 56060
rect 9356 56058 9412 56060
rect 9116 56006 9162 56058
rect 9162 56006 9172 56058
rect 9196 56006 9226 56058
rect 9226 56006 9238 56058
rect 9238 56006 9252 56058
rect 9276 56006 9290 56058
rect 9290 56006 9302 56058
rect 9302 56006 9332 56058
rect 9356 56006 9366 56058
rect 9366 56006 9412 56058
rect 9116 56004 9172 56006
rect 9196 56004 9252 56006
rect 9276 56004 9332 56006
rect 9356 56004 9412 56006
rect 9310 55700 9312 55720
rect 9312 55700 9364 55720
rect 9364 55700 9366 55720
rect 9310 55664 9366 55700
rect 9116 54970 9172 54972
rect 9196 54970 9252 54972
rect 9276 54970 9332 54972
rect 9356 54970 9412 54972
rect 9116 54918 9162 54970
rect 9162 54918 9172 54970
rect 9196 54918 9226 54970
rect 9226 54918 9238 54970
rect 9238 54918 9252 54970
rect 9276 54918 9290 54970
rect 9290 54918 9302 54970
rect 9302 54918 9332 54970
rect 9356 54918 9366 54970
rect 9366 54918 9412 54970
rect 9116 54916 9172 54918
rect 9196 54916 9252 54918
rect 9276 54916 9332 54918
rect 9356 54916 9412 54918
rect 9494 54848 9550 54904
rect 9116 53882 9172 53884
rect 9196 53882 9252 53884
rect 9276 53882 9332 53884
rect 9356 53882 9412 53884
rect 9116 53830 9162 53882
rect 9162 53830 9172 53882
rect 9196 53830 9226 53882
rect 9226 53830 9238 53882
rect 9238 53830 9252 53882
rect 9276 53830 9290 53882
rect 9290 53830 9302 53882
rect 9302 53830 9332 53882
rect 9356 53830 9366 53882
rect 9366 53830 9412 53882
rect 9116 53828 9172 53830
rect 9196 53828 9252 53830
rect 9276 53828 9332 53830
rect 9356 53828 9412 53830
rect 9116 52794 9172 52796
rect 9196 52794 9252 52796
rect 9276 52794 9332 52796
rect 9356 52794 9412 52796
rect 9116 52742 9162 52794
rect 9162 52742 9172 52794
rect 9196 52742 9226 52794
rect 9226 52742 9238 52794
rect 9238 52742 9252 52794
rect 9276 52742 9290 52794
rect 9290 52742 9302 52794
rect 9302 52742 9332 52794
rect 9356 52742 9366 52794
rect 9366 52742 9412 52794
rect 9116 52740 9172 52742
rect 9196 52740 9252 52742
rect 9276 52740 9332 52742
rect 9356 52740 9412 52742
rect 9116 51706 9172 51708
rect 9196 51706 9252 51708
rect 9276 51706 9332 51708
rect 9356 51706 9412 51708
rect 9116 51654 9162 51706
rect 9162 51654 9172 51706
rect 9196 51654 9226 51706
rect 9226 51654 9238 51706
rect 9238 51654 9252 51706
rect 9276 51654 9290 51706
rect 9290 51654 9302 51706
rect 9302 51654 9332 51706
rect 9356 51654 9366 51706
rect 9366 51654 9412 51706
rect 9116 51652 9172 51654
rect 9196 51652 9252 51654
rect 9276 51652 9332 51654
rect 9356 51652 9412 51654
rect 7484 42458 7540 42460
rect 7564 42458 7620 42460
rect 7644 42458 7700 42460
rect 7724 42458 7780 42460
rect 7484 42406 7530 42458
rect 7530 42406 7540 42458
rect 7564 42406 7594 42458
rect 7594 42406 7606 42458
rect 7606 42406 7620 42458
rect 7644 42406 7658 42458
rect 7658 42406 7670 42458
rect 7670 42406 7700 42458
rect 7724 42406 7734 42458
rect 7734 42406 7780 42458
rect 7484 42404 7540 42406
rect 7564 42404 7620 42406
rect 7644 42404 7700 42406
rect 7724 42404 7780 42406
rect 7484 41370 7540 41372
rect 7564 41370 7620 41372
rect 7644 41370 7700 41372
rect 7724 41370 7780 41372
rect 7484 41318 7530 41370
rect 7530 41318 7540 41370
rect 7564 41318 7594 41370
rect 7594 41318 7606 41370
rect 7606 41318 7620 41370
rect 7644 41318 7658 41370
rect 7658 41318 7670 41370
rect 7670 41318 7700 41370
rect 7724 41318 7734 41370
rect 7734 41318 7780 41370
rect 7484 41316 7540 41318
rect 7564 41316 7620 41318
rect 7644 41316 7700 41318
rect 7724 41316 7780 41318
rect 7484 40282 7540 40284
rect 7564 40282 7620 40284
rect 7644 40282 7700 40284
rect 7724 40282 7780 40284
rect 7484 40230 7530 40282
rect 7530 40230 7540 40282
rect 7564 40230 7594 40282
rect 7594 40230 7606 40282
rect 7606 40230 7620 40282
rect 7644 40230 7658 40282
rect 7658 40230 7670 40282
rect 7670 40230 7700 40282
rect 7724 40230 7734 40282
rect 7734 40230 7780 40282
rect 7484 40228 7540 40230
rect 7564 40228 7620 40230
rect 7644 40228 7700 40230
rect 7724 40228 7780 40230
rect 7484 39194 7540 39196
rect 7564 39194 7620 39196
rect 7644 39194 7700 39196
rect 7724 39194 7780 39196
rect 7484 39142 7530 39194
rect 7530 39142 7540 39194
rect 7564 39142 7594 39194
rect 7594 39142 7606 39194
rect 7606 39142 7620 39194
rect 7644 39142 7658 39194
rect 7658 39142 7670 39194
rect 7670 39142 7700 39194
rect 7724 39142 7734 39194
rect 7734 39142 7780 39194
rect 7484 39140 7540 39142
rect 7564 39140 7620 39142
rect 7644 39140 7700 39142
rect 7724 39140 7780 39142
rect 7484 38106 7540 38108
rect 7564 38106 7620 38108
rect 7644 38106 7700 38108
rect 7724 38106 7780 38108
rect 7484 38054 7530 38106
rect 7530 38054 7540 38106
rect 7564 38054 7594 38106
rect 7594 38054 7606 38106
rect 7606 38054 7620 38106
rect 7644 38054 7658 38106
rect 7658 38054 7670 38106
rect 7670 38054 7700 38106
rect 7724 38054 7734 38106
rect 7734 38054 7780 38106
rect 7484 38052 7540 38054
rect 7564 38052 7620 38054
rect 7644 38052 7700 38054
rect 7724 38052 7780 38054
rect 7484 37018 7540 37020
rect 7564 37018 7620 37020
rect 7644 37018 7700 37020
rect 7724 37018 7780 37020
rect 7484 36966 7530 37018
rect 7530 36966 7540 37018
rect 7564 36966 7594 37018
rect 7594 36966 7606 37018
rect 7606 36966 7620 37018
rect 7644 36966 7658 37018
rect 7658 36966 7670 37018
rect 7670 36966 7700 37018
rect 7724 36966 7734 37018
rect 7734 36966 7780 37018
rect 7484 36964 7540 36966
rect 7564 36964 7620 36966
rect 7644 36964 7700 36966
rect 7724 36964 7780 36966
rect 7484 35930 7540 35932
rect 7564 35930 7620 35932
rect 7644 35930 7700 35932
rect 7724 35930 7780 35932
rect 7484 35878 7530 35930
rect 7530 35878 7540 35930
rect 7564 35878 7594 35930
rect 7594 35878 7606 35930
rect 7606 35878 7620 35930
rect 7644 35878 7658 35930
rect 7658 35878 7670 35930
rect 7670 35878 7700 35930
rect 7724 35878 7734 35930
rect 7734 35878 7780 35930
rect 7484 35876 7540 35878
rect 7564 35876 7620 35878
rect 7644 35876 7700 35878
rect 7724 35876 7780 35878
rect 7484 34842 7540 34844
rect 7564 34842 7620 34844
rect 7644 34842 7700 34844
rect 7724 34842 7780 34844
rect 7484 34790 7530 34842
rect 7530 34790 7540 34842
rect 7564 34790 7594 34842
rect 7594 34790 7606 34842
rect 7606 34790 7620 34842
rect 7644 34790 7658 34842
rect 7658 34790 7670 34842
rect 7670 34790 7700 34842
rect 7724 34790 7734 34842
rect 7734 34790 7780 34842
rect 7484 34788 7540 34790
rect 7564 34788 7620 34790
rect 7644 34788 7700 34790
rect 7724 34788 7780 34790
rect 7484 33754 7540 33756
rect 7564 33754 7620 33756
rect 7644 33754 7700 33756
rect 7724 33754 7780 33756
rect 7484 33702 7530 33754
rect 7530 33702 7540 33754
rect 7564 33702 7594 33754
rect 7594 33702 7606 33754
rect 7606 33702 7620 33754
rect 7644 33702 7658 33754
rect 7658 33702 7670 33754
rect 7670 33702 7700 33754
rect 7724 33702 7734 33754
rect 7734 33702 7780 33754
rect 7484 33700 7540 33702
rect 7564 33700 7620 33702
rect 7644 33700 7700 33702
rect 7724 33700 7780 33702
rect 7484 32666 7540 32668
rect 7564 32666 7620 32668
rect 7644 32666 7700 32668
rect 7724 32666 7780 32668
rect 7484 32614 7530 32666
rect 7530 32614 7540 32666
rect 7564 32614 7594 32666
rect 7594 32614 7606 32666
rect 7606 32614 7620 32666
rect 7644 32614 7658 32666
rect 7658 32614 7670 32666
rect 7670 32614 7700 32666
rect 7724 32614 7734 32666
rect 7734 32614 7780 32666
rect 7484 32612 7540 32614
rect 7564 32612 7620 32614
rect 7644 32612 7700 32614
rect 7724 32612 7780 32614
rect 7484 31578 7540 31580
rect 7564 31578 7620 31580
rect 7644 31578 7700 31580
rect 7724 31578 7780 31580
rect 7484 31526 7530 31578
rect 7530 31526 7540 31578
rect 7564 31526 7594 31578
rect 7594 31526 7606 31578
rect 7606 31526 7620 31578
rect 7644 31526 7658 31578
rect 7658 31526 7670 31578
rect 7670 31526 7700 31578
rect 7724 31526 7734 31578
rect 7734 31526 7780 31578
rect 7484 31524 7540 31526
rect 7564 31524 7620 31526
rect 7644 31524 7700 31526
rect 7724 31524 7780 31526
rect 7484 30490 7540 30492
rect 7564 30490 7620 30492
rect 7644 30490 7700 30492
rect 7724 30490 7780 30492
rect 7484 30438 7530 30490
rect 7530 30438 7540 30490
rect 7564 30438 7594 30490
rect 7594 30438 7606 30490
rect 7606 30438 7620 30490
rect 7644 30438 7658 30490
rect 7658 30438 7670 30490
rect 7670 30438 7700 30490
rect 7724 30438 7734 30490
rect 7734 30438 7780 30490
rect 7484 30436 7540 30438
rect 7564 30436 7620 30438
rect 7644 30436 7700 30438
rect 7724 30436 7780 30438
rect 5852 29946 5908 29948
rect 5932 29946 5988 29948
rect 6012 29946 6068 29948
rect 6092 29946 6148 29948
rect 5852 29894 5898 29946
rect 5898 29894 5908 29946
rect 5932 29894 5962 29946
rect 5962 29894 5974 29946
rect 5974 29894 5988 29946
rect 6012 29894 6026 29946
rect 6026 29894 6038 29946
rect 6038 29894 6068 29946
rect 6092 29894 6102 29946
rect 6102 29894 6148 29946
rect 5852 29892 5908 29894
rect 5932 29892 5988 29894
rect 6012 29892 6068 29894
rect 6092 29892 6148 29894
rect 7484 29402 7540 29404
rect 7564 29402 7620 29404
rect 7644 29402 7700 29404
rect 7724 29402 7780 29404
rect 7484 29350 7530 29402
rect 7530 29350 7540 29402
rect 7564 29350 7594 29402
rect 7594 29350 7606 29402
rect 7606 29350 7620 29402
rect 7644 29350 7658 29402
rect 7658 29350 7670 29402
rect 7670 29350 7700 29402
rect 7724 29350 7734 29402
rect 7734 29350 7780 29402
rect 7484 29348 7540 29350
rect 7564 29348 7620 29350
rect 7644 29348 7700 29350
rect 7724 29348 7780 29350
rect 5852 28858 5908 28860
rect 5932 28858 5988 28860
rect 6012 28858 6068 28860
rect 6092 28858 6148 28860
rect 5852 28806 5898 28858
rect 5898 28806 5908 28858
rect 5932 28806 5962 28858
rect 5962 28806 5974 28858
rect 5974 28806 5988 28858
rect 6012 28806 6026 28858
rect 6026 28806 6038 28858
rect 6038 28806 6068 28858
rect 6092 28806 6102 28858
rect 6102 28806 6148 28858
rect 5852 28804 5908 28806
rect 5932 28804 5988 28806
rect 6012 28804 6068 28806
rect 6092 28804 6148 28806
rect 7484 28314 7540 28316
rect 7564 28314 7620 28316
rect 7644 28314 7700 28316
rect 7724 28314 7780 28316
rect 7484 28262 7530 28314
rect 7530 28262 7540 28314
rect 7564 28262 7594 28314
rect 7594 28262 7606 28314
rect 7606 28262 7620 28314
rect 7644 28262 7658 28314
rect 7658 28262 7670 28314
rect 7670 28262 7700 28314
rect 7724 28262 7734 28314
rect 7734 28262 7780 28314
rect 7484 28260 7540 28262
rect 7564 28260 7620 28262
rect 7644 28260 7700 28262
rect 7724 28260 7780 28262
rect 5852 27770 5908 27772
rect 5932 27770 5988 27772
rect 6012 27770 6068 27772
rect 6092 27770 6148 27772
rect 5852 27718 5898 27770
rect 5898 27718 5908 27770
rect 5932 27718 5962 27770
rect 5962 27718 5974 27770
rect 5974 27718 5988 27770
rect 6012 27718 6026 27770
rect 6026 27718 6038 27770
rect 6038 27718 6068 27770
rect 6092 27718 6102 27770
rect 6102 27718 6148 27770
rect 5852 27716 5908 27718
rect 5932 27716 5988 27718
rect 6012 27716 6068 27718
rect 6092 27716 6148 27718
rect 7484 27226 7540 27228
rect 7564 27226 7620 27228
rect 7644 27226 7700 27228
rect 7724 27226 7780 27228
rect 7484 27174 7530 27226
rect 7530 27174 7540 27226
rect 7564 27174 7594 27226
rect 7594 27174 7606 27226
rect 7606 27174 7620 27226
rect 7644 27174 7658 27226
rect 7658 27174 7670 27226
rect 7670 27174 7700 27226
rect 7724 27174 7734 27226
rect 7734 27174 7780 27226
rect 7484 27172 7540 27174
rect 7564 27172 7620 27174
rect 7644 27172 7700 27174
rect 7724 27172 7780 27174
rect 5852 26682 5908 26684
rect 5932 26682 5988 26684
rect 6012 26682 6068 26684
rect 6092 26682 6148 26684
rect 5852 26630 5898 26682
rect 5898 26630 5908 26682
rect 5932 26630 5962 26682
rect 5962 26630 5974 26682
rect 5974 26630 5988 26682
rect 6012 26630 6026 26682
rect 6026 26630 6038 26682
rect 6038 26630 6068 26682
rect 6092 26630 6102 26682
rect 6102 26630 6148 26682
rect 5852 26628 5908 26630
rect 5932 26628 5988 26630
rect 6012 26628 6068 26630
rect 6092 26628 6148 26630
rect 7484 26138 7540 26140
rect 7564 26138 7620 26140
rect 7644 26138 7700 26140
rect 7724 26138 7780 26140
rect 7484 26086 7530 26138
rect 7530 26086 7540 26138
rect 7564 26086 7594 26138
rect 7594 26086 7606 26138
rect 7606 26086 7620 26138
rect 7644 26086 7658 26138
rect 7658 26086 7670 26138
rect 7670 26086 7700 26138
rect 7724 26086 7734 26138
rect 7734 26086 7780 26138
rect 7484 26084 7540 26086
rect 7564 26084 7620 26086
rect 7644 26084 7700 26086
rect 7724 26084 7780 26086
rect 5852 25594 5908 25596
rect 5932 25594 5988 25596
rect 6012 25594 6068 25596
rect 6092 25594 6148 25596
rect 5852 25542 5898 25594
rect 5898 25542 5908 25594
rect 5932 25542 5962 25594
rect 5962 25542 5974 25594
rect 5974 25542 5988 25594
rect 6012 25542 6026 25594
rect 6026 25542 6038 25594
rect 6038 25542 6068 25594
rect 6092 25542 6102 25594
rect 6102 25542 6148 25594
rect 5852 25540 5908 25542
rect 5932 25540 5988 25542
rect 6012 25540 6068 25542
rect 6092 25540 6148 25542
rect 7484 25050 7540 25052
rect 7564 25050 7620 25052
rect 7644 25050 7700 25052
rect 7724 25050 7780 25052
rect 7484 24998 7530 25050
rect 7530 24998 7540 25050
rect 7564 24998 7594 25050
rect 7594 24998 7606 25050
rect 7606 24998 7620 25050
rect 7644 24998 7658 25050
rect 7658 24998 7670 25050
rect 7670 24998 7700 25050
rect 7724 24998 7734 25050
rect 7734 24998 7780 25050
rect 7484 24996 7540 24998
rect 7564 24996 7620 24998
rect 7644 24996 7700 24998
rect 7724 24996 7780 24998
rect 5852 24506 5908 24508
rect 5932 24506 5988 24508
rect 6012 24506 6068 24508
rect 6092 24506 6148 24508
rect 5852 24454 5898 24506
rect 5898 24454 5908 24506
rect 5932 24454 5962 24506
rect 5962 24454 5974 24506
rect 5974 24454 5988 24506
rect 6012 24454 6026 24506
rect 6026 24454 6038 24506
rect 6038 24454 6068 24506
rect 6092 24454 6102 24506
rect 6102 24454 6148 24506
rect 5852 24452 5908 24454
rect 5932 24452 5988 24454
rect 6012 24452 6068 24454
rect 6092 24452 6148 24454
rect 7484 23962 7540 23964
rect 7564 23962 7620 23964
rect 7644 23962 7700 23964
rect 7724 23962 7780 23964
rect 7484 23910 7530 23962
rect 7530 23910 7540 23962
rect 7564 23910 7594 23962
rect 7594 23910 7606 23962
rect 7606 23910 7620 23962
rect 7644 23910 7658 23962
rect 7658 23910 7670 23962
rect 7670 23910 7700 23962
rect 7724 23910 7734 23962
rect 7734 23910 7780 23962
rect 7484 23908 7540 23910
rect 7564 23908 7620 23910
rect 7644 23908 7700 23910
rect 7724 23908 7780 23910
rect 5852 23418 5908 23420
rect 5932 23418 5988 23420
rect 6012 23418 6068 23420
rect 6092 23418 6148 23420
rect 5852 23366 5898 23418
rect 5898 23366 5908 23418
rect 5932 23366 5962 23418
rect 5962 23366 5974 23418
rect 5974 23366 5988 23418
rect 6012 23366 6026 23418
rect 6026 23366 6038 23418
rect 6038 23366 6068 23418
rect 6092 23366 6102 23418
rect 6102 23366 6148 23418
rect 5852 23364 5908 23366
rect 5932 23364 5988 23366
rect 6012 23364 6068 23366
rect 6092 23364 6148 23366
rect 7484 22874 7540 22876
rect 7564 22874 7620 22876
rect 7644 22874 7700 22876
rect 7724 22874 7780 22876
rect 7484 22822 7530 22874
rect 7530 22822 7540 22874
rect 7564 22822 7594 22874
rect 7594 22822 7606 22874
rect 7606 22822 7620 22874
rect 7644 22822 7658 22874
rect 7658 22822 7670 22874
rect 7670 22822 7700 22874
rect 7724 22822 7734 22874
rect 7734 22822 7780 22874
rect 7484 22820 7540 22822
rect 7564 22820 7620 22822
rect 7644 22820 7700 22822
rect 7724 22820 7780 22822
rect 5852 22330 5908 22332
rect 5932 22330 5988 22332
rect 6012 22330 6068 22332
rect 6092 22330 6148 22332
rect 5852 22278 5898 22330
rect 5898 22278 5908 22330
rect 5932 22278 5962 22330
rect 5962 22278 5974 22330
rect 5974 22278 5988 22330
rect 6012 22278 6026 22330
rect 6026 22278 6038 22330
rect 6038 22278 6068 22330
rect 6092 22278 6102 22330
rect 6102 22278 6148 22330
rect 5852 22276 5908 22278
rect 5932 22276 5988 22278
rect 6012 22276 6068 22278
rect 6092 22276 6148 22278
rect 7484 21786 7540 21788
rect 7564 21786 7620 21788
rect 7644 21786 7700 21788
rect 7724 21786 7780 21788
rect 7484 21734 7530 21786
rect 7530 21734 7540 21786
rect 7564 21734 7594 21786
rect 7594 21734 7606 21786
rect 7606 21734 7620 21786
rect 7644 21734 7658 21786
rect 7658 21734 7670 21786
rect 7670 21734 7700 21786
rect 7724 21734 7734 21786
rect 7734 21734 7780 21786
rect 7484 21732 7540 21734
rect 7564 21732 7620 21734
rect 7644 21732 7700 21734
rect 7724 21732 7780 21734
rect 5852 21242 5908 21244
rect 5932 21242 5988 21244
rect 6012 21242 6068 21244
rect 6092 21242 6148 21244
rect 5852 21190 5898 21242
rect 5898 21190 5908 21242
rect 5932 21190 5962 21242
rect 5962 21190 5974 21242
rect 5974 21190 5988 21242
rect 6012 21190 6026 21242
rect 6026 21190 6038 21242
rect 6038 21190 6068 21242
rect 6092 21190 6102 21242
rect 6102 21190 6148 21242
rect 5852 21188 5908 21190
rect 5932 21188 5988 21190
rect 6012 21188 6068 21190
rect 6092 21188 6148 21190
rect 7484 20698 7540 20700
rect 7564 20698 7620 20700
rect 7644 20698 7700 20700
rect 7724 20698 7780 20700
rect 7484 20646 7530 20698
rect 7530 20646 7540 20698
rect 7564 20646 7594 20698
rect 7594 20646 7606 20698
rect 7606 20646 7620 20698
rect 7644 20646 7658 20698
rect 7658 20646 7670 20698
rect 7670 20646 7700 20698
rect 7724 20646 7734 20698
rect 7734 20646 7780 20698
rect 7484 20644 7540 20646
rect 7564 20644 7620 20646
rect 7644 20644 7700 20646
rect 7724 20644 7780 20646
rect 5852 20154 5908 20156
rect 5932 20154 5988 20156
rect 6012 20154 6068 20156
rect 6092 20154 6148 20156
rect 5852 20102 5898 20154
rect 5898 20102 5908 20154
rect 5932 20102 5962 20154
rect 5962 20102 5974 20154
rect 5974 20102 5988 20154
rect 6012 20102 6026 20154
rect 6026 20102 6038 20154
rect 6038 20102 6068 20154
rect 6092 20102 6102 20154
rect 6102 20102 6148 20154
rect 5852 20100 5908 20102
rect 5932 20100 5988 20102
rect 6012 20100 6068 20102
rect 6092 20100 6148 20102
rect 7484 19610 7540 19612
rect 7564 19610 7620 19612
rect 7644 19610 7700 19612
rect 7724 19610 7780 19612
rect 7484 19558 7530 19610
rect 7530 19558 7540 19610
rect 7564 19558 7594 19610
rect 7594 19558 7606 19610
rect 7606 19558 7620 19610
rect 7644 19558 7658 19610
rect 7658 19558 7670 19610
rect 7670 19558 7700 19610
rect 7724 19558 7734 19610
rect 7734 19558 7780 19610
rect 7484 19556 7540 19558
rect 7564 19556 7620 19558
rect 7644 19556 7700 19558
rect 7724 19556 7780 19558
rect 5852 19066 5908 19068
rect 5932 19066 5988 19068
rect 6012 19066 6068 19068
rect 6092 19066 6148 19068
rect 5852 19014 5898 19066
rect 5898 19014 5908 19066
rect 5932 19014 5962 19066
rect 5962 19014 5974 19066
rect 5974 19014 5988 19066
rect 6012 19014 6026 19066
rect 6026 19014 6038 19066
rect 6038 19014 6068 19066
rect 6092 19014 6102 19066
rect 6102 19014 6148 19066
rect 5852 19012 5908 19014
rect 5932 19012 5988 19014
rect 6012 19012 6068 19014
rect 6092 19012 6148 19014
rect 7484 18522 7540 18524
rect 7564 18522 7620 18524
rect 7644 18522 7700 18524
rect 7724 18522 7780 18524
rect 7484 18470 7530 18522
rect 7530 18470 7540 18522
rect 7564 18470 7594 18522
rect 7594 18470 7606 18522
rect 7606 18470 7620 18522
rect 7644 18470 7658 18522
rect 7658 18470 7670 18522
rect 7670 18470 7700 18522
rect 7724 18470 7734 18522
rect 7734 18470 7780 18522
rect 7484 18468 7540 18470
rect 7564 18468 7620 18470
rect 7644 18468 7700 18470
rect 7724 18468 7780 18470
rect 5852 17978 5908 17980
rect 5932 17978 5988 17980
rect 6012 17978 6068 17980
rect 6092 17978 6148 17980
rect 5852 17926 5898 17978
rect 5898 17926 5908 17978
rect 5932 17926 5962 17978
rect 5962 17926 5974 17978
rect 5974 17926 5988 17978
rect 6012 17926 6026 17978
rect 6026 17926 6038 17978
rect 6038 17926 6068 17978
rect 6092 17926 6102 17978
rect 6102 17926 6148 17978
rect 5852 17924 5908 17926
rect 5932 17924 5988 17926
rect 6012 17924 6068 17926
rect 6092 17924 6148 17926
rect 7484 17434 7540 17436
rect 7564 17434 7620 17436
rect 7644 17434 7700 17436
rect 7724 17434 7780 17436
rect 7484 17382 7530 17434
rect 7530 17382 7540 17434
rect 7564 17382 7594 17434
rect 7594 17382 7606 17434
rect 7606 17382 7620 17434
rect 7644 17382 7658 17434
rect 7658 17382 7670 17434
rect 7670 17382 7700 17434
rect 7724 17382 7734 17434
rect 7734 17382 7780 17434
rect 7484 17380 7540 17382
rect 7564 17380 7620 17382
rect 7644 17380 7700 17382
rect 7724 17380 7780 17382
rect 5852 16890 5908 16892
rect 5932 16890 5988 16892
rect 6012 16890 6068 16892
rect 6092 16890 6148 16892
rect 5852 16838 5898 16890
rect 5898 16838 5908 16890
rect 5932 16838 5962 16890
rect 5962 16838 5974 16890
rect 5974 16838 5988 16890
rect 6012 16838 6026 16890
rect 6026 16838 6038 16890
rect 6038 16838 6068 16890
rect 6092 16838 6102 16890
rect 6102 16838 6148 16890
rect 5852 16836 5908 16838
rect 5932 16836 5988 16838
rect 6012 16836 6068 16838
rect 6092 16836 6148 16838
rect 7484 16346 7540 16348
rect 7564 16346 7620 16348
rect 7644 16346 7700 16348
rect 7724 16346 7780 16348
rect 7484 16294 7530 16346
rect 7530 16294 7540 16346
rect 7564 16294 7594 16346
rect 7594 16294 7606 16346
rect 7606 16294 7620 16346
rect 7644 16294 7658 16346
rect 7658 16294 7670 16346
rect 7670 16294 7700 16346
rect 7724 16294 7734 16346
rect 7734 16294 7780 16346
rect 7484 16292 7540 16294
rect 7564 16292 7620 16294
rect 7644 16292 7700 16294
rect 7724 16292 7780 16294
rect 5852 15802 5908 15804
rect 5932 15802 5988 15804
rect 6012 15802 6068 15804
rect 6092 15802 6148 15804
rect 5852 15750 5898 15802
rect 5898 15750 5908 15802
rect 5932 15750 5962 15802
rect 5962 15750 5974 15802
rect 5974 15750 5988 15802
rect 6012 15750 6026 15802
rect 6026 15750 6038 15802
rect 6038 15750 6068 15802
rect 6092 15750 6102 15802
rect 6102 15750 6148 15802
rect 5852 15748 5908 15750
rect 5932 15748 5988 15750
rect 6012 15748 6068 15750
rect 6092 15748 6148 15750
rect 7484 15258 7540 15260
rect 7564 15258 7620 15260
rect 7644 15258 7700 15260
rect 7724 15258 7780 15260
rect 7484 15206 7530 15258
rect 7530 15206 7540 15258
rect 7564 15206 7594 15258
rect 7594 15206 7606 15258
rect 7606 15206 7620 15258
rect 7644 15206 7658 15258
rect 7658 15206 7670 15258
rect 7670 15206 7700 15258
rect 7724 15206 7734 15258
rect 7734 15206 7780 15258
rect 7484 15204 7540 15206
rect 7564 15204 7620 15206
rect 7644 15204 7700 15206
rect 7724 15204 7780 15206
rect 5852 14714 5908 14716
rect 5932 14714 5988 14716
rect 6012 14714 6068 14716
rect 6092 14714 6148 14716
rect 5852 14662 5898 14714
rect 5898 14662 5908 14714
rect 5932 14662 5962 14714
rect 5962 14662 5974 14714
rect 5974 14662 5988 14714
rect 6012 14662 6026 14714
rect 6026 14662 6038 14714
rect 6038 14662 6068 14714
rect 6092 14662 6102 14714
rect 6102 14662 6148 14714
rect 5852 14660 5908 14662
rect 5932 14660 5988 14662
rect 6012 14660 6068 14662
rect 6092 14660 6148 14662
rect 7484 14170 7540 14172
rect 7564 14170 7620 14172
rect 7644 14170 7700 14172
rect 7724 14170 7780 14172
rect 7484 14118 7530 14170
rect 7530 14118 7540 14170
rect 7564 14118 7594 14170
rect 7594 14118 7606 14170
rect 7606 14118 7620 14170
rect 7644 14118 7658 14170
rect 7658 14118 7670 14170
rect 7670 14118 7700 14170
rect 7724 14118 7734 14170
rect 7734 14118 7780 14170
rect 7484 14116 7540 14118
rect 7564 14116 7620 14118
rect 7644 14116 7700 14118
rect 7724 14116 7780 14118
rect 5852 13626 5908 13628
rect 5932 13626 5988 13628
rect 6012 13626 6068 13628
rect 6092 13626 6148 13628
rect 5852 13574 5898 13626
rect 5898 13574 5908 13626
rect 5932 13574 5962 13626
rect 5962 13574 5974 13626
rect 5974 13574 5988 13626
rect 6012 13574 6026 13626
rect 6026 13574 6038 13626
rect 6038 13574 6068 13626
rect 6092 13574 6102 13626
rect 6102 13574 6148 13626
rect 5852 13572 5908 13574
rect 5932 13572 5988 13574
rect 6012 13572 6068 13574
rect 6092 13572 6148 13574
rect 7484 13082 7540 13084
rect 7564 13082 7620 13084
rect 7644 13082 7700 13084
rect 7724 13082 7780 13084
rect 7484 13030 7530 13082
rect 7530 13030 7540 13082
rect 7564 13030 7594 13082
rect 7594 13030 7606 13082
rect 7606 13030 7620 13082
rect 7644 13030 7658 13082
rect 7658 13030 7670 13082
rect 7670 13030 7700 13082
rect 7724 13030 7734 13082
rect 7734 13030 7780 13082
rect 7484 13028 7540 13030
rect 7564 13028 7620 13030
rect 7644 13028 7700 13030
rect 7724 13028 7780 13030
rect 5852 12538 5908 12540
rect 5932 12538 5988 12540
rect 6012 12538 6068 12540
rect 6092 12538 6148 12540
rect 5852 12486 5898 12538
rect 5898 12486 5908 12538
rect 5932 12486 5962 12538
rect 5962 12486 5974 12538
rect 5974 12486 5988 12538
rect 6012 12486 6026 12538
rect 6026 12486 6038 12538
rect 6038 12486 6068 12538
rect 6092 12486 6102 12538
rect 6102 12486 6148 12538
rect 5852 12484 5908 12486
rect 5932 12484 5988 12486
rect 6012 12484 6068 12486
rect 6092 12484 6148 12486
rect 7484 11994 7540 11996
rect 7564 11994 7620 11996
rect 7644 11994 7700 11996
rect 7724 11994 7780 11996
rect 7484 11942 7530 11994
rect 7530 11942 7540 11994
rect 7564 11942 7594 11994
rect 7594 11942 7606 11994
rect 7606 11942 7620 11994
rect 7644 11942 7658 11994
rect 7658 11942 7670 11994
rect 7670 11942 7700 11994
rect 7724 11942 7734 11994
rect 7734 11942 7780 11994
rect 7484 11940 7540 11942
rect 7564 11940 7620 11942
rect 7644 11940 7700 11942
rect 7724 11940 7780 11942
rect 5852 11450 5908 11452
rect 5932 11450 5988 11452
rect 6012 11450 6068 11452
rect 6092 11450 6148 11452
rect 5852 11398 5898 11450
rect 5898 11398 5908 11450
rect 5932 11398 5962 11450
rect 5962 11398 5974 11450
rect 5974 11398 5988 11450
rect 6012 11398 6026 11450
rect 6026 11398 6038 11450
rect 6038 11398 6068 11450
rect 6092 11398 6102 11450
rect 6102 11398 6148 11450
rect 5852 11396 5908 11398
rect 5932 11396 5988 11398
rect 6012 11396 6068 11398
rect 6092 11396 6148 11398
rect 7484 10906 7540 10908
rect 7564 10906 7620 10908
rect 7644 10906 7700 10908
rect 7724 10906 7780 10908
rect 7484 10854 7530 10906
rect 7530 10854 7540 10906
rect 7564 10854 7594 10906
rect 7594 10854 7606 10906
rect 7606 10854 7620 10906
rect 7644 10854 7658 10906
rect 7658 10854 7670 10906
rect 7670 10854 7700 10906
rect 7724 10854 7734 10906
rect 7734 10854 7780 10906
rect 7484 10852 7540 10854
rect 7564 10852 7620 10854
rect 7644 10852 7700 10854
rect 7724 10852 7780 10854
rect 5852 10362 5908 10364
rect 5932 10362 5988 10364
rect 6012 10362 6068 10364
rect 6092 10362 6148 10364
rect 5852 10310 5898 10362
rect 5898 10310 5908 10362
rect 5932 10310 5962 10362
rect 5962 10310 5974 10362
rect 5974 10310 5988 10362
rect 6012 10310 6026 10362
rect 6026 10310 6038 10362
rect 6038 10310 6068 10362
rect 6092 10310 6102 10362
rect 6102 10310 6148 10362
rect 5852 10308 5908 10310
rect 5932 10308 5988 10310
rect 6012 10308 6068 10310
rect 6092 10308 6148 10310
rect 7484 9818 7540 9820
rect 7564 9818 7620 9820
rect 7644 9818 7700 9820
rect 7724 9818 7780 9820
rect 7484 9766 7530 9818
rect 7530 9766 7540 9818
rect 7564 9766 7594 9818
rect 7594 9766 7606 9818
rect 7606 9766 7620 9818
rect 7644 9766 7658 9818
rect 7658 9766 7670 9818
rect 7670 9766 7700 9818
rect 7724 9766 7734 9818
rect 7734 9766 7780 9818
rect 7484 9764 7540 9766
rect 7564 9764 7620 9766
rect 7644 9764 7700 9766
rect 7724 9764 7780 9766
rect 9116 50618 9172 50620
rect 9196 50618 9252 50620
rect 9276 50618 9332 50620
rect 9356 50618 9412 50620
rect 9116 50566 9162 50618
rect 9162 50566 9172 50618
rect 9196 50566 9226 50618
rect 9226 50566 9238 50618
rect 9238 50566 9252 50618
rect 9276 50566 9290 50618
rect 9290 50566 9302 50618
rect 9302 50566 9332 50618
rect 9356 50566 9366 50618
rect 9366 50566 9412 50618
rect 9116 50564 9172 50566
rect 9196 50564 9252 50566
rect 9276 50564 9332 50566
rect 9356 50564 9412 50566
rect 9116 49530 9172 49532
rect 9196 49530 9252 49532
rect 9276 49530 9332 49532
rect 9356 49530 9412 49532
rect 9116 49478 9162 49530
rect 9162 49478 9172 49530
rect 9196 49478 9226 49530
rect 9226 49478 9238 49530
rect 9238 49478 9252 49530
rect 9276 49478 9290 49530
rect 9290 49478 9302 49530
rect 9302 49478 9332 49530
rect 9356 49478 9366 49530
rect 9366 49478 9412 49530
rect 9116 49476 9172 49478
rect 9196 49476 9252 49478
rect 9276 49476 9332 49478
rect 9356 49476 9412 49478
rect 9586 49408 9642 49464
rect 9116 48442 9172 48444
rect 9196 48442 9252 48444
rect 9276 48442 9332 48444
rect 9356 48442 9412 48444
rect 9116 48390 9162 48442
rect 9162 48390 9172 48442
rect 9196 48390 9226 48442
rect 9226 48390 9238 48442
rect 9238 48390 9252 48442
rect 9276 48390 9290 48442
rect 9290 48390 9302 48442
rect 9302 48390 9332 48442
rect 9356 48390 9366 48442
rect 9366 48390 9412 48442
rect 9116 48388 9172 48390
rect 9196 48388 9252 48390
rect 9276 48388 9332 48390
rect 9356 48388 9412 48390
rect 9116 47354 9172 47356
rect 9196 47354 9252 47356
rect 9276 47354 9332 47356
rect 9356 47354 9412 47356
rect 9116 47302 9162 47354
rect 9162 47302 9172 47354
rect 9196 47302 9226 47354
rect 9226 47302 9238 47354
rect 9238 47302 9252 47354
rect 9276 47302 9290 47354
rect 9290 47302 9302 47354
rect 9302 47302 9332 47354
rect 9356 47302 9366 47354
rect 9366 47302 9412 47354
rect 9116 47300 9172 47302
rect 9196 47300 9252 47302
rect 9276 47300 9332 47302
rect 9356 47300 9412 47302
rect 9116 46266 9172 46268
rect 9196 46266 9252 46268
rect 9276 46266 9332 46268
rect 9356 46266 9412 46268
rect 9116 46214 9162 46266
rect 9162 46214 9172 46266
rect 9196 46214 9226 46266
rect 9226 46214 9238 46266
rect 9238 46214 9252 46266
rect 9276 46214 9290 46266
rect 9290 46214 9302 46266
rect 9302 46214 9332 46266
rect 9356 46214 9366 46266
rect 9366 46214 9412 46266
rect 9116 46212 9172 46214
rect 9196 46212 9252 46214
rect 9276 46212 9332 46214
rect 9356 46212 9412 46214
rect 9116 45178 9172 45180
rect 9196 45178 9252 45180
rect 9276 45178 9332 45180
rect 9356 45178 9412 45180
rect 9116 45126 9162 45178
rect 9162 45126 9172 45178
rect 9196 45126 9226 45178
rect 9226 45126 9238 45178
rect 9238 45126 9252 45178
rect 9276 45126 9290 45178
rect 9290 45126 9302 45178
rect 9302 45126 9332 45178
rect 9356 45126 9366 45178
rect 9366 45126 9412 45178
rect 9116 45124 9172 45126
rect 9196 45124 9252 45126
rect 9276 45124 9332 45126
rect 9356 45124 9412 45126
rect 9116 44090 9172 44092
rect 9196 44090 9252 44092
rect 9276 44090 9332 44092
rect 9356 44090 9412 44092
rect 9116 44038 9162 44090
rect 9162 44038 9172 44090
rect 9196 44038 9226 44090
rect 9226 44038 9238 44090
rect 9238 44038 9252 44090
rect 9276 44038 9290 44090
rect 9290 44038 9302 44090
rect 9302 44038 9332 44090
rect 9356 44038 9366 44090
rect 9366 44038 9412 44090
rect 9116 44036 9172 44038
rect 9196 44036 9252 44038
rect 9276 44036 9332 44038
rect 9356 44036 9412 44038
rect 9116 43002 9172 43004
rect 9196 43002 9252 43004
rect 9276 43002 9332 43004
rect 9356 43002 9412 43004
rect 9116 42950 9162 43002
rect 9162 42950 9172 43002
rect 9196 42950 9226 43002
rect 9226 42950 9238 43002
rect 9238 42950 9252 43002
rect 9276 42950 9290 43002
rect 9290 42950 9302 43002
rect 9302 42950 9332 43002
rect 9356 42950 9366 43002
rect 9366 42950 9412 43002
rect 9116 42948 9172 42950
rect 9196 42948 9252 42950
rect 9276 42948 9332 42950
rect 9356 42948 9412 42950
rect 9116 41914 9172 41916
rect 9196 41914 9252 41916
rect 9276 41914 9332 41916
rect 9356 41914 9412 41916
rect 9116 41862 9162 41914
rect 9162 41862 9172 41914
rect 9196 41862 9226 41914
rect 9226 41862 9238 41914
rect 9238 41862 9252 41914
rect 9276 41862 9290 41914
rect 9290 41862 9302 41914
rect 9302 41862 9332 41914
rect 9356 41862 9366 41914
rect 9366 41862 9412 41914
rect 9116 41860 9172 41862
rect 9196 41860 9252 41862
rect 9276 41860 9332 41862
rect 9356 41860 9412 41862
rect 9116 40826 9172 40828
rect 9196 40826 9252 40828
rect 9276 40826 9332 40828
rect 9356 40826 9412 40828
rect 9116 40774 9162 40826
rect 9162 40774 9172 40826
rect 9196 40774 9226 40826
rect 9226 40774 9238 40826
rect 9238 40774 9252 40826
rect 9276 40774 9290 40826
rect 9290 40774 9302 40826
rect 9302 40774 9332 40826
rect 9356 40774 9366 40826
rect 9366 40774 9412 40826
rect 9116 40772 9172 40774
rect 9196 40772 9252 40774
rect 9276 40772 9332 40774
rect 9356 40772 9412 40774
rect 10138 76372 10140 76392
rect 10140 76372 10192 76392
rect 10192 76372 10194 76392
rect 10138 76336 10194 76372
rect 10138 75656 10194 75712
rect 10138 74840 10194 74896
rect 10138 74024 10194 74080
rect 10138 73344 10194 73400
rect 10138 72528 10194 72584
rect 10138 71712 10194 71768
rect 10138 71032 10194 71088
rect 10138 70216 10194 70272
rect 10138 69400 10194 69456
rect 10138 68756 10140 68776
rect 10140 68756 10192 68776
rect 10192 68756 10194 68776
rect 10138 68720 10194 68756
rect 10138 67904 10194 67960
rect 10138 67088 10194 67144
rect 10138 66408 10194 66464
rect 10138 65592 10194 65648
rect 10138 64776 10194 64832
rect 10138 64096 10194 64152
rect 10138 62464 10194 62520
rect 10138 61784 10194 61840
rect 10138 60968 10194 61024
rect 10138 60288 10194 60344
rect 10138 58656 10194 58712
rect 10138 57976 10194 58032
rect 10046 54052 10102 54088
rect 10046 54032 10048 54052
rect 10048 54032 10100 54052
rect 10100 54032 10102 54052
rect 10046 53388 10048 53408
rect 10048 53388 10100 53408
rect 10100 53388 10102 53408
rect 10046 53352 10102 53388
rect 10046 52536 10102 52592
rect 10046 51756 10048 51776
rect 10048 51756 10100 51776
rect 10100 51756 10102 51776
rect 10046 51720 10102 51756
rect 10046 51040 10102 51096
rect 10046 50224 10102 50280
rect 10046 48728 10102 48784
rect 10046 47948 10048 47968
rect 10048 47948 10100 47968
rect 10100 47948 10102 47968
rect 10046 47912 10102 47948
rect 10046 47096 10102 47152
rect 10046 46436 10102 46472
rect 10046 46416 10048 46436
rect 10048 46416 10100 46436
rect 10100 46416 10102 46436
rect 10046 45600 10102 45656
rect 10046 44784 10102 44840
rect 10046 44140 10048 44160
rect 10048 44140 10100 44160
rect 10100 44140 10102 44160
rect 10046 44104 10102 44140
rect 10046 43288 10102 43344
rect 10046 42508 10048 42528
rect 10048 42508 10100 42528
rect 10100 42508 10102 42528
rect 10046 42472 10102 42508
rect 10046 41792 10102 41848
rect 9116 39738 9172 39740
rect 9196 39738 9252 39740
rect 9276 39738 9332 39740
rect 9356 39738 9412 39740
rect 9116 39686 9162 39738
rect 9162 39686 9172 39738
rect 9196 39686 9226 39738
rect 9226 39686 9238 39738
rect 9238 39686 9252 39738
rect 9276 39686 9290 39738
rect 9290 39686 9302 39738
rect 9302 39686 9332 39738
rect 9356 39686 9366 39738
rect 9366 39686 9412 39738
rect 9116 39684 9172 39686
rect 9196 39684 9252 39686
rect 9276 39684 9332 39686
rect 9356 39684 9412 39686
rect 9116 38650 9172 38652
rect 9196 38650 9252 38652
rect 9276 38650 9332 38652
rect 9356 38650 9412 38652
rect 9116 38598 9162 38650
rect 9162 38598 9172 38650
rect 9196 38598 9226 38650
rect 9226 38598 9238 38650
rect 9238 38598 9252 38650
rect 9276 38598 9290 38650
rect 9290 38598 9302 38650
rect 9302 38598 9332 38650
rect 9356 38598 9366 38650
rect 9366 38598 9412 38650
rect 9116 38596 9172 38598
rect 9196 38596 9252 38598
rect 9276 38596 9332 38598
rect 9356 38596 9412 38598
rect 9116 37562 9172 37564
rect 9196 37562 9252 37564
rect 9276 37562 9332 37564
rect 9356 37562 9412 37564
rect 9116 37510 9162 37562
rect 9162 37510 9172 37562
rect 9196 37510 9226 37562
rect 9226 37510 9238 37562
rect 9238 37510 9252 37562
rect 9276 37510 9290 37562
rect 9290 37510 9302 37562
rect 9302 37510 9332 37562
rect 9356 37510 9366 37562
rect 9366 37510 9412 37562
rect 9116 37508 9172 37510
rect 9196 37508 9252 37510
rect 9276 37508 9332 37510
rect 9356 37508 9412 37510
rect 9116 36474 9172 36476
rect 9196 36474 9252 36476
rect 9276 36474 9332 36476
rect 9356 36474 9412 36476
rect 9116 36422 9162 36474
rect 9162 36422 9172 36474
rect 9196 36422 9226 36474
rect 9226 36422 9238 36474
rect 9238 36422 9252 36474
rect 9276 36422 9290 36474
rect 9290 36422 9302 36474
rect 9302 36422 9332 36474
rect 9356 36422 9366 36474
rect 9366 36422 9412 36474
rect 9116 36420 9172 36422
rect 9196 36420 9252 36422
rect 9276 36420 9332 36422
rect 9356 36420 9412 36422
rect 9116 35386 9172 35388
rect 9196 35386 9252 35388
rect 9276 35386 9332 35388
rect 9356 35386 9412 35388
rect 9116 35334 9162 35386
rect 9162 35334 9172 35386
rect 9196 35334 9226 35386
rect 9226 35334 9238 35386
rect 9238 35334 9252 35386
rect 9276 35334 9290 35386
rect 9290 35334 9302 35386
rect 9302 35334 9332 35386
rect 9356 35334 9366 35386
rect 9366 35334 9412 35386
rect 9116 35332 9172 35334
rect 9196 35332 9252 35334
rect 9276 35332 9332 35334
rect 9356 35332 9412 35334
rect 9116 34298 9172 34300
rect 9196 34298 9252 34300
rect 9276 34298 9332 34300
rect 9356 34298 9412 34300
rect 9116 34246 9162 34298
rect 9162 34246 9172 34298
rect 9196 34246 9226 34298
rect 9226 34246 9238 34298
rect 9238 34246 9252 34298
rect 9276 34246 9290 34298
rect 9290 34246 9302 34298
rect 9302 34246 9332 34298
rect 9356 34246 9366 34298
rect 9366 34246 9412 34298
rect 9116 34244 9172 34246
rect 9196 34244 9252 34246
rect 9276 34244 9332 34246
rect 9356 34244 9412 34246
rect 9586 34040 9642 34096
rect 9116 33210 9172 33212
rect 9196 33210 9252 33212
rect 9276 33210 9332 33212
rect 9356 33210 9412 33212
rect 9116 33158 9162 33210
rect 9162 33158 9172 33210
rect 9196 33158 9226 33210
rect 9226 33158 9238 33210
rect 9238 33158 9252 33210
rect 9276 33158 9290 33210
rect 9290 33158 9302 33210
rect 9302 33158 9332 33210
rect 9356 33158 9366 33210
rect 9366 33158 9412 33210
rect 9116 33156 9172 33158
rect 9196 33156 9252 33158
rect 9276 33156 9332 33158
rect 9356 33156 9412 33158
rect 10046 40996 10102 41032
rect 10046 40976 10048 40996
rect 10048 40976 10100 40996
rect 10100 40976 10102 40996
rect 10046 40332 10048 40352
rect 10048 40332 10100 40352
rect 10100 40332 10102 40352
rect 10046 40296 10102 40332
rect 10046 39480 10102 39536
rect 10046 38700 10048 38720
rect 10048 38700 10100 38720
rect 10100 38700 10102 38720
rect 10046 38664 10102 38700
rect 10046 37984 10102 38040
rect 10046 37168 10102 37224
rect 10046 36352 10102 36408
rect 10046 35672 10102 35728
rect 10046 34892 10048 34912
rect 10048 34892 10100 34912
rect 10100 34892 10102 34912
rect 10046 34856 10102 34892
rect 9116 32122 9172 32124
rect 9196 32122 9252 32124
rect 9276 32122 9332 32124
rect 9356 32122 9412 32124
rect 9116 32070 9162 32122
rect 9162 32070 9172 32122
rect 9196 32070 9226 32122
rect 9226 32070 9238 32122
rect 9238 32070 9252 32122
rect 9276 32070 9290 32122
rect 9290 32070 9302 32122
rect 9302 32070 9332 32122
rect 9356 32070 9366 32122
rect 9366 32070 9412 32122
rect 9116 32068 9172 32070
rect 9196 32068 9252 32070
rect 9276 32068 9332 32070
rect 9356 32068 9412 32070
rect 9116 31034 9172 31036
rect 9196 31034 9252 31036
rect 9276 31034 9332 31036
rect 9356 31034 9412 31036
rect 9116 30982 9162 31034
rect 9162 30982 9172 31034
rect 9196 30982 9226 31034
rect 9226 30982 9238 31034
rect 9238 30982 9252 31034
rect 9276 30982 9290 31034
rect 9290 30982 9302 31034
rect 9302 30982 9332 31034
rect 9356 30982 9366 31034
rect 9366 30982 9412 31034
rect 9116 30980 9172 30982
rect 9196 30980 9252 30982
rect 9276 30980 9332 30982
rect 9356 30980 9412 30982
rect 9116 29946 9172 29948
rect 9196 29946 9252 29948
rect 9276 29946 9332 29948
rect 9356 29946 9412 29948
rect 9116 29894 9162 29946
rect 9162 29894 9172 29946
rect 9196 29894 9226 29946
rect 9226 29894 9238 29946
rect 9238 29894 9252 29946
rect 9276 29894 9290 29946
rect 9290 29894 9302 29946
rect 9302 29894 9332 29946
rect 9356 29894 9366 29946
rect 9366 29894 9412 29946
rect 9116 29892 9172 29894
rect 9196 29892 9252 29894
rect 9276 29892 9332 29894
rect 9356 29892 9412 29894
rect 9116 28858 9172 28860
rect 9196 28858 9252 28860
rect 9276 28858 9332 28860
rect 9356 28858 9412 28860
rect 9116 28806 9162 28858
rect 9162 28806 9172 28858
rect 9196 28806 9226 28858
rect 9226 28806 9238 28858
rect 9238 28806 9252 28858
rect 9276 28806 9290 28858
rect 9290 28806 9302 28858
rect 9302 28806 9332 28858
rect 9356 28806 9366 28858
rect 9366 28806 9412 28858
rect 9116 28804 9172 28806
rect 9196 28804 9252 28806
rect 9276 28804 9332 28806
rect 9356 28804 9412 28806
rect 10046 33380 10102 33416
rect 10046 33360 10048 33380
rect 10048 33360 10100 33380
rect 10100 33360 10102 33380
rect 10046 32544 10102 32600
rect 10046 31728 10102 31784
rect 10046 31084 10048 31104
rect 10048 31084 10100 31104
rect 10100 31084 10102 31104
rect 10046 31048 10102 31084
rect 10046 30232 10102 30288
rect 10138 29416 10194 29472
rect 10138 28736 10194 28792
rect 9954 27956 9956 27976
rect 9956 27956 10008 27976
rect 10008 27956 10010 27976
rect 9954 27920 10010 27956
rect 9116 27770 9172 27772
rect 9196 27770 9252 27772
rect 9276 27770 9332 27772
rect 9356 27770 9412 27772
rect 9116 27718 9162 27770
rect 9162 27718 9172 27770
rect 9196 27718 9226 27770
rect 9226 27718 9238 27770
rect 9238 27718 9252 27770
rect 9276 27718 9290 27770
rect 9290 27718 9302 27770
rect 9302 27718 9332 27770
rect 9356 27718 9366 27770
rect 9366 27718 9412 27770
rect 9116 27716 9172 27718
rect 9196 27716 9252 27718
rect 9276 27716 9332 27718
rect 9356 27716 9412 27718
rect 9954 27104 10010 27160
rect 9116 26682 9172 26684
rect 9196 26682 9252 26684
rect 9276 26682 9332 26684
rect 9356 26682 9412 26684
rect 9116 26630 9162 26682
rect 9162 26630 9172 26682
rect 9196 26630 9226 26682
rect 9226 26630 9238 26682
rect 9238 26630 9252 26682
rect 9276 26630 9290 26682
rect 9290 26630 9302 26682
rect 9302 26630 9332 26682
rect 9356 26630 9366 26682
rect 9366 26630 9412 26682
rect 9116 26628 9172 26630
rect 9196 26628 9252 26630
rect 9276 26628 9332 26630
rect 9356 26628 9412 26630
rect 10138 26424 10194 26480
rect 10138 25644 10140 25664
rect 10140 25644 10192 25664
rect 10192 25644 10194 25664
rect 10138 25608 10194 25644
rect 9116 25594 9172 25596
rect 9196 25594 9252 25596
rect 9276 25594 9332 25596
rect 9356 25594 9412 25596
rect 9116 25542 9162 25594
rect 9162 25542 9172 25594
rect 9196 25542 9226 25594
rect 9226 25542 9238 25594
rect 9238 25542 9252 25594
rect 9276 25542 9290 25594
rect 9290 25542 9302 25594
rect 9302 25542 9332 25594
rect 9356 25542 9366 25594
rect 9366 25542 9412 25594
rect 9116 25540 9172 25542
rect 9196 25540 9252 25542
rect 9276 25540 9332 25542
rect 9356 25540 9412 25542
rect 10138 24792 10194 24848
rect 9116 24506 9172 24508
rect 9196 24506 9252 24508
rect 9276 24506 9332 24508
rect 9356 24506 9412 24508
rect 9116 24454 9162 24506
rect 9162 24454 9172 24506
rect 9196 24454 9226 24506
rect 9226 24454 9238 24506
rect 9238 24454 9252 24506
rect 9276 24454 9290 24506
rect 9290 24454 9302 24506
rect 9302 24454 9332 24506
rect 9356 24454 9366 24506
rect 9366 24454 9412 24506
rect 9116 24452 9172 24454
rect 9196 24452 9252 24454
rect 9276 24452 9332 24454
rect 9356 24452 9412 24454
rect 10138 24148 10140 24168
rect 10140 24148 10192 24168
rect 10192 24148 10194 24168
rect 10138 24112 10194 24148
rect 9116 23418 9172 23420
rect 9196 23418 9252 23420
rect 9276 23418 9332 23420
rect 9356 23418 9412 23420
rect 9116 23366 9162 23418
rect 9162 23366 9172 23418
rect 9196 23366 9226 23418
rect 9226 23366 9238 23418
rect 9238 23366 9252 23418
rect 9276 23366 9290 23418
rect 9290 23366 9302 23418
rect 9302 23366 9332 23418
rect 9356 23366 9366 23418
rect 9366 23366 9412 23418
rect 9116 23364 9172 23366
rect 9196 23364 9252 23366
rect 9276 23364 9332 23366
rect 9356 23364 9412 23366
rect 10138 23296 10194 23352
rect 10138 22500 10194 22536
rect 10138 22480 10140 22500
rect 10140 22480 10192 22500
rect 10192 22480 10194 22500
rect 9116 22330 9172 22332
rect 9196 22330 9252 22332
rect 9276 22330 9332 22332
rect 9356 22330 9412 22332
rect 9116 22278 9162 22330
rect 9162 22278 9172 22330
rect 9196 22278 9226 22330
rect 9226 22278 9238 22330
rect 9238 22278 9252 22330
rect 9276 22278 9290 22330
rect 9290 22278 9302 22330
rect 9302 22278 9332 22330
rect 9356 22278 9366 22330
rect 9366 22278 9412 22330
rect 9116 22276 9172 22278
rect 9196 22276 9252 22278
rect 9276 22276 9332 22278
rect 9356 22276 9412 22278
rect 10138 21800 10194 21856
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 9276 21242 9332 21244
rect 9356 21242 9412 21244
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9238 21242
rect 9238 21190 9252 21242
rect 9276 21190 9290 21242
rect 9290 21190 9302 21242
rect 9302 21190 9332 21242
rect 9356 21190 9366 21242
rect 9366 21190 9412 21242
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 9276 21188 9332 21190
rect 9356 21188 9412 21190
rect 10138 20984 10194 21040
rect 10046 20324 10102 20360
rect 10046 20304 10048 20324
rect 10048 20304 10100 20324
rect 10100 20304 10102 20324
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 9276 20154 9332 20156
rect 9356 20154 9412 20156
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9238 20154
rect 9238 20102 9252 20154
rect 9276 20102 9290 20154
rect 9290 20102 9302 20154
rect 9302 20102 9332 20154
rect 9356 20102 9366 20154
rect 9366 20102 9412 20154
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 9276 20100 9332 20102
rect 9356 20100 9412 20102
rect 10046 19488 10102 19544
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 9276 19066 9332 19068
rect 9356 19066 9412 19068
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9238 19066
rect 9238 19014 9252 19066
rect 9276 19014 9290 19066
rect 9290 19014 9302 19066
rect 9302 19014 9332 19066
rect 9356 19014 9366 19066
rect 9366 19014 9412 19066
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 9276 19012 9332 19014
rect 9356 19012 9412 19014
rect 10046 18672 10102 18728
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 9276 17978 9332 17980
rect 9356 17978 9412 17980
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9238 17978
rect 9238 17926 9252 17978
rect 9276 17926 9290 17978
rect 9290 17926 9302 17978
rect 9302 17926 9332 17978
rect 9356 17926 9366 17978
rect 9366 17926 9412 17978
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 9276 17924 9332 17926
rect 9356 17924 9412 17926
rect 10046 18028 10048 18048
rect 10048 18028 10100 18048
rect 10100 18028 10102 18048
rect 10046 17992 10102 18028
rect 10046 17176 10102 17232
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 9276 16890 9332 16892
rect 9356 16890 9412 16892
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9238 16890
rect 9238 16838 9252 16890
rect 9276 16838 9290 16890
rect 9290 16838 9302 16890
rect 9302 16838 9332 16890
rect 9356 16838 9366 16890
rect 9366 16838 9412 16890
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 9276 16836 9332 16838
rect 9356 16836 9412 16838
rect 10046 16396 10048 16416
rect 10048 16396 10100 16416
rect 10100 16396 10102 16416
rect 10046 16360 10102 16396
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 9276 15802 9332 15804
rect 9356 15802 9412 15804
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9238 15802
rect 9238 15750 9252 15802
rect 9276 15750 9290 15802
rect 9290 15750 9302 15802
rect 9302 15750 9332 15802
rect 9356 15750 9366 15802
rect 9366 15750 9412 15802
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 9276 15748 9332 15750
rect 9356 15748 9412 15750
rect 10046 15680 10102 15736
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 9276 14714 9332 14716
rect 9356 14714 9412 14716
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9238 14714
rect 9238 14662 9252 14714
rect 9276 14662 9290 14714
rect 9290 14662 9302 14714
rect 9302 14662 9332 14714
rect 9356 14662 9366 14714
rect 9366 14662 9412 14714
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 9276 14660 9332 14662
rect 9356 14660 9412 14662
rect 10046 14884 10102 14920
rect 10046 14864 10048 14884
rect 10048 14864 10100 14884
rect 10100 14864 10102 14884
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 9276 13626 9332 13628
rect 9356 13626 9412 13628
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9238 13626
rect 9238 13574 9252 13626
rect 9276 13574 9290 13626
rect 9290 13574 9302 13626
rect 9302 13574 9332 13626
rect 9356 13574 9366 13626
rect 9366 13574 9412 13626
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 9276 13572 9332 13574
rect 9356 13572 9412 13574
rect 10046 14048 10102 14104
rect 9586 13368 9642 13424
rect 10046 12588 10048 12608
rect 10048 12588 10100 12608
rect 10100 12588 10102 12608
rect 10046 12552 10102 12588
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 9276 12538 9332 12540
rect 9356 12538 9412 12540
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9238 12538
rect 9238 12486 9252 12538
rect 9276 12486 9290 12538
rect 9290 12486 9302 12538
rect 9302 12486 9332 12538
rect 9356 12486 9366 12538
rect 9366 12486 9412 12538
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 9276 12484 9332 12486
rect 9356 12484 9412 12486
rect 10046 11736 10102 11792
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 9276 11450 9332 11452
rect 9356 11450 9412 11452
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9238 11450
rect 9238 11398 9252 11450
rect 9276 11398 9290 11450
rect 9290 11398 9302 11450
rect 9302 11398 9332 11450
rect 9356 11398 9366 11450
rect 9366 11398 9412 11450
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 9276 11396 9332 11398
rect 9356 11396 9412 11398
rect 10046 11056 10102 11112
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 9276 10362 9332 10364
rect 9356 10362 9412 10364
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9238 10362
rect 9238 10310 9252 10362
rect 9276 10310 9290 10362
rect 9290 10310 9302 10362
rect 9302 10310 9332 10362
rect 9356 10310 9366 10362
rect 9366 10310 9412 10362
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 9276 10308 9332 10310
rect 9356 10308 9412 10310
rect 10046 10240 10102 10296
rect 10046 9444 10102 9480
rect 10046 9424 10048 9444
rect 10048 9424 10100 9444
rect 10100 9424 10102 9444
rect 5852 9274 5908 9276
rect 5932 9274 5988 9276
rect 6012 9274 6068 9276
rect 6092 9274 6148 9276
rect 5852 9222 5898 9274
rect 5898 9222 5908 9274
rect 5932 9222 5962 9274
rect 5962 9222 5974 9274
rect 5974 9222 5988 9274
rect 6012 9222 6026 9274
rect 6026 9222 6038 9274
rect 6038 9222 6068 9274
rect 6092 9222 6102 9274
rect 6102 9222 6148 9274
rect 5852 9220 5908 9222
rect 5932 9220 5988 9222
rect 6012 9220 6068 9222
rect 6092 9220 6148 9222
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 9276 9274 9332 9276
rect 9356 9274 9412 9276
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9238 9274
rect 9238 9222 9252 9274
rect 9276 9222 9290 9274
rect 9290 9222 9302 9274
rect 9302 9222 9332 9274
rect 9356 9222 9366 9274
rect 9366 9222 9412 9274
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 9276 9220 9332 9222
rect 9356 9220 9412 9222
rect 10046 8780 10048 8800
rect 10048 8780 10100 8800
rect 10100 8780 10102 8800
rect 10046 8744 10102 8780
rect 7484 8730 7540 8732
rect 7564 8730 7620 8732
rect 7644 8730 7700 8732
rect 7724 8730 7780 8732
rect 7484 8678 7530 8730
rect 7530 8678 7540 8730
rect 7564 8678 7594 8730
rect 7594 8678 7606 8730
rect 7606 8678 7620 8730
rect 7644 8678 7658 8730
rect 7658 8678 7670 8730
rect 7670 8678 7700 8730
rect 7724 8678 7734 8730
rect 7734 8678 7780 8730
rect 7484 8676 7540 8678
rect 7564 8676 7620 8678
rect 7644 8676 7700 8678
rect 7724 8676 7780 8678
rect 5852 8186 5908 8188
rect 5932 8186 5988 8188
rect 6012 8186 6068 8188
rect 6092 8186 6148 8188
rect 5852 8134 5898 8186
rect 5898 8134 5908 8186
rect 5932 8134 5962 8186
rect 5962 8134 5974 8186
rect 5974 8134 5988 8186
rect 6012 8134 6026 8186
rect 6026 8134 6038 8186
rect 6038 8134 6068 8186
rect 6092 8134 6102 8186
rect 6102 8134 6148 8186
rect 5852 8132 5908 8134
rect 5932 8132 5988 8134
rect 6012 8132 6068 8134
rect 6092 8132 6148 8134
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 9276 8186 9332 8188
rect 9356 8186 9412 8188
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9238 8186
rect 9238 8134 9252 8186
rect 9276 8134 9290 8186
rect 9290 8134 9302 8186
rect 9302 8134 9332 8186
rect 9356 8134 9366 8186
rect 9366 8134 9412 8186
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 9276 8132 9332 8134
rect 9356 8132 9412 8134
rect 10046 7928 10102 7984
rect 7484 7642 7540 7644
rect 7564 7642 7620 7644
rect 7644 7642 7700 7644
rect 7724 7642 7780 7644
rect 7484 7590 7530 7642
rect 7530 7590 7540 7642
rect 7564 7590 7594 7642
rect 7594 7590 7606 7642
rect 7606 7590 7620 7642
rect 7644 7590 7658 7642
rect 7658 7590 7670 7642
rect 7670 7590 7700 7642
rect 7724 7590 7734 7642
rect 7734 7590 7780 7642
rect 7484 7588 7540 7590
rect 7564 7588 7620 7590
rect 7644 7588 7700 7590
rect 7724 7588 7780 7590
rect 10046 7148 10048 7168
rect 10048 7148 10100 7168
rect 10100 7148 10102 7168
rect 5852 7098 5908 7100
rect 5932 7098 5988 7100
rect 6012 7098 6068 7100
rect 6092 7098 6148 7100
rect 5852 7046 5898 7098
rect 5898 7046 5908 7098
rect 5932 7046 5962 7098
rect 5962 7046 5974 7098
rect 5974 7046 5988 7098
rect 6012 7046 6026 7098
rect 6026 7046 6038 7098
rect 6038 7046 6068 7098
rect 6092 7046 6102 7098
rect 6102 7046 6148 7098
rect 5852 7044 5908 7046
rect 5932 7044 5988 7046
rect 6012 7044 6068 7046
rect 6092 7044 6148 7046
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 9276 7098 9332 7100
rect 9356 7098 9412 7100
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9238 7098
rect 9238 7046 9252 7098
rect 9276 7046 9290 7098
rect 9290 7046 9302 7098
rect 9302 7046 9332 7098
rect 9356 7046 9366 7098
rect 9366 7046 9412 7098
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 9276 7044 9332 7046
rect 9356 7044 9412 7046
rect 10046 7112 10102 7148
rect 7484 6554 7540 6556
rect 7564 6554 7620 6556
rect 7644 6554 7700 6556
rect 7724 6554 7780 6556
rect 7484 6502 7530 6554
rect 7530 6502 7540 6554
rect 7564 6502 7594 6554
rect 7594 6502 7606 6554
rect 7606 6502 7620 6554
rect 7644 6502 7658 6554
rect 7658 6502 7670 6554
rect 7670 6502 7700 6554
rect 7724 6502 7734 6554
rect 7734 6502 7780 6554
rect 7484 6500 7540 6502
rect 7564 6500 7620 6502
rect 7644 6500 7700 6502
rect 7724 6500 7780 6502
rect 10046 6432 10102 6488
rect 5852 6010 5908 6012
rect 5932 6010 5988 6012
rect 6012 6010 6068 6012
rect 6092 6010 6148 6012
rect 5852 5958 5898 6010
rect 5898 5958 5908 6010
rect 5932 5958 5962 6010
rect 5962 5958 5974 6010
rect 5974 5958 5988 6010
rect 6012 5958 6026 6010
rect 6026 5958 6038 6010
rect 6038 5958 6068 6010
rect 6092 5958 6102 6010
rect 6102 5958 6148 6010
rect 5852 5956 5908 5958
rect 5932 5956 5988 5958
rect 6012 5956 6068 5958
rect 6092 5956 6148 5958
rect 7484 5466 7540 5468
rect 7564 5466 7620 5468
rect 7644 5466 7700 5468
rect 7724 5466 7780 5468
rect 7484 5414 7530 5466
rect 7530 5414 7540 5466
rect 7564 5414 7594 5466
rect 7594 5414 7606 5466
rect 7606 5414 7620 5466
rect 7644 5414 7658 5466
rect 7658 5414 7670 5466
rect 7670 5414 7700 5466
rect 7724 5414 7734 5466
rect 7734 5414 7780 5466
rect 7484 5412 7540 5414
rect 7564 5412 7620 5414
rect 7644 5412 7700 5414
rect 7724 5412 7780 5414
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 9276 6010 9332 6012
rect 9356 6010 9412 6012
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9238 6010
rect 9238 5958 9252 6010
rect 9276 5958 9290 6010
rect 9290 5958 9302 6010
rect 9302 5958 9332 6010
rect 9356 5958 9366 6010
rect 9366 5958 9412 6010
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 9276 5956 9332 5958
rect 9356 5956 9412 5958
rect 10046 5616 10102 5672
rect 5852 4922 5908 4924
rect 5932 4922 5988 4924
rect 6012 4922 6068 4924
rect 6092 4922 6148 4924
rect 5852 4870 5898 4922
rect 5898 4870 5908 4922
rect 5932 4870 5962 4922
rect 5962 4870 5974 4922
rect 5974 4870 5988 4922
rect 6012 4870 6026 4922
rect 6026 4870 6038 4922
rect 6038 4870 6068 4922
rect 6092 4870 6102 4922
rect 6102 4870 6148 4922
rect 5852 4868 5908 4870
rect 5932 4868 5988 4870
rect 6012 4868 6068 4870
rect 6092 4868 6148 4870
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 9276 4922 9332 4924
rect 9356 4922 9412 4924
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9238 4922
rect 9238 4870 9252 4922
rect 9276 4870 9290 4922
rect 9290 4870 9302 4922
rect 9302 4870 9332 4922
rect 9356 4870 9366 4922
rect 9366 4870 9412 4922
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 9276 4868 9332 4870
rect 9356 4868 9412 4870
rect 4066 4664 4122 4720
rect 10046 4800 10102 4856
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4266 4378
rect 4266 4326 4276 4378
rect 4300 4326 4330 4378
rect 4330 4326 4342 4378
rect 4342 4326 4356 4378
rect 4380 4326 4394 4378
rect 4394 4326 4406 4378
rect 4406 4326 4436 4378
rect 4460 4326 4470 4378
rect 4470 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 7484 4378 7540 4380
rect 7564 4378 7620 4380
rect 7644 4378 7700 4380
rect 7724 4378 7780 4380
rect 7484 4326 7530 4378
rect 7530 4326 7540 4378
rect 7564 4326 7594 4378
rect 7594 4326 7606 4378
rect 7606 4326 7620 4378
rect 7644 4326 7658 4378
rect 7658 4326 7670 4378
rect 7670 4326 7700 4378
rect 7724 4326 7734 4378
rect 7734 4326 7780 4378
rect 7484 4324 7540 4326
rect 7564 4324 7620 4326
rect 7644 4324 7700 4326
rect 7724 4324 7780 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4266 3290
rect 4266 3238 4276 3290
rect 4300 3238 4330 3290
rect 4330 3238 4342 3290
rect 4342 3238 4356 3290
rect 4380 3238 4394 3290
rect 4394 3238 4406 3290
rect 4406 3238 4436 3290
rect 4460 3238 4470 3290
rect 4470 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 5852 3834 5908 3836
rect 5932 3834 5988 3836
rect 6012 3834 6068 3836
rect 6092 3834 6148 3836
rect 5852 3782 5898 3834
rect 5898 3782 5908 3834
rect 5932 3782 5962 3834
rect 5962 3782 5974 3834
rect 5974 3782 5988 3834
rect 6012 3782 6026 3834
rect 6026 3782 6038 3834
rect 6038 3782 6068 3834
rect 6092 3782 6102 3834
rect 6102 3782 6148 3834
rect 5852 3780 5908 3782
rect 5932 3780 5988 3782
rect 6012 3780 6068 3782
rect 6092 3780 6148 3782
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 9276 3834 9332 3836
rect 9356 3834 9412 3836
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9238 3834
rect 9238 3782 9252 3834
rect 9276 3782 9290 3834
rect 9290 3782 9302 3834
rect 9302 3782 9332 3834
rect 9356 3782 9366 3834
rect 9366 3782 9412 3834
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 9276 3780 9332 3782
rect 9356 3780 9412 3782
rect 3514 2488 3570 2544
rect 10046 4120 10102 4176
rect 7484 3290 7540 3292
rect 7564 3290 7620 3292
rect 7644 3290 7700 3292
rect 7724 3290 7780 3292
rect 7484 3238 7530 3290
rect 7530 3238 7540 3290
rect 7564 3238 7594 3290
rect 7594 3238 7606 3290
rect 7606 3238 7620 3290
rect 7644 3238 7658 3290
rect 7658 3238 7670 3290
rect 7670 3238 7700 3290
rect 7724 3238 7734 3290
rect 7734 3238 7780 3290
rect 7484 3236 7540 3238
rect 7564 3236 7620 3238
rect 7644 3236 7700 3238
rect 7724 3236 7780 3238
rect 5852 2746 5908 2748
rect 5932 2746 5988 2748
rect 6012 2746 6068 2748
rect 6092 2746 6148 2748
rect 5852 2694 5898 2746
rect 5898 2694 5908 2746
rect 5932 2694 5962 2746
rect 5962 2694 5974 2746
rect 5974 2694 5988 2746
rect 6012 2694 6026 2746
rect 6026 2694 6038 2746
rect 6038 2694 6068 2746
rect 6092 2694 6102 2746
rect 6102 2694 6148 2746
rect 5852 2692 5908 2694
rect 5932 2692 5988 2694
rect 6012 2692 6068 2694
rect 6092 2692 6148 2694
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 9276 2746 9332 2748
rect 9356 2746 9412 2748
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9238 2746
rect 9238 2694 9252 2746
rect 9276 2694 9290 2746
rect 9290 2694 9302 2746
rect 9302 2694 9332 2746
rect 9356 2694 9366 2746
rect 9366 2694 9412 2746
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 9276 2692 9332 2694
rect 9356 2692 9412 2694
rect 2962 2216 3018 2272
rect 2870 1400 2926 1456
rect 2870 1028 2872 1048
rect 2872 1028 2924 1048
rect 2924 1028 2926 1048
rect 2870 992 2926 1028
rect 2778 584 2834 640
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4266 2202
rect 4266 2150 4276 2202
rect 4300 2150 4330 2202
rect 4330 2150 4342 2202
rect 4342 2150 4356 2202
rect 4380 2150 4394 2202
rect 4394 2150 4406 2202
rect 4406 2150 4436 2202
rect 4460 2150 4470 2202
rect 4470 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 7484 2202 7540 2204
rect 7564 2202 7620 2204
rect 7644 2202 7700 2204
rect 7724 2202 7780 2204
rect 7484 2150 7530 2202
rect 7530 2150 7540 2202
rect 7564 2150 7594 2202
rect 7594 2150 7606 2202
rect 7606 2150 7620 2202
rect 7644 2150 7658 2202
rect 7658 2150 7670 2202
rect 7670 2150 7700 2202
rect 7724 2150 7734 2202
rect 7734 2150 7780 2202
rect 7484 2148 7540 2150
rect 7564 2148 7620 2150
rect 7644 2148 7700 2150
rect 7724 2148 7780 2150
rect 10046 3340 10048 3360
rect 10048 3340 10100 3360
rect 10100 3340 10102 3360
rect 10046 3304 10102 3340
rect 10046 2488 10102 2544
rect 9494 1808 9550 1864
rect 9586 992 9642 1048
rect 9310 312 9366 368
rect 3974 176 4030 232
<< metal3 >>
rect 0 79568 800 79688
rect 9949 79522 10015 79525
rect 11200 79522 12000 79552
rect 9949 79520 12000 79522
rect 9949 79464 9954 79520
rect 10010 79464 12000 79520
rect 9949 79462 12000 79464
rect 9949 79459 10015 79462
rect 11200 79432 12000 79462
rect 0 79250 800 79280
rect 1393 79250 1459 79253
rect 0 79248 1459 79250
rect 0 79192 1398 79248
rect 1454 79192 1459 79248
rect 0 79190 1459 79192
rect 0 79160 800 79190
rect 1393 79187 1459 79190
rect 0 78842 800 78872
rect 1301 78842 1367 78845
rect 0 78840 1367 78842
rect 0 78784 1306 78840
rect 1362 78784 1367 78840
rect 0 78782 1367 78784
rect 0 78752 800 78782
rect 1301 78779 1367 78782
rect 9581 78706 9647 78709
rect 11200 78706 12000 78736
rect 9581 78704 12000 78706
rect 9581 78648 9586 78704
rect 9642 78648 12000 78704
rect 9581 78646 12000 78648
rect 9581 78643 9647 78646
rect 11200 78616 12000 78646
rect 0 78434 800 78464
rect 3877 78434 3943 78437
rect 0 78432 3943 78434
rect 0 78376 3882 78432
rect 3938 78376 3943 78432
rect 0 78374 3943 78376
rect 0 78344 800 78374
rect 3877 78371 3943 78374
rect 0 78026 800 78056
rect 4061 78026 4127 78029
rect 0 78024 4127 78026
rect 0 77968 4066 78024
rect 4122 77968 4127 78024
rect 0 77966 4127 77968
rect 0 77936 800 77966
rect 4061 77963 4127 77966
rect 9489 78026 9555 78029
rect 11200 78026 12000 78056
rect 9489 78024 12000 78026
rect 9489 77968 9494 78024
rect 9550 77968 12000 78024
rect 9489 77966 12000 77968
rect 9489 77963 9555 77966
rect 11200 77936 12000 77966
rect 2576 77824 2896 77825
rect 2576 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2576 77759 2896 77760
rect 5840 77824 6160 77825
rect 5840 77760 5848 77824
rect 5912 77760 5928 77824
rect 5992 77760 6008 77824
rect 6072 77760 6088 77824
rect 6152 77760 6160 77824
rect 5840 77759 6160 77760
rect 9104 77824 9424 77825
rect 9104 77760 9112 77824
rect 9176 77760 9192 77824
rect 9256 77760 9272 77824
rect 9336 77760 9352 77824
rect 9416 77760 9424 77824
rect 9104 77759 9424 77760
rect 0 77618 800 77648
rect 3601 77618 3667 77621
rect 0 77616 3667 77618
rect 0 77560 3606 77616
rect 3662 77560 3667 77616
rect 0 77558 3667 77560
rect 0 77528 800 77558
rect 3601 77555 3667 77558
rect 4208 77280 4528 77281
rect 0 77210 800 77240
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 77215 4528 77216
rect 7472 77280 7792 77281
rect 7472 77216 7480 77280
rect 7544 77216 7560 77280
rect 7624 77216 7640 77280
rect 7704 77216 7720 77280
rect 7784 77216 7792 77280
rect 7472 77215 7792 77216
rect 3969 77210 4035 77213
rect 0 77208 4035 77210
rect 0 77152 3974 77208
rect 4030 77152 4035 77208
rect 0 77150 4035 77152
rect 0 77120 800 77150
rect 3969 77147 4035 77150
rect 9397 77210 9463 77213
rect 11200 77210 12000 77240
rect 9397 77208 12000 77210
rect 9397 77152 9402 77208
rect 9458 77152 12000 77208
rect 9397 77150 12000 77152
rect 9397 77147 9463 77150
rect 11200 77120 12000 77150
rect 2865 76938 2931 76941
rect 1350 76936 2931 76938
rect 1350 76880 2870 76936
rect 2926 76880 2931 76936
rect 1350 76878 2931 76880
rect 0 76666 800 76696
rect 1350 76666 1410 76878
rect 2865 76875 2931 76878
rect 2576 76736 2896 76737
rect 2576 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2576 76671 2896 76672
rect 5840 76736 6160 76737
rect 5840 76672 5848 76736
rect 5912 76672 5928 76736
rect 5992 76672 6008 76736
rect 6072 76672 6088 76736
rect 6152 76672 6160 76736
rect 5840 76671 6160 76672
rect 9104 76736 9424 76737
rect 9104 76672 9112 76736
rect 9176 76672 9192 76736
rect 9256 76672 9272 76736
rect 9336 76672 9352 76736
rect 9416 76672 9424 76736
rect 9104 76671 9424 76672
rect 0 76606 1410 76666
rect 0 76576 800 76606
rect 10133 76394 10199 76397
rect 11200 76394 12000 76424
rect 10133 76392 12000 76394
rect 10133 76336 10138 76392
rect 10194 76336 12000 76392
rect 10133 76334 12000 76336
rect 10133 76331 10199 76334
rect 11200 76304 12000 76334
rect 0 76258 800 76288
rect 2957 76258 3023 76261
rect 0 76256 3023 76258
rect 0 76200 2962 76256
rect 3018 76200 3023 76256
rect 0 76198 3023 76200
rect 0 76168 800 76198
rect 2957 76195 3023 76198
rect 4208 76192 4528 76193
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 76127 4528 76128
rect 7472 76192 7792 76193
rect 7472 76128 7480 76192
rect 7544 76128 7560 76192
rect 7624 76128 7640 76192
rect 7704 76128 7720 76192
rect 7784 76128 7792 76192
rect 7472 76127 7792 76128
rect 0 75850 800 75880
rect 1485 75850 1551 75853
rect 0 75848 1551 75850
rect 0 75792 1490 75848
rect 1546 75792 1551 75848
rect 0 75790 1551 75792
rect 0 75760 800 75790
rect 1485 75787 1551 75790
rect 10133 75714 10199 75717
rect 11200 75714 12000 75744
rect 10133 75712 12000 75714
rect 10133 75656 10138 75712
rect 10194 75656 12000 75712
rect 10133 75654 12000 75656
rect 10133 75651 10199 75654
rect 2576 75648 2896 75649
rect 2576 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2576 75583 2896 75584
rect 5840 75648 6160 75649
rect 5840 75584 5848 75648
rect 5912 75584 5928 75648
rect 5992 75584 6008 75648
rect 6072 75584 6088 75648
rect 6152 75584 6160 75648
rect 5840 75583 6160 75584
rect 9104 75648 9424 75649
rect 9104 75584 9112 75648
rect 9176 75584 9192 75648
rect 9256 75584 9272 75648
rect 9336 75584 9352 75648
rect 9416 75584 9424 75648
rect 11200 75624 12000 75654
rect 9104 75583 9424 75584
rect 0 75442 800 75472
rect 3601 75442 3667 75445
rect 0 75440 3667 75442
rect 0 75384 3606 75440
rect 3662 75384 3667 75440
rect 0 75382 3667 75384
rect 0 75352 800 75382
rect 3601 75379 3667 75382
rect 4208 75104 4528 75105
rect 0 75034 800 75064
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 75039 4528 75040
rect 7472 75104 7792 75105
rect 7472 75040 7480 75104
rect 7544 75040 7560 75104
rect 7624 75040 7640 75104
rect 7704 75040 7720 75104
rect 7784 75040 7792 75104
rect 7472 75039 7792 75040
rect 3233 75034 3299 75037
rect 0 75032 3299 75034
rect 0 74976 3238 75032
rect 3294 74976 3299 75032
rect 0 74974 3299 74976
rect 0 74944 800 74974
rect 3233 74971 3299 74974
rect 10133 74898 10199 74901
rect 11200 74898 12000 74928
rect 10133 74896 12000 74898
rect 10133 74840 10138 74896
rect 10194 74840 12000 74896
rect 10133 74838 12000 74840
rect 10133 74835 10199 74838
rect 11200 74808 12000 74838
rect 1945 74762 2011 74765
rect 2078 74762 2084 74764
rect 1945 74760 2084 74762
rect 1945 74704 1950 74760
rect 2006 74704 2084 74760
rect 1945 74702 2084 74704
rect 1945 74699 2011 74702
rect 2078 74700 2084 74702
rect 2148 74700 2154 74764
rect 0 74626 800 74656
rect 1577 74626 1643 74629
rect 0 74624 1643 74626
rect 0 74568 1582 74624
rect 1638 74568 1643 74624
rect 0 74566 1643 74568
rect 0 74536 800 74566
rect 1577 74563 1643 74566
rect 2576 74560 2896 74561
rect 2576 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2576 74495 2896 74496
rect 5840 74560 6160 74561
rect 5840 74496 5848 74560
rect 5912 74496 5928 74560
rect 5992 74496 6008 74560
rect 6072 74496 6088 74560
rect 6152 74496 6160 74560
rect 5840 74495 6160 74496
rect 9104 74560 9424 74561
rect 9104 74496 9112 74560
rect 9176 74496 9192 74560
rect 9256 74496 9272 74560
rect 9336 74496 9352 74560
rect 9416 74496 9424 74560
rect 9104 74495 9424 74496
rect 0 74218 800 74248
rect 3233 74218 3299 74221
rect 0 74216 3299 74218
rect 0 74160 3238 74216
rect 3294 74160 3299 74216
rect 0 74158 3299 74160
rect 0 74128 800 74158
rect 3233 74155 3299 74158
rect 10133 74082 10199 74085
rect 11200 74082 12000 74112
rect 10133 74080 12000 74082
rect 10133 74024 10138 74080
rect 10194 74024 12000 74080
rect 10133 74022 12000 74024
rect 10133 74019 10199 74022
rect 4208 74016 4528 74017
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 73951 4528 73952
rect 7472 74016 7792 74017
rect 7472 73952 7480 74016
rect 7544 73952 7560 74016
rect 7624 73952 7640 74016
rect 7704 73952 7720 74016
rect 7784 73952 7792 74016
rect 11200 73992 12000 74022
rect 7472 73951 7792 73952
rect 0 73810 800 73840
rect 2957 73810 3023 73813
rect 0 73808 3023 73810
rect 0 73752 2962 73808
rect 3018 73752 3023 73808
rect 0 73750 3023 73752
rect 0 73720 800 73750
rect 2957 73747 3023 73750
rect 2576 73472 2896 73473
rect 2576 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2576 73407 2896 73408
rect 5840 73472 6160 73473
rect 5840 73408 5848 73472
rect 5912 73408 5928 73472
rect 5992 73408 6008 73472
rect 6072 73408 6088 73472
rect 6152 73408 6160 73472
rect 5840 73407 6160 73408
rect 9104 73472 9424 73473
rect 9104 73408 9112 73472
rect 9176 73408 9192 73472
rect 9256 73408 9272 73472
rect 9336 73408 9352 73472
rect 9416 73408 9424 73472
rect 9104 73407 9424 73408
rect 10133 73402 10199 73405
rect 11200 73402 12000 73432
rect 10133 73400 12000 73402
rect 10133 73344 10138 73400
rect 10194 73344 12000 73400
rect 10133 73342 12000 73344
rect 10133 73339 10199 73342
rect 11200 73312 12000 73342
rect 0 73266 800 73296
rect 2221 73266 2287 73269
rect 0 73264 2287 73266
rect 0 73208 2226 73264
rect 2282 73208 2287 73264
rect 0 73206 2287 73208
rect 0 73176 800 73206
rect 2221 73203 2287 73206
rect 4208 72928 4528 72929
rect 0 72858 800 72888
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 72863 4528 72864
rect 7472 72928 7792 72929
rect 7472 72864 7480 72928
rect 7544 72864 7560 72928
rect 7624 72864 7640 72928
rect 7704 72864 7720 72928
rect 7784 72864 7792 72928
rect 7472 72863 7792 72864
rect 1577 72858 1643 72861
rect 0 72856 1643 72858
rect 0 72800 1582 72856
rect 1638 72800 1643 72856
rect 0 72798 1643 72800
rect 0 72768 800 72798
rect 1577 72795 1643 72798
rect 1894 72660 1900 72724
rect 1964 72722 1970 72724
rect 2497 72722 2563 72725
rect 1964 72720 2563 72722
rect 1964 72664 2502 72720
rect 2558 72664 2563 72720
rect 1964 72662 2563 72664
rect 1964 72660 1970 72662
rect 2497 72659 2563 72662
rect 2865 72586 2931 72589
rect 1350 72584 2931 72586
rect 1350 72528 2870 72584
rect 2926 72528 2931 72584
rect 1350 72526 2931 72528
rect 0 72450 800 72480
rect 1350 72450 1410 72526
rect 2865 72523 2931 72526
rect 10133 72586 10199 72589
rect 11200 72586 12000 72616
rect 10133 72584 12000 72586
rect 10133 72528 10138 72584
rect 10194 72528 12000 72584
rect 10133 72526 12000 72528
rect 10133 72523 10199 72526
rect 11200 72496 12000 72526
rect 0 72390 1410 72450
rect 0 72360 800 72390
rect 2576 72384 2896 72385
rect 2576 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2576 72319 2896 72320
rect 5840 72384 6160 72385
rect 5840 72320 5848 72384
rect 5912 72320 5928 72384
rect 5992 72320 6008 72384
rect 6072 72320 6088 72384
rect 6152 72320 6160 72384
rect 5840 72319 6160 72320
rect 9104 72384 9424 72385
rect 9104 72320 9112 72384
rect 9176 72320 9192 72384
rect 9256 72320 9272 72384
rect 9336 72320 9352 72384
rect 9416 72320 9424 72384
rect 9104 72319 9424 72320
rect 1577 72180 1643 72181
rect 1526 72178 1532 72180
rect 1486 72118 1532 72178
rect 1596 72176 1643 72180
rect 1638 72120 1643 72176
rect 1526 72116 1532 72118
rect 1596 72116 1643 72120
rect 1577 72115 1643 72116
rect 0 72042 800 72072
rect 2221 72042 2287 72045
rect 0 72040 2287 72042
rect 0 71984 2226 72040
rect 2282 71984 2287 72040
rect 0 71982 2287 71984
rect 0 71952 800 71982
rect 2221 71979 2287 71982
rect 4208 71840 4528 71841
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 71775 4528 71776
rect 7472 71840 7792 71841
rect 7472 71776 7480 71840
rect 7544 71776 7560 71840
rect 7624 71776 7640 71840
rect 7704 71776 7720 71840
rect 7784 71776 7792 71840
rect 7472 71775 7792 71776
rect 10133 71770 10199 71773
rect 11200 71770 12000 71800
rect 10133 71768 12000 71770
rect 10133 71712 10138 71768
rect 10194 71712 12000 71768
rect 10133 71710 12000 71712
rect 10133 71707 10199 71710
rect 11200 71680 12000 71710
rect 0 71634 800 71664
rect 1393 71634 1459 71637
rect 0 71632 1459 71634
rect 0 71576 1398 71632
rect 1454 71576 1459 71632
rect 0 71574 1459 71576
rect 0 71544 800 71574
rect 1393 71571 1459 71574
rect 2576 71296 2896 71297
rect 0 71226 800 71256
rect 2576 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2576 71231 2896 71232
rect 5840 71296 6160 71297
rect 5840 71232 5848 71296
rect 5912 71232 5928 71296
rect 5992 71232 6008 71296
rect 6072 71232 6088 71296
rect 6152 71232 6160 71296
rect 5840 71231 6160 71232
rect 9104 71296 9424 71297
rect 9104 71232 9112 71296
rect 9176 71232 9192 71296
rect 9256 71232 9272 71296
rect 9336 71232 9352 71296
rect 9416 71232 9424 71296
rect 9104 71231 9424 71232
rect 1577 71226 1643 71229
rect 0 71224 1643 71226
rect 0 71168 1582 71224
rect 1638 71168 1643 71224
rect 0 71166 1643 71168
rect 0 71136 800 71166
rect 1577 71163 1643 71166
rect 10133 71090 10199 71093
rect 11200 71090 12000 71120
rect 10133 71088 12000 71090
rect 10133 71032 10138 71088
rect 10194 71032 12000 71088
rect 10133 71030 12000 71032
rect 10133 71027 10199 71030
rect 11200 71000 12000 71030
rect 0 70818 800 70848
rect 2221 70818 2287 70821
rect 0 70816 2287 70818
rect 0 70760 2226 70816
rect 2282 70760 2287 70816
rect 0 70758 2287 70760
rect 0 70728 800 70758
rect 2221 70755 2287 70758
rect 4208 70752 4528 70753
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 70687 4528 70688
rect 7472 70752 7792 70753
rect 7472 70688 7480 70752
rect 7544 70688 7560 70752
rect 7624 70688 7640 70752
rect 7704 70688 7720 70752
rect 7784 70688 7792 70752
rect 7472 70687 7792 70688
rect 1853 70682 1919 70685
rect 2262 70682 2268 70684
rect 1853 70680 2268 70682
rect 1853 70624 1858 70680
rect 1914 70624 2268 70680
rect 1853 70622 2268 70624
rect 1853 70619 1919 70622
rect 2262 70620 2268 70622
rect 2332 70620 2338 70684
rect 0 70410 800 70440
rect 933 70410 999 70413
rect 0 70408 999 70410
rect 0 70352 938 70408
rect 994 70352 999 70408
rect 0 70350 999 70352
rect 0 70320 800 70350
rect 933 70347 999 70350
rect 1485 70412 1551 70413
rect 1485 70408 1532 70412
rect 1596 70410 1602 70412
rect 1485 70352 1490 70408
rect 1485 70348 1532 70352
rect 1596 70350 1642 70410
rect 1596 70348 1602 70350
rect 1485 70347 1551 70348
rect 1945 70276 2011 70277
rect 2313 70276 2379 70277
rect 1894 70274 1900 70276
rect 1854 70214 1900 70274
rect 1964 70272 2011 70276
rect 2262 70274 2268 70276
rect 2006 70216 2011 70272
rect 1894 70212 1900 70214
rect 1964 70212 2011 70216
rect 2222 70214 2268 70274
rect 2332 70272 2379 70276
rect 2374 70216 2379 70272
rect 2262 70212 2268 70214
rect 2332 70212 2379 70216
rect 1945 70211 2011 70212
rect 2313 70211 2379 70212
rect 10133 70274 10199 70277
rect 11200 70274 12000 70304
rect 10133 70272 12000 70274
rect 10133 70216 10138 70272
rect 10194 70216 12000 70272
rect 10133 70214 12000 70216
rect 10133 70211 10199 70214
rect 2576 70208 2896 70209
rect 2576 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2576 70143 2896 70144
rect 5840 70208 6160 70209
rect 5840 70144 5848 70208
rect 5912 70144 5928 70208
rect 5992 70144 6008 70208
rect 6072 70144 6088 70208
rect 6152 70144 6160 70208
rect 5840 70143 6160 70144
rect 9104 70208 9424 70209
rect 9104 70144 9112 70208
rect 9176 70144 9192 70208
rect 9256 70144 9272 70208
rect 9336 70144 9352 70208
rect 9416 70144 9424 70208
rect 11200 70184 12000 70214
rect 9104 70143 9424 70144
rect 1761 70138 1827 70141
rect 2262 70138 2268 70140
rect 1761 70136 2268 70138
rect 1761 70080 1766 70136
rect 1822 70080 2268 70136
rect 1761 70078 2268 70080
rect 1761 70075 1827 70078
rect 2262 70076 2268 70078
rect 2332 70076 2338 70140
rect 1393 70004 1459 70005
rect 1342 69940 1348 70004
rect 1412 70002 1459 70004
rect 1412 70000 1504 70002
rect 1454 69944 1504 70000
rect 1412 69942 1504 69944
rect 1412 69940 1459 69942
rect 1393 69939 1459 69940
rect 0 69866 800 69896
rect 1577 69866 1643 69869
rect 0 69864 1643 69866
rect 0 69808 1582 69864
rect 1638 69808 1643 69864
rect 0 69806 1643 69808
rect 0 69776 800 69806
rect 1577 69803 1643 69806
rect 4208 69664 4528 69665
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 69599 4528 69600
rect 7472 69664 7792 69665
rect 7472 69600 7480 69664
rect 7544 69600 7560 69664
rect 7624 69600 7640 69664
rect 7704 69600 7720 69664
rect 7784 69600 7792 69664
rect 7472 69599 7792 69600
rect 0 69458 800 69488
rect 1669 69458 1735 69461
rect 0 69456 1735 69458
rect 0 69400 1674 69456
rect 1730 69400 1735 69456
rect 0 69398 1735 69400
rect 0 69368 800 69398
rect 1669 69395 1735 69398
rect 10133 69458 10199 69461
rect 11200 69458 12000 69488
rect 10133 69456 12000 69458
rect 10133 69400 10138 69456
rect 10194 69400 12000 69456
rect 10133 69398 12000 69400
rect 10133 69395 10199 69398
rect 11200 69368 12000 69398
rect 2576 69120 2896 69121
rect 0 69050 800 69080
rect 2576 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2576 69055 2896 69056
rect 5840 69120 6160 69121
rect 5840 69056 5848 69120
rect 5912 69056 5928 69120
rect 5992 69056 6008 69120
rect 6072 69056 6088 69120
rect 6152 69056 6160 69120
rect 5840 69055 6160 69056
rect 9104 69120 9424 69121
rect 9104 69056 9112 69120
rect 9176 69056 9192 69120
rect 9256 69056 9272 69120
rect 9336 69056 9352 69120
rect 9416 69056 9424 69120
rect 9104 69055 9424 69056
rect 2221 69050 2287 69053
rect 0 69048 2287 69050
rect 0 68992 2226 69048
rect 2282 68992 2287 69048
rect 0 68990 2287 68992
rect 0 68960 800 68990
rect 2221 68987 2287 68990
rect 10133 68778 10199 68781
rect 11200 68778 12000 68808
rect 10133 68776 12000 68778
rect 10133 68720 10138 68776
rect 10194 68720 12000 68776
rect 10133 68718 12000 68720
rect 10133 68715 10199 68718
rect 11200 68688 12000 68718
rect 0 68642 800 68672
rect 2773 68642 2839 68645
rect 0 68640 2839 68642
rect 0 68584 2778 68640
rect 2834 68584 2839 68640
rect 0 68582 2839 68584
rect 0 68552 800 68582
rect 2773 68579 2839 68582
rect 4208 68576 4528 68577
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 68511 4528 68512
rect 7472 68576 7792 68577
rect 7472 68512 7480 68576
rect 7544 68512 7560 68576
rect 7624 68512 7640 68576
rect 7704 68512 7720 68576
rect 7784 68512 7792 68576
rect 7472 68511 7792 68512
rect 0 68234 800 68264
rect 1577 68234 1643 68237
rect 0 68232 1643 68234
rect 0 68176 1582 68232
rect 1638 68176 1643 68232
rect 0 68174 1643 68176
rect 0 68144 800 68174
rect 1577 68171 1643 68174
rect 2576 68032 2896 68033
rect 2576 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2576 67967 2896 67968
rect 5840 68032 6160 68033
rect 5840 67968 5848 68032
rect 5912 67968 5928 68032
rect 5992 67968 6008 68032
rect 6072 67968 6088 68032
rect 6152 67968 6160 68032
rect 5840 67967 6160 67968
rect 9104 68032 9424 68033
rect 9104 67968 9112 68032
rect 9176 67968 9192 68032
rect 9256 67968 9272 68032
rect 9336 67968 9352 68032
rect 9416 67968 9424 68032
rect 9104 67967 9424 67968
rect 10133 67962 10199 67965
rect 11200 67962 12000 67992
rect 10133 67960 12000 67962
rect 10133 67904 10138 67960
rect 10194 67904 12000 67960
rect 10133 67902 12000 67904
rect 10133 67899 10199 67902
rect 11200 67872 12000 67902
rect 0 67826 800 67856
rect 2957 67826 3023 67829
rect 0 67824 3023 67826
rect 0 67768 2962 67824
rect 3018 67768 3023 67824
rect 0 67766 3023 67768
rect 0 67736 800 67766
rect 2957 67763 3023 67766
rect 2773 67690 2839 67693
rect 3325 67690 3391 67693
rect 2773 67688 3391 67690
rect 2773 67632 2778 67688
rect 2834 67632 3330 67688
rect 3386 67632 3391 67688
rect 2773 67630 3391 67632
rect 2773 67627 2839 67630
rect 3325 67627 3391 67630
rect 4208 67488 4528 67489
rect 0 67418 800 67448
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 67423 4528 67424
rect 7472 67488 7792 67489
rect 7472 67424 7480 67488
rect 7544 67424 7560 67488
rect 7624 67424 7640 67488
rect 7704 67424 7720 67488
rect 7784 67424 7792 67488
rect 7472 67423 7792 67424
rect 1577 67418 1643 67421
rect 0 67416 1643 67418
rect 0 67360 1582 67416
rect 1638 67360 1643 67416
rect 0 67358 1643 67360
rect 0 67328 800 67358
rect 1577 67355 1643 67358
rect 10133 67146 10199 67149
rect 11200 67146 12000 67176
rect 10133 67144 12000 67146
rect 10133 67088 10138 67144
rect 10194 67088 12000 67144
rect 10133 67086 12000 67088
rect 10133 67083 10199 67086
rect 11200 67056 12000 67086
rect 0 67010 800 67040
rect 1393 67010 1459 67013
rect 0 67008 1459 67010
rect 0 66952 1398 67008
rect 1454 66952 1459 67008
rect 0 66950 1459 66952
rect 0 66920 800 66950
rect 1393 66947 1459 66950
rect 2576 66944 2896 66945
rect 2576 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2576 66879 2896 66880
rect 5840 66944 6160 66945
rect 5840 66880 5848 66944
rect 5912 66880 5928 66944
rect 5992 66880 6008 66944
rect 6072 66880 6088 66944
rect 6152 66880 6160 66944
rect 5840 66879 6160 66880
rect 9104 66944 9424 66945
rect 9104 66880 9112 66944
rect 9176 66880 9192 66944
rect 9256 66880 9272 66944
rect 9336 66880 9352 66944
rect 9416 66880 9424 66944
rect 9104 66879 9424 66880
rect 0 66466 800 66496
rect 1393 66466 1459 66469
rect 0 66464 1459 66466
rect 0 66408 1398 66464
rect 1454 66408 1459 66464
rect 0 66406 1459 66408
rect 0 66376 800 66406
rect 1393 66403 1459 66406
rect 10133 66466 10199 66469
rect 11200 66466 12000 66496
rect 10133 66464 12000 66466
rect 10133 66408 10138 66464
rect 10194 66408 12000 66464
rect 10133 66406 12000 66408
rect 10133 66403 10199 66406
rect 4208 66400 4528 66401
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 66335 4528 66336
rect 7472 66400 7792 66401
rect 7472 66336 7480 66400
rect 7544 66336 7560 66400
rect 7624 66336 7640 66400
rect 7704 66336 7720 66400
rect 7784 66336 7792 66400
rect 11200 66376 12000 66406
rect 7472 66335 7792 66336
rect 1526 66268 1532 66332
rect 1596 66330 1602 66332
rect 1669 66330 1735 66333
rect 1596 66328 1735 66330
rect 1596 66272 1674 66328
rect 1730 66272 1735 66328
rect 1596 66270 1735 66272
rect 1596 66268 1602 66270
rect 1669 66267 1735 66270
rect 0 66058 800 66088
rect 1301 66058 1367 66061
rect 0 66056 1367 66058
rect 0 66000 1306 66056
rect 1362 66000 1367 66056
rect 0 65998 1367 66000
rect 0 65968 800 65998
rect 1301 65995 1367 65998
rect 2773 66058 2839 66061
rect 3734 66058 3740 66060
rect 2773 66056 3740 66058
rect 2773 66000 2778 66056
rect 2834 66000 3740 66056
rect 2773 65998 3740 66000
rect 2773 65995 2839 65998
rect 3734 65996 3740 65998
rect 3804 65996 3810 66060
rect 2576 65856 2896 65857
rect 2576 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2576 65791 2896 65792
rect 5840 65856 6160 65857
rect 5840 65792 5848 65856
rect 5912 65792 5928 65856
rect 5992 65792 6008 65856
rect 6072 65792 6088 65856
rect 6152 65792 6160 65856
rect 5840 65791 6160 65792
rect 9104 65856 9424 65857
rect 9104 65792 9112 65856
rect 9176 65792 9192 65856
rect 9256 65792 9272 65856
rect 9336 65792 9352 65856
rect 9416 65792 9424 65856
rect 9104 65791 9424 65792
rect 0 65650 800 65680
rect 1393 65650 1459 65653
rect 0 65648 1459 65650
rect 0 65592 1398 65648
rect 1454 65592 1459 65648
rect 0 65590 1459 65592
rect 0 65560 800 65590
rect 1393 65587 1459 65590
rect 10133 65650 10199 65653
rect 11200 65650 12000 65680
rect 10133 65648 12000 65650
rect 10133 65592 10138 65648
rect 10194 65592 12000 65648
rect 10133 65590 12000 65592
rect 10133 65587 10199 65590
rect 11200 65560 12000 65590
rect 4208 65312 4528 65313
rect 0 65242 800 65272
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 65247 4528 65248
rect 7472 65312 7792 65313
rect 7472 65248 7480 65312
rect 7544 65248 7560 65312
rect 7624 65248 7640 65312
rect 7704 65248 7720 65312
rect 7784 65248 7792 65312
rect 7472 65247 7792 65248
rect 3969 65242 4035 65245
rect 0 65240 4035 65242
rect 0 65184 3974 65240
rect 4030 65184 4035 65240
rect 0 65182 4035 65184
rect 0 65152 800 65182
rect 3969 65179 4035 65182
rect 1393 65106 1459 65109
rect 1577 65106 1643 65109
rect 1393 65104 1643 65106
rect 1393 65048 1398 65104
rect 1454 65048 1582 65104
rect 1638 65048 1643 65104
rect 1393 65046 1643 65048
rect 1393 65043 1459 65046
rect 1577 65043 1643 65046
rect 3049 65106 3115 65109
rect 3550 65106 3556 65108
rect 3049 65104 3556 65106
rect 3049 65048 3054 65104
rect 3110 65048 3556 65104
rect 3049 65046 3556 65048
rect 3049 65043 3115 65046
rect 3550 65044 3556 65046
rect 3620 65044 3626 65108
rect 1669 64972 1735 64973
rect 1669 64968 1716 64972
rect 1780 64970 1786 64972
rect 1669 64912 1674 64968
rect 1669 64908 1716 64912
rect 1780 64910 1826 64970
rect 1780 64908 1786 64910
rect 1669 64907 1735 64908
rect 0 64834 800 64864
rect 3325 64834 3391 64837
rect 0 64774 1410 64834
rect 0 64744 800 64774
rect 1350 64562 1410 64774
rect 3190 64832 3391 64834
rect 3190 64776 3330 64832
rect 3386 64776 3391 64832
rect 3190 64774 3391 64776
rect 2576 64768 2896 64769
rect 2576 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2576 64703 2896 64704
rect 3190 64562 3250 64774
rect 3325 64771 3391 64774
rect 10133 64834 10199 64837
rect 11200 64834 12000 64864
rect 10133 64832 12000 64834
rect 10133 64776 10138 64832
rect 10194 64776 12000 64832
rect 10133 64774 12000 64776
rect 10133 64771 10199 64774
rect 5840 64768 6160 64769
rect 5840 64704 5848 64768
rect 5912 64704 5928 64768
rect 5992 64704 6008 64768
rect 6072 64704 6088 64768
rect 6152 64704 6160 64768
rect 5840 64703 6160 64704
rect 9104 64768 9424 64769
rect 9104 64704 9112 64768
rect 9176 64704 9192 64768
rect 9256 64704 9272 64768
rect 9336 64704 9352 64768
rect 9416 64704 9424 64768
rect 11200 64744 12000 64774
rect 9104 64703 9424 64704
rect 1350 64502 3250 64562
rect 0 64426 800 64456
rect 3049 64426 3115 64429
rect 0 64424 3115 64426
rect 0 64368 3054 64424
rect 3110 64368 3115 64424
rect 0 64366 3115 64368
rect 0 64336 800 64366
rect 3049 64363 3115 64366
rect 4208 64224 4528 64225
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 64159 4528 64160
rect 7472 64224 7792 64225
rect 7472 64160 7480 64224
rect 7544 64160 7560 64224
rect 7624 64160 7640 64224
rect 7704 64160 7720 64224
rect 7784 64160 7792 64224
rect 7472 64159 7792 64160
rect 10133 64154 10199 64157
rect 11200 64154 12000 64184
rect 10133 64152 12000 64154
rect 10133 64096 10138 64152
rect 10194 64096 12000 64152
rect 10133 64094 12000 64096
rect 10133 64091 10199 64094
rect 11200 64064 12000 64094
rect 0 64018 800 64048
rect 3141 64018 3207 64021
rect 0 64016 3207 64018
rect 0 63960 3146 64016
rect 3202 63960 3207 64016
rect 0 63958 3207 63960
rect 0 63928 800 63958
rect 3141 63955 3207 63958
rect 2497 63882 2563 63885
rect 2998 63882 3004 63884
rect 2497 63880 3004 63882
rect 2497 63824 2502 63880
rect 2558 63824 3004 63880
rect 2497 63822 3004 63824
rect 2497 63819 2563 63822
rect 2998 63820 3004 63822
rect 3068 63820 3074 63884
rect 2576 63680 2896 63681
rect 0 63610 800 63640
rect 2576 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2576 63615 2896 63616
rect 5840 63680 6160 63681
rect 5840 63616 5848 63680
rect 5912 63616 5928 63680
rect 5992 63616 6008 63680
rect 6072 63616 6088 63680
rect 6152 63616 6160 63680
rect 5840 63615 6160 63616
rect 9104 63680 9424 63681
rect 9104 63616 9112 63680
rect 9176 63616 9192 63680
rect 9256 63616 9272 63680
rect 9336 63616 9352 63680
rect 9416 63616 9424 63680
rect 9104 63615 9424 63616
rect 1577 63610 1643 63613
rect 0 63608 1643 63610
rect 0 63552 1582 63608
rect 1638 63552 1643 63608
rect 0 63550 1643 63552
rect 0 63520 800 63550
rect 1577 63547 1643 63550
rect 3049 63608 3115 63613
rect 3049 63552 3054 63608
rect 3110 63552 3115 63608
rect 3049 63547 3115 63552
rect 2865 63474 2931 63477
rect 3052 63474 3112 63547
rect 2865 63472 3112 63474
rect 2865 63416 2870 63472
rect 2926 63416 3112 63472
rect 2865 63414 3112 63416
rect 2865 63411 2931 63414
rect 9305 63338 9371 63341
rect 11200 63338 12000 63368
rect 9305 63336 12000 63338
rect 9305 63280 9310 63336
rect 9366 63280 12000 63336
rect 9305 63278 12000 63280
rect 9305 63275 9371 63278
rect 11200 63248 12000 63278
rect 4208 63136 4528 63137
rect 0 63066 800 63096
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 63071 4528 63072
rect 7472 63136 7792 63137
rect 7472 63072 7480 63136
rect 7544 63072 7560 63136
rect 7624 63072 7640 63136
rect 7704 63072 7720 63136
rect 7784 63072 7792 63136
rect 7472 63071 7792 63072
rect 3325 63066 3391 63069
rect 0 63064 3391 63066
rect 0 63008 3330 63064
rect 3386 63008 3391 63064
rect 0 63006 3391 63008
rect 0 62976 800 63006
rect 3325 63003 3391 63006
rect 2262 62868 2268 62932
rect 2332 62930 2338 62932
rect 2589 62930 2655 62933
rect 2332 62928 2655 62930
rect 2332 62872 2594 62928
rect 2650 62872 2655 62928
rect 2332 62870 2655 62872
rect 2332 62868 2338 62870
rect 2589 62867 2655 62870
rect 3693 62794 3759 62797
rect 1350 62792 3759 62794
rect 1350 62736 3698 62792
rect 3754 62736 3759 62792
rect 1350 62734 3759 62736
rect 0 62658 800 62688
rect 1350 62658 1410 62734
rect 3693 62731 3759 62734
rect 0 62598 1410 62658
rect 1669 62658 1735 62661
rect 1894 62658 1900 62660
rect 1669 62656 1900 62658
rect 1669 62600 1674 62656
rect 1730 62600 1900 62656
rect 1669 62598 1900 62600
rect 0 62568 800 62598
rect 1669 62595 1735 62598
rect 1894 62596 1900 62598
rect 1964 62596 1970 62660
rect 3693 62658 3759 62661
rect 3969 62658 4035 62661
rect 3693 62656 4035 62658
rect 3693 62600 3698 62656
rect 3754 62600 3974 62656
rect 4030 62600 4035 62656
rect 3693 62598 4035 62600
rect 3693 62595 3759 62598
rect 3969 62595 4035 62598
rect 2576 62592 2896 62593
rect 2576 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2576 62527 2896 62528
rect 5840 62592 6160 62593
rect 5840 62528 5848 62592
rect 5912 62528 5928 62592
rect 5992 62528 6008 62592
rect 6072 62528 6088 62592
rect 6152 62528 6160 62592
rect 5840 62527 6160 62528
rect 9104 62592 9424 62593
rect 9104 62528 9112 62592
rect 9176 62528 9192 62592
rect 9256 62528 9272 62592
rect 9336 62528 9352 62592
rect 9416 62528 9424 62592
rect 9104 62527 9424 62528
rect 10133 62522 10199 62525
rect 11200 62522 12000 62552
rect 10133 62520 12000 62522
rect 10133 62464 10138 62520
rect 10194 62464 12000 62520
rect 10133 62462 12000 62464
rect 10133 62459 10199 62462
rect 11200 62432 12000 62462
rect 0 62250 800 62280
rect 2773 62250 2839 62253
rect 0 62248 2839 62250
rect 0 62192 2778 62248
rect 2834 62192 2839 62248
rect 0 62190 2839 62192
rect 0 62160 800 62190
rect 2773 62187 2839 62190
rect 4208 62048 4528 62049
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 61983 4528 61984
rect 7472 62048 7792 62049
rect 7472 61984 7480 62048
rect 7544 61984 7560 62048
rect 7624 61984 7640 62048
rect 7704 61984 7720 62048
rect 7784 61984 7792 62048
rect 7472 61983 7792 61984
rect 0 61842 800 61872
rect 2313 61842 2379 61845
rect 0 61840 2379 61842
rect 0 61784 2318 61840
rect 2374 61784 2379 61840
rect 0 61782 2379 61784
rect 0 61752 800 61782
rect 2313 61779 2379 61782
rect 10133 61842 10199 61845
rect 11200 61842 12000 61872
rect 10133 61840 12000 61842
rect 10133 61784 10138 61840
rect 10194 61784 12000 61840
rect 10133 61782 12000 61784
rect 10133 61779 10199 61782
rect 11200 61752 12000 61782
rect 2589 61706 2655 61709
rect 3182 61706 3188 61708
rect 2589 61704 3188 61706
rect 2589 61648 2594 61704
rect 2650 61648 3188 61704
rect 2589 61646 3188 61648
rect 2589 61643 2655 61646
rect 3182 61644 3188 61646
rect 3252 61644 3258 61708
rect 2576 61504 2896 61505
rect 0 61434 800 61464
rect 2576 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2576 61439 2896 61440
rect 5840 61504 6160 61505
rect 5840 61440 5848 61504
rect 5912 61440 5928 61504
rect 5992 61440 6008 61504
rect 6072 61440 6088 61504
rect 6152 61440 6160 61504
rect 5840 61439 6160 61440
rect 9104 61504 9424 61505
rect 9104 61440 9112 61504
rect 9176 61440 9192 61504
rect 9256 61440 9272 61504
rect 9336 61440 9352 61504
rect 9416 61440 9424 61504
rect 9104 61439 9424 61440
rect 1577 61434 1643 61437
rect 0 61432 1643 61434
rect 0 61376 1582 61432
rect 1638 61376 1643 61432
rect 0 61374 1643 61376
rect 0 61344 800 61374
rect 1577 61371 1643 61374
rect 2129 61162 2195 61165
rect 2262 61162 2268 61164
rect 2129 61160 2268 61162
rect 2129 61104 2134 61160
rect 2190 61104 2268 61160
rect 2129 61102 2268 61104
rect 2129 61099 2195 61102
rect 2262 61100 2268 61102
rect 2332 61100 2338 61164
rect 0 61026 800 61056
rect 2313 61026 2379 61029
rect 0 61024 2379 61026
rect 0 60968 2318 61024
rect 2374 60968 2379 61024
rect 0 60966 2379 60968
rect 0 60936 800 60966
rect 2313 60963 2379 60966
rect 10133 61026 10199 61029
rect 11200 61026 12000 61056
rect 10133 61024 12000 61026
rect 10133 60968 10138 61024
rect 10194 60968 12000 61024
rect 10133 60966 12000 60968
rect 10133 60963 10199 60966
rect 4208 60960 4528 60961
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 60895 4528 60896
rect 7472 60960 7792 60961
rect 7472 60896 7480 60960
rect 7544 60896 7560 60960
rect 7624 60896 7640 60960
rect 7704 60896 7720 60960
rect 7784 60896 7792 60960
rect 11200 60936 12000 60966
rect 7472 60895 7792 60896
rect 2313 60890 2379 60893
rect 3969 60892 4035 60893
rect 3182 60890 3188 60892
rect 2313 60888 3188 60890
rect 2313 60832 2318 60888
rect 2374 60832 3188 60888
rect 2313 60830 3188 60832
rect 2313 60827 2379 60830
rect 3182 60828 3188 60830
rect 3252 60828 3258 60892
rect 3918 60828 3924 60892
rect 3988 60890 4035 60892
rect 3988 60888 4080 60890
rect 4030 60832 4080 60888
rect 3988 60830 4080 60832
rect 3988 60828 4035 60830
rect 3969 60827 4035 60828
rect 3049 60754 3115 60757
rect 3969 60754 4035 60757
rect 3049 60752 4035 60754
rect 3049 60696 3054 60752
rect 3110 60696 3974 60752
rect 4030 60696 4035 60752
rect 3049 60694 4035 60696
rect 3049 60691 3115 60694
rect 3969 60691 4035 60694
rect 0 60618 800 60648
rect 2773 60618 2839 60621
rect 3969 60620 4035 60621
rect 3918 60618 3924 60620
rect 0 60616 2839 60618
rect 0 60560 2778 60616
rect 2834 60560 2839 60616
rect 0 60558 2839 60560
rect 3878 60558 3924 60618
rect 3988 60616 4035 60620
rect 4030 60560 4035 60616
rect 0 60528 800 60558
rect 2773 60555 2839 60558
rect 3918 60556 3924 60558
rect 3988 60556 4035 60560
rect 3969 60555 4035 60556
rect 1945 60482 2011 60485
rect 2262 60482 2268 60484
rect 1945 60480 2268 60482
rect 1945 60424 1950 60480
rect 2006 60424 2268 60480
rect 1945 60422 2268 60424
rect 1945 60419 2011 60422
rect 2262 60420 2268 60422
rect 2332 60420 2338 60484
rect 2576 60416 2896 60417
rect 2576 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2576 60351 2896 60352
rect 5840 60416 6160 60417
rect 5840 60352 5848 60416
rect 5912 60352 5928 60416
rect 5992 60352 6008 60416
rect 6072 60352 6088 60416
rect 6152 60352 6160 60416
rect 5840 60351 6160 60352
rect 9104 60416 9424 60417
rect 9104 60352 9112 60416
rect 9176 60352 9192 60416
rect 9256 60352 9272 60416
rect 9336 60352 9352 60416
rect 9416 60352 9424 60416
rect 9104 60351 9424 60352
rect 1342 60284 1348 60348
rect 1412 60346 1418 60348
rect 2262 60346 2268 60348
rect 1412 60286 2268 60346
rect 1412 60284 1418 60286
rect 2262 60284 2268 60286
rect 2332 60284 2338 60348
rect 10133 60346 10199 60349
rect 11200 60346 12000 60376
rect 10133 60344 12000 60346
rect 10133 60288 10138 60344
rect 10194 60288 12000 60344
rect 10133 60286 12000 60288
rect 10133 60283 10199 60286
rect 11200 60256 12000 60286
rect 0 60210 800 60240
rect 1577 60210 1643 60213
rect 0 60208 1643 60210
rect 0 60152 1582 60208
rect 1638 60152 1643 60208
rect 0 60150 1643 60152
rect 0 60120 800 60150
rect 1577 60147 1643 60150
rect 2078 60148 2084 60212
rect 2148 60210 2154 60212
rect 2497 60210 2563 60213
rect 2148 60208 2563 60210
rect 2148 60152 2502 60208
rect 2558 60152 2563 60208
rect 2148 60150 2563 60152
rect 2148 60148 2154 60150
rect 2497 60147 2563 60150
rect 2078 60012 2084 60076
rect 2148 60074 2154 60076
rect 2589 60074 2655 60077
rect 2148 60072 2655 60074
rect 2148 60016 2594 60072
rect 2650 60016 2655 60072
rect 2148 60014 2655 60016
rect 2148 60012 2154 60014
rect 2589 60011 2655 60014
rect 473 59938 539 59941
rect 3366 59938 3372 59940
rect 473 59936 3372 59938
rect 473 59880 478 59936
rect 534 59880 3372 59936
rect 473 59878 3372 59880
rect 473 59875 539 59878
rect 3366 59876 3372 59878
rect 3436 59876 3442 59940
rect 4208 59872 4528 59873
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 59807 4528 59808
rect 7472 59872 7792 59873
rect 7472 59808 7480 59872
rect 7544 59808 7560 59872
rect 7624 59808 7640 59872
rect 7704 59808 7720 59872
rect 7784 59808 7792 59872
rect 7472 59807 7792 59808
rect 0 59666 800 59696
rect 2313 59666 2379 59669
rect 0 59664 2379 59666
rect 0 59608 2318 59664
rect 2374 59608 2379 59664
rect 0 59606 2379 59608
rect 0 59576 800 59606
rect 2313 59603 2379 59606
rect 9305 59530 9371 59533
rect 11200 59530 12000 59560
rect 9305 59528 12000 59530
rect 9305 59472 9310 59528
rect 9366 59472 12000 59528
rect 9305 59470 12000 59472
rect 9305 59467 9371 59470
rect 11200 59440 12000 59470
rect 2576 59328 2896 59329
rect 0 59258 800 59288
rect 2576 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2576 59263 2896 59264
rect 5840 59328 6160 59329
rect 5840 59264 5848 59328
rect 5912 59264 5928 59328
rect 5992 59264 6008 59328
rect 6072 59264 6088 59328
rect 6152 59264 6160 59328
rect 5840 59263 6160 59264
rect 9104 59328 9424 59329
rect 9104 59264 9112 59328
rect 9176 59264 9192 59328
rect 9256 59264 9272 59328
rect 9336 59264 9352 59328
rect 9416 59264 9424 59328
rect 9104 59263 9424 59264
rect 1577 59258 1643 59261
rect 3550 59258 3556 59260
rect 0 59256 1643 59258
rect 0 59200 1582 59256
rect 1638 59200 1643 59256
rect 0 59198 1643 59200
rect 0 59168 800 59198
rect 1577 59195 1643 59198
rect 3006 59198 3556 59258
rect 2681 59122 2747 59125
rect 3006 59122 3066 59198
rect 3550 59196 3556 59198
rect 3620 59196 3626 59260
rect 2681 59120 3066 59122
rect 2681 59064 2686 59120
rect 2742 59064 3066 59120
rect 2681 59062 3066 59064
rect 3141 59122 3207 59125
rect 3550 59122 3556 59124
rect 3141 59120 3556 59122
rect 3141 59064 3146 59120
rect 3202 59064 3556 59120
rect 3141 59062 3556 59064
rect 2681 59059 2747 59062
rect 3141 59059 3207 59062
rect 3550 59060 3556 59062
rect 3620 59060 3626 59124
rect 0 58850 800 58880
rect 3049 58850 3115 58853
rect 0 58848 3115 58850
rect 0 58792 3054 58848
rect 3110 58792 3115 58848
rect 0 58790 3115 58792
rect 0 58760 800 58790
rect 3049 58787 3115 58790
rect 4208 58784 4528 58785
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 58719 4528 58720
rect 7472 58784 7792 58785
rect 7472 58720 7480 58784
rect 7544 58720 7560 58784
rect 7624 58720 7640 58784
rect 7704 58720 7720 58784
rect 7784 58720 7792 58784
rect 7472 58719 7792 58720
rect 10133 58714 10199 58717
rect 11200 58714 12000 58744
rect 10133 58712 12000 58714
rect 10133 58656 10138 58712
rect 10194 58656 12000 58712
rect 10133 58654 12000 58656
rect 10133 58651 10199 58654
rect 11200 58624 12000 58654
rect 0 58442 800 58472
rect 2313 58442 2379 58445
rect 2681 58442 2747 58445
rect 3182 58442 3188 58444
rect 0 58440 2379 58442
rect 0 58384 2318 58440
rect 2374 58384 2379 58440
rect 0 58382 2379 58384
rect 0 58352 800 58382
rect 2313 58379 2379 58382
rect 2454 58440 3188 58442
rect 2454 58384 2686 58440
rect 2742 58384 3188 58440
rect 2454 58382 3188 58384
rect 2313 58306 2379 58309
rect 2454 58306 2514 58382
rect 2681 58379 2747 58382
rect 3182 58380 3188 58382
rect 3252 58380 3258 58444
rect 2313 58304 2514 58306
rect 2313 58248 2318 58304
rect 2374 58248 2514 58304
rect 2313 58246 2514 58248
rect 2313 58243 2379 58246
rect 2576 58240 2896 58241
rect 2576 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2576 58175 2896 58176
rect 5840 58240 6160 58241
rect 5840 58176 5848 58240
rect 5912 58176 5928 58240
rect 5992 58176 6008 58240
rect 6072 58176 6088 58240
rect 6152 58176 6160 58240
rect 5840 58175 6160 58176
rect 9104 58240 9424 58241
rect 9104 58176 9112 58240
rect 9176 58176 9192 58240
rect 9256 58176 9272 58240
rect 9336 58176 9352 58240
rect 9416 58176 9424 58240
rect 9104 58175 9424 58176
rect 0 58034 800 58064
rect 1393 58034 1459 58037
rect 0 58032 1459 58034
rect 0 57976 1398 58032
rect 1454 57976 1459 58032
rect 0 57974 1459 57976
rect 0 57944 800 57974
rect 1393 57971 1459 57974
rect 2078 57972 2084 58036
rect 2148 58034 2154 58036
rect 2589 58034 2655 58037
rect 2148 58032 2655 58034
rect 2148 57976 2594 58032
rect 2650 57976 2655 58032
rect 2148 57974 2655 57976
rect 2148 57972 2154 57974
rect 2589 57971 2655 57974
rect 2773 58034 2839 58037
rect 3734 58034 3740 58036
rect 2773 58032 3740 58034
rect 2773 57976 2778 58032
rect 2834 57976 3740 58032
rect 2773 57974 3740 57976
rect 2773 57971 2839 57974
rect 3734 57972 3740 57974
rect 3804 57972 3810 58036
rect 10133 58034 10199 58037
rect 11200 58034 12000 58064
rect 10133 58032 12000 58034
rect 10133 57976 10138 58032
rect 10194 57976 12000 58032
rect 10133 57974 12000 57976
rect 10133 57971 10199 57974
rect 11200 57944 12000 57974
rect 974 57836 980 57900
rect 1044 57898 1050 57900
rect 1853 57898 1919 57901
rect 1044 57896 1919 57898
rect 1044 57840 1858 57896
rect 1914 57840 1919 57896
rect 1044 57838 1919 57840
rect 1044 57836 1050 57838
rect 1853 57835 1919 57838
rect 1158 57700 1164 57764
rect 1228 57762 1234 57764
rect 2405 57762 2471 57765
rect 1228 57760 2471 57762
rect 1228 57704 2410 57760
rect 2466 57704 2471 57760
rect 1228 57702 2471 57704
rect 1228 57700 1234 57702
rect 2405 57699 2471 57702
rect 3049 57762 3115 57765
rect 3734 57762 3740 57764
rect 3049 57760 3740 57762
rect 3049 57704 3054 57760
rect 3110 57704 3740 57760
rect 3049 57702 3740 57704
rect 3049 57699 3115 57702
rect 3734 57700 3740 57702
rect 3804 57700 3810 57764
rect 4208 57696 4528 57697
rect 0 57626 800 57656
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 57631 4528 57632
rect 7472 57696 7792 57697
rect 7472 57632 7480 57696
rect 7544 57632 7560 57696
rect 7624 57632 7640 57696
rect 7704 57632 7720 57696
rect 7784 57632 7792 57696
rect 7472 57631 7792 57632
rect 1577 57626 1643 57629
rect 0 57624 1643 57626
rect 0 57568 1582 57624
rect 1638 57568 1643 57624
rect 0 57566 1643 57568
rect 0 57536 800 57566
rect 1577 57563 1643 57566
rect 2078 57564 2084 57628
rect 2148 57626 2154 57628
rect 2681 57626 2747 57629
rect 2148 57624 2747 57626
rect 2148 57568 2686 57624
rect 2742 57568 2747 57624
rect 2148 57566 2747 57568
rect 2148 57564 2154 57566
rect 2681 57563 2747 57566
rect 3141 57628 3207 57629
rect 3141 57624 3188 57628
rect 3252 57626 3258 57628
rect 3141 57568 3146 57624
rect 3141 57564 3188 57568
rect 3252 57566 3298 57626
rect 3252 57564 3258 57566
rect 3141 57563 3207 57564
rect 1342 57428 1348 57492
rect 1412 57490 1418 57492
rect 1577 57490 1643 57493
rect 6913 57490 6979 57493
rect 1412 57488 1643 57490
rect 1412 57432 1582 57488
rect 1638 57432 1643 57488
rect 1412 57430 1643 57432
rect 1412 57428 1418 57430
rect 1577 57427 1643 57430
rect 1856 57488 6979 57490
rect 1856 57432 6918 57488
rect 6974 57432 6979 57488
rect 1856 57430 6979 57432
rect 1485 57354 1551 57357
rect 1856 57354 1916 57430
rect 6913 57427 6979 57430
rect 2589 57354 2655 57357
rect 1485 57352 1916 57354
rect 1485 57296 1490 57352
rect 1546 57296 1916 57352
rect 1485 57294 1916 57296
rect 2454 57352 2655 57354
rect 2454 57296 2594 57352
rect 2650 57296 2655 57352
rect 2454 57294 2655 57296
rect 1485 57291 1551 57294
rect 0 57218 800 57248
rect 1158 57218 1164 57220
rect 0 57158 1164 57218
rect 0 57128 800 57158
rect 1158 57156 1164 57158
rect 1228 57156 1234 57220
rect 1342 57020 1348 57084
rect 1412 57082 1418 57084
rect 1761 57082 1827 57085
rect 1412 57080 1827 57082
rect 1412 57024 1766 57080
rect 1822 57024 1827 57080
rect 1412 57022 1827 57024
rect 1412 57020 1418 57022
rect 1761 57019 1827 57022
rect 2454 56949 2514 57294
rect 2589 57291 2655 57294
rect 3049 57354 3115 57357
rect 5574 57354 5580 57356
rect 3049 57352 5580 57354
rect 3049 57296 3054 57352
rect 3110 57296 5580 57352
rect 3049 57294 5580 57296
rect 3049 57291 3115 57294
rect 5574 57292 5580 57294
rect 5644 57292 5650 57356
rect 9489 57218 9555 57221
rect 11200 57218 12000 57248
rect 9489 57216 12000 57218
rect 9489 57160 9494 57216
rect 9550 57160 12000 57216
rect 9489 57158 12000 57160
rect 9489 57155 9555 57158
rect 2576 57152 2896 57153
rect 2576 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2576 57087 2896 57088
rect 5840 57152 6160 57153
rect 5840 57088 5848 57152
rect 5912 57088 5928 57152
rect 5992 57088 6008 57152
rect 6072 57088 6088 57152
rect 6152 57088 6160 57152
rect 5840 57087 6160 57088
rect 9104 57152 9424 57153
rect 9104 57088 9112 57152
rect 9176 57088 9192 57152
rect 9256 57088 9272 57152
rect 9336 57088 9352 57152
rect 9416 57088 9424 57152
rect 11200 57128 12000 57158
rect 9104 57087 9424 57088
rect 657 56946 723 56949
rect 790 56946 796 56948
rect 657 56944 796 56946
rect 657 56888 662 56944
rect 718 56888 796 56944
rect 657 56886 796 56888
rect 657 56883 723 56886
rect 790 56884 796 56886
rect 860 56884 866 56948
rect 2454 56944 2563 56949
rect 2454 56888 2502 56944
rect 2558 56888 2563 56944
rect 2454 56886 2563 56888
rect 2497 56883 2563 56886
rect 1209 56812 1275 56813
rect 1158 56748 1164 56812
rect 1228 56810 1275 56812
rect 2313 56810 2379 56813
rect 5390 56810 5396 56812
rect 1228 56808 1320 56810
rect 1270 56752 1320 56808
rect 1228 56750 1320 56752
rect 2313 56808 5396 56810
rect 2313 56752 2318 56808
rect 2374 56752 5396 56808
rect 2313 56750 5396 56752
rect 1228 56748 1275 56750
rect 1209 56747 1275 56748
rect 2313 56747 2379 56750
rect 5390 56748 5396 56750
rect 5460 56748 5466 56812
rect 0 56674 800 56704
rect 1577 56674 1643 56677
rect 0 56672 1643 56674
rect 0 56616 1582 56672
rect 1638 56616 1643 56672
rect 0 56614 1643 56616
rect 0 56584 800 56614
rect 1577 56611 1643 56614
rect 2262 56612 2268 56676
rect 2332 56674 2338 56676
rect 2497 56674 2563 56677
rect 2332 56672 2563 56674
rect 2332 56616 2502 56672
rect 2558 56616 2563 56672
rect 2332 56614 2563 56616
rect 2332 56612 2338 56614
rect 2497 56611 2563 56614
rect 4208 56608 4528 56609
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 56543 4528 56544
rect 7472 56608 7792 56609
rect 7472 56544 7480 56608
rect 7544 56544 7560 56608
rect 7624 56544 7640 56608
rect 7704 56544 7720 56608
rect 7784 56544 7792 56608
rect 7472 56543 7792 56544
rect 2078 56476 2084 56540
rect 2148 56538 2154 56540
rect 2589 56538 2655 56541
rect 2773 56538 2839 56541
rect 2148 56536 2839 56538
rect 2148 56480 2594 56536
rect 2650 56480 2778 56536
rect 2834 56480 2839 56536
rect 2148 56478 2839 56480
rect 2148 56476 2154 56478
rect 2589 56475 2655 56478
rect 2773 56475 2839 56478
rect 2957 56404 3023 56405
rect 2957 56400 3004 56404
rect 3068 56402 3074 56404
rect 9305 56402 9371 56405
rect 11200 56402 12000 56432
rect 2957 56344 2962 56400
rect 2957 56340 3004 56344
rect 3068 56342 3114 56402
rect 9305 56400 12000 56402
rect 9305 56344 9310 56400
rect 9366 56344 12000 56400
rect 9305 56342 12000 56344
rect 3068 56340 3074 56342
rect 2957 56339 3023 56340
rect 9305 56339 9371 56342
rect 11200 56312 12000 56342
rect 0 56266 800 56296
rect 0 56176 858 56266
rect 798 56130 858 56176
rect 798 56099 904 56130
rect 798 56094 907 56099
rect 798 56070 846 56094
rect 841 56038 846 56070
rect 902 56038 907 56094
rect 841 56033 907 56038
rect 2576 56064 2896 56065
rect 2576 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2576 55999 2896 56000
rect 5840 56064 6160 56065
rect 5840 56000 5848 56064
rect 5912 56000 5928 56064
rect 5992 56000 6008 56064
rect 6072 56000 6088 56064
rect 6152 56000 6160 56064
rect 5840 55999 6160 56000
rect 9104 56064 9424 56065
rect 9104 56000 9112 56064
rect 9176 56000 9192 56064
rect 9256 56000 9272 56064
rect 9336 56000 9352 56064
rect 9416 56000 9424 56064
rect 9104 55999 9424 56000
rect 0 55858 800 55888
rect 3049 55858 3115 55861
rect 0 55856 3115 55858
rect 0 55800 3054 55856
rect 3110 55800 3115 55856
rect 0 55798 3115 55800
rect 0 55768 800 55798
rect 3049 55795 3115 55798
rect 3918 55796 3924 55860
rect 3988 55858 3994 55860
rect 4153 55858 4219 55861
rect 3988 55856 4219 55858
rect 3988 55800 4158 55856
rect 4214 55800 4219 55856
rect 3988 55798 4219 55800
rect 3988 55796 3994 55798
rect 4153 55795 4219 55798
rect 4613 55858 4679 55861
rect 4797 55858 4863 55861
rect 4613 55856 4863 55858
rect 4613 55800 4618 55856
rect 4674 55800 4802 55856
rect 4858 55800 4863 55856
rect 4613 55798 4863 55800
rect 4613 55795 4679 55798
rect 4797 55795 4863 55798
rect 2497 55722 2563 55725
rect 5717 55722 5783 55725
rect 2497 55720 5783 55722
rect 2497 55664 2502 55720
rect 2558 55664 5722 55720
rect 5778 55664 5783 55720
rect 2497 55662 5783 55664
rect 2497 55659 2563 55662
rect 5717 55659 5783 55662
rect 9305 55722 9371 55725
rect 11200 55722 12000 55752
rect 9305 55720 12000 55722
rect 9305 55664 9310 55720
rect 9366 55664 12000 55720
rect 9305 55662 12000 55664
rect 9305 55659 9371 55662
rect 11200 55632 12000 55662
rect 1894 55524 1900 55588
rect 1964 55586 1970 55588
rect 3049 55586 3115 55589
rect 1964 55584 3115 55586
rect 1964 55528 3054 55584
rect 3110 55528 3115 55584
rect 1964 55526 3115 55528
rect 1964 55524 1970 55526
rect 3049 55523 3115 55526
rect 4208 55520 4528 55521
rect 0 55450 800 55480
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 55455 4528 55456
rect 7472 55520 7792 55521
rect 7472 55456 7480 55520
rect 7544 55456 7560 55520
rect 7624 55456 7640 55520
rect 7704 55456 7720 55520
rect 7784 55456 7792 55520
rect 7472 55455 7792 55456
rect 3969 55450 4035 55453
rect 0 55448 4035 55450
rect 0 55392 3974 55448
rect 4030 55392 4035 55448
rect 0 55390 4035 55392
rect 0 55360 800 55390
rect 3969 55387 4035 55390
rect 2313 55316 2379 55317
rect 2262 55314 2268 55316
rect 2222 55254 2268 55314
rect 2332 55312 2379 55316
rect 2374 55256 2379 55312
rect 2262 55252 2268 55254
rect 2332 55252 2379 55256
rect 2313 55251 2379 55252
rect 4153 55314 4219 55317
rect 6310 55314 6316 55316
rect 4153 55312 6316 55314
rect 4153 55256 4158 55312
rect 4214 55256 6316 55312
rect 4153 55254 6316 55256
rect 4153 55251 4219 55254
rect 6310 55252 6316 55254
rect 6380 55252 6386 55316
rect 3417 55178 3483 55181
rect 1350 55176 3483 55178
rect 1350 55120 3422 55176
rect 3478 55120 3483 55176
rect 1350 55118 3483 55120
rect 0 55042 800 55072
rect 1350 55042 1410 55118
rect 3417 55115 3483 55118
rect 0 54982 1410 55042
rect 0 54952 800 54982
rect 2576 54976 2896 54977
rect 2576 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2576 54911 2896 54912
rect 5840 54976 6160 54977
rect 5840 54912 5848 54976
rect 5912 54912 5928 54976
rect 5992 54912 6008 54976
rect 6072 54912 6088 54976
rect 6152 54912 6160 54976
rect 5840 54911 6160 54912
rect 9104 54976 9424 54977
rect 9104 54912 9112 54976
rect 9176 54912 9192 54976
rect 9256 54912 9272 54976
rect 9336 54912 9352 54976
rect 9416 54912 9424 54976
rect 9104 54911 9424 54912
rect 1342 54844 1348 54908
rect 1412 54906 1418 54908
rect 1485 54906 1551 54909
rect 1412 54904 1551 54906
rect 1412 54848 1490 54904
rect 1546 54848 1551 54904
rect 1412 54846 1551 54848
rect 1412 54844 1418 54846
rect 1485 54843 1551 54846
rect 1894 54844 1900 54908
rect 1964 54906 1970 54908
rect 2078 54906 2084 54908
rect 1964 54846 2084 54906
rect 1964 54844 1970 54846
rect 2078 54844 2084 54846
rect 2148 54906 2154 54908
rect 2313 54906 2379 54909
rect 2148 54904 2379 54906
rect 2148 54848 2318 54904
rect 2374 54848 2379 54904
rect 2148 54846 2379 54848
rect 2148 54844 2154 54846
rect 2313 54843 2379 54846
rect 9489 54906 9555 54909
rect 11200 54906 12000 54936
rect 9489 54904 12000 54906
rect 9489 54848 9494 54904
rect 9550 54848 12000 54904
rect 9489 54846 12000 54848
rect 9489 54843 9555 54846
rect 11200 54816 12000 54846
rect 0 54634 800 54664
rect 2497 54634 2563 54637
rect 0 54632 2563 54634
rect 0 54576 2502 54632
rect 2558 54576 2563 54632
rect 0 54574 2563 54576
rect 0 54544 800 54574
rect 2497 54571 2563 54574
rect 2262 54436 2268 54500
rect 2332 54498 2338 54500
rect 3182 54498 3188 54500
rect 2332 54438 3188 54498
rect 2332 54436 2338 54438
rect 3182 54436 3188 54438
rect 3252 54436 3258 54500
rect 4208 54432 4528 54433
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 54367 4528 54368
rect 7472 54432 7792 54433
rect 7472 54368 7480 54432
rect 7544 54368 7560 54432
rect 7624 54368 7640 54432
rect 7704 54368 7720 54432
rect 7784 54368 7792 54432
rect 7472 54367 7792 54368
rect 2957 54362 3023 54365
rect 3918 54362 3924 54364
rect 2957 54360 3924 54362
rect 2957 54304 2962 54360
rect 3018 54304 3924 54360
rect 2957 54302 3924 54304
rect 2957 54299 3023 54302
rect 3918 54300 3924 54302
rect 3988 54300 3994 54364
rect 0 54226 800 54256
rect 2773 54226 2839 54229
rect 0 54224 2839 54226
rect 0 54168 2778 54224
rect 2834 54168 2839 54224
rect 0 54166 2839 54168
rect 0 54136 800 54166
rect 2773 54163 2839 54166
rect 2681 54090 2747 54093
rect 3182 54090 3188 54092
rect 2681 54088 3188 54090
rect 2681 54032 2686 54088
rect 2742 54032 3188 54088
rect 2681 54030 3188 54032
rect 2681 54027 2747 54030
rect 3182 54028 3188 54030
rect 3252 54028 3258 54092
rect 10041 54090 10107 54093
rect 11200 54090 12000 54120
rect 10041 54088 12000 54090
rect 10041 54032 10046 54088
rect 10102 54032 12000 54088
rect 10041 54030 12000 54032
rect 10041 54027 10107 54030
rect 11200 54000 12000 54030
rect 2576 53888 2896 53889
rect 0 53818 800 53848
rect 2576 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2576 53823 2896 53824
rect 5840 53888 6160 53889
rect 5840 53824 5848 53888
rect 5912 53824 5928 53888
rect 5992 53824 6008 53888
rect 6072 53824 6088 53888
rect 6152 53824 6160 53888
rect 5840 53823 6160 53824
rect 9104 53888 9424 53889
rect 9104 53824 9112 53888
rect 9176 53824 9192 53888
rect 9256 53824 9272 53888
rect 9336 53824 9352 53888
rect 9416 53824 9424 53888
rect 9104 53823 9424 53824
rect 2313 53818 2379 53821
rect 0 53816 2379 53818
rect 0 53760 2318 53816
rect 2374 53760 2379 53816
rect 0 53758 2379 53760
rect 0 53728 800 53758
rect 2313 53755 2379 53758
rect 3233 53682 3299 53685
rect 844 53680 3299 53682
rect 844 53624 3238 53680
rect 3294 53624 3299 53680
rect 844 53622 3299 53624
rect 238 53484 244 53548
rect 308 53546 314 53548
rect 844 53546 904 53622
rect 3233 53619 3299 53622
rect 4429 53682 4495 53685
rect 5206 53682 5212 53684
rect 4429 53680 5212 53682
rect 4429 53624 4434 53680
rect 4490 53624 5212 53680
rect 4429 53622 5212 53624
rect 4429 53619 4495 53622
rect 5206 53620 5212 53622
rect 5276 53620 5282 53684
rect 308 53486 904 53546
rect 4521 53546 4587 53549
rect 4654 53546 4660 53548
rect 4521 53544 4660 53546
rect 4521 53488 4526 53544
rect 4582 53488 4660 53544
rect 4521 53486 4660 53488
rect 308 53484 314 53486
rect 4521 53483 4587 53486
rect 4654 53484 4660 53486
rect 4724 53484 4730 53548
rect 10041 53410 10107 53413
rect 11200 53410 12000 53440
rect 10041 53408 12000 53410
rect 10041 53352 10046 53408
rect 10102 53352 12000 53408
rect 10041 53350 12000 53352
rect 10041 53347 10107 53350
rect 4208 53344 4528 53345
rect 0 53274 800 53304
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 53279 4528 53280
rect 7472 53344 7792 53345
rect 7472 53280 7480 53344
rect 7544 53280 7560 53344
rect 7624 53280 7640 53344
rect 7704 53280 7720 53344
rect 7784 53280 7792 53344
rect 11200 53320 12000 53350
rect 7472 53279 7792 53280
rect 1393 53274 1459 53277
rect 0 53272 1459 53274
rect 0 53216 1398 53272
rect 1454 53216 1459 53272
rect 0 53214 1459 53216
rect 0 53184 800 53214
rect 1393 53211 1459 53214
rect 2078 53076 2084 53140
rect 2148 53138 2154 53140
rect 2313 53138 2379 53141
rect 5073 53140 5139 53141
rect 5022 53138 5028 53140
rect 2148 53136 2379 53138
rect 2148 53080 2318 53136
rect 2374 53080 2379 53136
rect 2148 53078 2379 53080
rect 4982 53078 5028 53138
rect 5092 53136 5139 53140
rect 5134 53080 5139 53136
rect 2148 53076 2154 53078
rect 2313 53075 2379 53078
rect 5022 53076 5028 53078
rect 5092 53076 5139 53080
rect 5073 53075 5139 53076
rect 0 52866 800 52896
rect 1577 52866 1643 52869
rect 0 52864 1643 52866
rect 0 52808 1582 52864
rect 1638 52808 1643 52864
rect 0 52806 1643 52808
rect 0 52776 800 52806
rect 1577 52803 1643 52806
rect 2576 52800 2896 52801
rect 2576 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2576 52735 2896 52736
rect 5840 52800 6160 52801
rect 5840 52736 5848 52800
rect 5912 52736 5928 52800
rect 5992 52736 6008 52800
rect 6072 52736 6088 52800
rect 6152 52736 6160 52800
rect 5840 52735 6160 52736
rect 9104 52800 9424 52801
rect 9104 52736 9112 52800
rect 9176 52736 9192 52800
rect 9256 52736 9272 52800
rect 9336 52736 9352 52800
rect 9416 52736 9424 52800
rect 9104 52735 9424 52736
rect 974 52532 980 52596
rect 1044 52594 1050 52596
rect 1485 52594 1551 52597
rect 1044 52592 1551 52594
rect 1044 52536 1490 52592
rect 1546 52536 1551 52592
rect 1044 52534 1551 52536
rect 1044 52532 1050 52534
rect 1485 52531 1551 52534
rect 10041 52594 10107 52597
rect 11200 52594 12000 52624
rect 10041 52592 12000 52594
rect 10041 52536 10046 52592
rect 10102 52536 12000 52592
rect 10041 52534 12000 52536
rect 10041 52531 10107 52534
rect 11200 52504 12000 52534
rect 0 52458 800 52488
rect 2313 52458 2379 52461
rect 0 52456 2379 52458
rect 0 52400 2318 52456
rect 2374 52400 2379 52456
rect 0 52398 2379 52400
rect 0 52368 800 52398
rect 2313 52395 2379 52398
rect 4208 52256 4528 52257
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 52191 4528 52192
rect 7472 52256 7792 52257
rect 7472 52192 7480 52256
rect 7544 52192 7560 52256
rect 7624 52192 7640 52256
rect 7704 52192 7720 52256
rect 7784 52192 7792 52256
rect 7472 52191 7792 52192
rect 2262 52124 2268 52188
rect 2332 52186 2338 52188
rect 2405 52186 2471 52189
rect 2332 52184 2471 52186
rect 2332 52128 2410 52184
rect 2466 52128 2471 52184
rect 2332 52126 2471 52128
rect 2332 52124 2338 52126
rect 2405 52123 2471 52126
rect 0 52050 800 52080
rect 1393 52050 1459 52053
rect 0 52048 1459 52050
rect 0 51992 1398 52048
rect 1454 51992 1459 52048
rect 0 51990 1459 51992
rect 0 51960 800 51990
rect 1393 51987 1459 51990
rect 2078 51988 2084 52052
rect 2148 52050 2154 52052
rect 2313 52050 2379 52053
rect 2148 52048 2379 52050
rect 2148 51992 2318 52048
rect 2374 51992 2379 52048
rect 2148 51990 2379 51992
rect 2148 51988 2154 51990
rect 2313 51987 2379 51990
rect 2078 51852 2084 51916
rect 2148 51914 2154 51916
rect 2497 51914 2563 51917
rect 2148 51912 2563 51914
rect 2148 51856 2502 51912
rect 2558 51856 2563 51912
rect 2148 51854 2563 51856
rect 2148 51852 2154 51854
rect 2497 51851 2563 51854
rect 10041 51778 10107 51781
rect 11200 51778 12000 51808
rect 10041 51776 12000 51778
rect 10041 51720 10046 51776
rect 10102 51720 12000 51776
rect 10041 51718 12000 51720
rect 10041 51715 10107 51718
rect 2576 51712 2896 51713
rect 0 51642 800 51672
rect 2576 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2576 51647 2896 51648
rect 5840 51712 6160 51713
rect 5840 51648 5848 51712
rect 5912 51648 5928 51712
rect 5992 51648 6008 51712
rect 6072 51648 6088 51712
rect 6152 51648 6160 51712
rect 5840 51647 6160 51648
rect 9104 51712 9424 51713
rect 9104 51648 9112 51712
rect 9176 51648 9192 51712
rect 9256 51648 9272 51712
rect 9336 51648 9352 51712
rect 9416 51648 9424 51712
rect 11200 51688 12000 51718
rect 9104 51647 9424 51648
rect 1577 51642 1643 51645
rect 0 51640 1643 51642
rect 0 51584 1582 51640
rect 1638 51584 1643 51640
rect 0 51582 1643 51584
rect 0 51552 800 51582
rect 1577 51579 1643 51582
rect 3049 51508 3115 51509
rect 1158 51444 1164 51508
rect 1228 51506 1234 51508
rect 1228 51446 2376 51506
rect 1228 51444 1234 51446
rect 2316 51373 2376 51446
rect 2998 51444 3004 51508
rect 3068 51506 3115 51508
rect 3068 51504 3160 51506
rect 3110 51448 3160 51504
rect 3068 51446 3160 51448
rect 3068 51444 3115 51446
rect 3049 51443 3115 51444
rect 1761 51370 1827 51373
rect 1894 51370 1900 51372
rect 1761 51368 1900 51370
rect 1761 51312 1766 51368
rect 1822 51312 1900 51368
rect 1761 51310 1900 51312
rect 1761 51307 1827 51310
rect 1894 51308 1900 51310
rect 1964 51308 1970 51372
rect 2313 51368 2379 51373
rect 3141 51370 3207 51373
rect 2313 51312 2318 51368
rect 2374 51312 2379 51368
rect 2313 51307 2379 51312
rect 2822 51368 3207 51370
rect 2822 51312 3146 51368
rect 3202 51312 3207 51368
rect 2822 51310 3207 51312
rect 0 51234 800 51264
rect 1485 51234 1551 51237
rect 1945 51236 2011 51237
rect 1894 51234 1900 51236
rect 0 51232 1551 51234
rect 0 51176 1490 51232
rect 1546 51176 1551 51232
rect 0 51174 1551 51176
rect 1854 51174 1900 51234
rect 1964 51232 2011 51236
rect 2006 51176 2011 51232
rect 0 51144 800 51174
rect 1485 51171 1551 51174
rect 1894 51172 1900 51174
rect 1964 51172 2011 51176
rect 1945 51171 2011 51172
rect 606 50934 612 50998
rect 676 50996 682 50998
rect 676 50962 904 50996
rect 1301 50962 1367 50965
rect 676 50960 1367 50962
rect 676 50936 1306 50960
rect 676 50934 682 50936
rect 844 50904 1306 50936
rect 1362 50904 1367 50960
rect 844 50902 1367 50904
rect 1301 50899 1367 50902
rect 1577 50962 1643 50965
rect 2262 50962 2268 50964
rect 1577 50960 2268 50962
rect 1577 50904 1582 50960
rect 1638 50904 2268 50960
rect 1577 50902 2268 50904
rect 1577 50899 1643 50902
rect 2262 50900 2268 50902
rect 2332 50900 2338 50964
rect 0 50826 800 50856
rect 1945 50826 2011 50829
rect 0 50824 2011 50826
rect 0 50768 1950 50824
rect 2006 50768 2011 50824
rect 0 50766 2011 50768
rect 2822 50826 2882 51310
rect 3141 51307 3207 51310
rect 4838 51172 4844 51236
rect 4908 51234 4914 51236
rect 5073 51234 5139 51237
rect 4908 51232 5139 51234
rect 4908 51176 5078 51232
rect 5134 51176 5139 51232
rect 4908 51174 5139 51176
rect 4908 51172 4914 51174
rect 5073 51171 5139 51174
rect 4208 51168 4528 51169
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 51103 4528 51104
rect 7472 51168 7792 51169
rect 7472 51104 7480 51168
rect 7544 51104 7560 51168
rect 7624 51104 7640 51168
rect 7704 51104 7720 51168
rect 7784 51104 7792 51168
rect 7472 51103 7792 51104
rect 5073 51100 5139 51101
rect 5022 51036 5028 51100
rect 5092 51098 5139 51100
rect 5441 51098 5507 51101
rect 5625 51098 5691 51101
rect 5092 51096 5184 51098
rect 5134 51040 5184 51096
rect 5092 51038 5184 51040
rect 5441 51096 5691 51098
rect 5441 51040 5446 51096
rect 5502 51040 5630 51096
rect 5686 51040 5691 51096
rect 5441 51038 5691 51040
rect 5092 51036 5139 51038
rect 5073 51035 5139 51036
rect 5441 51035 5507 51038
rect 5625 51035 5691 51038
rect 10041 51098 10107 51101
rect 11200 51098 12000 51128
rect 10041 51096 12000 51098
rect 10041 51040 10046 51096
rect 10102 51040 12000 51096
rect 10041 51038 12000 51040
rect 10041 51035 10107 51038
rect 11200 51008 12000 51038
rect 4838 50900 4844 50964
rect 4908 50962 4914 50964
rect 5165 50962 5231 50965
rect 4908 50960 5231 50962
rect 4908 50904 5170 50960
rect 5226 50904 5231 50960
rect 4908 50902 5231 50904
rect 4908 50900 4914 50902
rect 5165 50899 5231 50902
rect 5533 50962 5599 50965
rect 5533 50960 5642 50962
rect 5533 50904 5538 50960
rect 5594 50904 5642 50960
rect 5533 50899 5642 50904
rect 3233 50826 3299 50829
rect 2822 50824 3299 50826
rect 2822 50768 3238 50824
rect 3294 50768 3299 50824
rect 2822 50766 3299 50768
rect 0 50736 800 50766
rect 1945 50763 2011 50766
rect 3233 50763 3299 50766
rect 4654 50764 4660 50828
rect 4724 50826 4730 50828
rect 5349 50826 5415 50829
rect 4724 50824 5415 50826
rect 4724 50768 5354 50824
rect 5410 50768 5415 50824
rect 4724 50766 5415 50768
rect 4724 50764 4730 50766
rect 5349 50763 5415 50766
rect 5257 50690 5323 50693
rect 5582 50690 5642 50899
rect 5257 50688 5642 50690
rect 5257 50632 5262 50688
rect 5318 50632 5642 50688
rect 5257 50630 5642 50632
rect 5257 50627 5323 50630
rect 2576 50624 2896 50625
rect 2576 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2576 50559 2896 50560
rect 5840 50624 6160 50625
rect 5840 50560 5848 50624
rect 5912 50560 5928 50624
rect 5992 50560 6008 50624
rect 6072 50560 6088 50624
rect 6152 50560 6160 50624
rect 5840 50559 6160 50560
rect 9104 50624 9424 50625
rect 9104 50560 9112 50624
rect 9176 50560 9192 50624
rect 9256 50560 9272 50624
rect 9336 50560 9352 50624
rect 9416 50560 9424 50624
rect 9104 50559 9424 50560
rect 1485 50554 1551 50557
rect 798 50552 1551 50554
rect 798 50496 1490 50552
rect 1546 50496 1551 50552
rect 798 50494 1551 50496
rect 798 50448 858 50494
rect 1485 50491 1551 50494
rect 1669 50554 1735 50557
rect 1945 50554 2011 50557
rect 1669 50552 2011 50554
rect 1669 50496 1674 50552
rect 1730 50496 1950 50552
rect 2006 50496 2011 50552
rect 1669 50494 2011 50496
rect 1669 50491 1735 50494
rect 1945 50491 2011 50494
rect 0 50358 858 50448
rect 0 50328 800 50358
rect 1526 50356 1532 50420
rect 1596 50418 1602 50420
rect 1669 50418 1735 50421
rect 1596 50416 1735 50418
rect 1596 50360 1674 50416
rect 1730 50360 1735 50416
rect 1596 50358 1735 50360
rect 1596 50356 1602 50358
rect 1669 50355 1735 50358
rect 3734 50356 3740 50420
rect 3804 50418 3810 50420
rect 4245 50418 4311 50421
rect 3804 50416 4311 50418
rect 3804 50360 4250 50416
rect 4306 50360 4311 50416
rect 3804 50358 4311 50360
rect 3804 50356 3810 50358
rect 4245 50355 4311 50358
rect 4981 50282 5047 50285
rect 5206 50282 5212 50284
rect 4981 50280 5212 50282
rect 4981 50224 4986 50280
rect 5042 50224 5212 50280
rect 4981 50222 5212 50224
rect 4981 50219 5047 50222
rect 5206 50220 5212 50222
rect 5276 50220 5282 50284
rect 10041 50282 10107 50285
rect 11200 50282 12000 50312
rect 10041 50280 12000 50282
rect 10041 50224 10046 50280
rect 10102 50224 12000 50280
rect 10041 50222 12000 50224
rect 10041 50219 10107 50222
rect 11200 50192 12000 50222
rect 422 50084 428 50148
rect 492 50146 498 50148
rect 1526 50146 1532 50148
rect 492 50086 1532 50146
rect 492 50084 498 50086
rect 1526 50084 1532 50086
rect 1596 50084 1602 50148
rect 4208 50080 4528 50081
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 50015 4528 50016
rect 7472 50080 7792 50081
rect 7472 50016 7480 50080
rect 7544 50016 7560 50080
rect 7624 50016 7640 50080
rect 7704 50016 7720 50080
rect 7784 50016 7792 50080
rect 7472 50015 7792 50016
rect 2313 50012 2379 50013
rect 2262 49948 2268 50012
rect 2332 50010 2379 50012
rect 2332 50008 2424 50010
rect 2374 49952 2424 50008
rect 2332 49950 2424 49952
rect 2332 49948 2379 49950
rect 2313 49947 2379 49948
rect 0 49874 800 49904
rect 2773 49874 2839 49877
rect 0 49872 2839 49874
rect 0 49816 2778 49872
rect 2834 49816 2839 49872
rect 0 49814 2839 49816
rect 0 49784 800 49814
rect 2773 49811 2839 49814
rect 1158 49676 1164 49740
rect 1228 49738 1234 49740
rect 1945 49738 2011 49741
rect 1228 49736 2011 49738
rect 1228 49680 1950 49736
rect 2006 49680 2011 49736
rect 1228 49678 2011 49680
rect 1228 49676 1234 49678
rect 1945 49675 2011 49678
rect 1669 49604 1735 49605
rect 1669 49600 1716 49604
rect 1780 49602 1786 49604
rect 1669 49544 1674 49600
rect 1669 49540 1716 49544
rect 1780 49542 1826 49602
rect 1780 49540 1786 49542
rect 1669 49539 1735 49540
rect 2576 49536 2896 49537
rect 0 49466 800 49496
rect 2576 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2576 49471 2896 49472
rect 5840 49536 6160 49537
rect 5840 49472 5848 49536
rect 5912 49472 5928 49536
rect 5992 49472 6008 49536
rect 6072 49472 6088 49536
rect 6152 49472 6160 49536
rect 5840 49471 6160 49472
rect 9104 49536 9424 49537
rect 9104 49472 9112 49536
rect 9176 49472 9192 49536
rect 9256 49472 9272 49536
rect 9336 49472 9352 49536
rect 9416 49472 9424 49536
rect 9104 49471 9424 49472
rect 1393 49466 1459 49469
rect 0 49464 1459 49466
rect 0 49408 1398 49464
rect 1454 49408 1459 49464
rect 0 49406 1459 49408
rect 0 49376 800 49406
rect 1393 49403 1459 49406
rect 3877 49466 3943 49469
rect 4654 49466 4660 49468
rect 3877 49464 4660 49466
rect 3877 49408 3882 49464
rect 3938 49408 4660 49464
rect 3877 49406 4660 49408
rect 3877 49403 3943 49406
rect 4654 49404 4660 49406
rect 4724 49404 4730 49468
rect 9581 49466 9647 49469
rect 11200 49466 12000 49496
rect 9581 49464 12000 49466
rect 9581 49408 9586 49464
rect 9642 49408 12000 49464
rect 9581 49406 12000 49408
rect 9581 49403 9647 49406
rect 11200 49376 12000 49406
rect 3325 49330 3391 49333
rect 3918 49330 3924 49332
rect 3325 49328 3924 49330
rect 3325 49272 3330 49328
rect 3386 49272 3924 49328
rect 3325 49270 3924 49272
rect 3325 49267 3391 49270
rect 3918 49268 3924 49270
rect 3988 49268 3994 49332
rect 3969 49196 4035 49197
rect 1710 49132 1716 49196
rect 1780 49194 1786 49196
rect 3550 49194 3556 49196
rect 1780 49134 3556 49194
rect 1780 49132 1786 49134
rect 3550 49132 3556 49134
rect 3620 49132 3626 49196
rect 3918 49194 3924 49196
rect 3878 49134 3924 49194
rect 3988 49192 4035 49196
rect 4030 49136 4035 49192
rect 3918 49132 3924 49134
rect 3988 49132 4035 49136
rect 3969 49131 4035 49132
rect 4521 49194 4587 49197
rect 5206 49194 5212 49196
rect 4521 49192 5212 49194
rect 4521 49136 4526 49192
rect 4582 49136 5212 49192
rect 4521 49134 5212 49136
rect 4521 49131 4587 49134
rect 5206 49132 5212 49134
rect 5276 49132 5282 49196
rect 0 49058 800 49088
rect 3969 49058 4035 49061
rect 0 49056 4035 49058
rect 0 49000 3974 49056
rect 4030 49000 4035 49056
rect 0 48998 4035 49000
rect 0 48968 800 48998
rect 3969 48995 4035 48998
rect 4208 48992 4528 48993
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 48927 4528 48928
rect 7472 48992 7792 48993
rect 7472 48928 7480 48992
rect 7544 48928 7560 48992
rect 7624 48928 7640 48992
rect 7704 48928 7720 48992
rect 7784 48928 7792 48992
rect 7472 48927 7792 48928
rect 1669 48922 1735 48925
rect 2681 48922 2747 48925
rect 1669 48920 2747 48922
rect 1669 48864 1674 48920
rect 1730 48864 2686 48920
rect 2742 48864 2747 48920
rect 1669 48862 2747 48864
rect 1669 48859 1735 48862
rect 2681 48859 2747 48862
rect 3049 48922 3115 48925
rect 3969 48922 4035 48925
rect 3049 48920 4035 48922
rect 3049 48864 3054 48920
rect 3110 48864 3974 48920
rect 4030 48864 4035 48920
rect 3049 48862 4035 48864
rect 3049 48859 3115 48862
rect 3969 48859 4035 48862
rect 10041 48786 10107 48789
rect 11200 48786 12000 48816
rect 10041 48784 12000 48786
rect 10041 48728 10046 48784
rect 10102 48728 12000 48784
rect 10041 48726 12000 48728
rect 10041 48723 10107 48726
rect 11200 48696 12000 48726
rect 0 48650 800 48680
rect 2221 48650 2287 48653
rect 0 48648 2287 48650
rect 0 48592 2226 48648
rect 2282 48592 2287 48648
rect 0 48590 2287 48592
rect 0 48560 800 48590
rect 2221 48587 2287 48590
rect 2773 48650 2839 48653
rect 2773 48648 3020 48650
rect 2773 48592 2778 48648
rect 2834 48592 3020 48648
rect 2773 48590 3020 48592
rect 2773 48587 2839 48590
rect 1526 48452 1532 48516
rect 1596 48452 1602 48516
rect 1761 48514 1827 48517
rect 1894 48514 1900 48516
rect 1761 48512 1900 48514
rect 1761 48456 1766 48512
rect 1822 48456 1900 48512
rect 1761 48454 1900 48456
rect 1534 48378 1594 48452
rect 1761 48451 1827 48454
rect 1894 48452 1900 48454
rect 1964 48452 1970 48516
rect 2576 48448 2896 48449
rect 2576 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2576 48383 2896 48384
rect 2960 48381 3020 48590
rect 3550 48588 3556 48652
rect 3620 48650 3626 48652
rect 3969 48650 4035 48653
rect 3620 48648 4035 48650
rect 3620 48592 3974 48648
rect 4030 48592 4035 48648
rect 3620 48590 4035 48592
rect 3620 48588 3626 48590
rect 3969 48587 4035 48590
rect 5840 48448 6160 48449
rect 5840 48384 5848 48448
rect 5912 48384 5928 48448
rect 5992 48384 6008 48448
rect 6072 48384 6088 48448
rect 6152 48384 6160 48448
rect 5840 48383 6160 48384
rect 9104 48448 9424 48449
rect 9104 48384 9112 48448
rect 9176 48384 9192 48448
rect 9256 48384 9272 48448
rect 9336 48384 9352 48448
rect 9416 48384 9424 48448
rect 9104 48383 9424 48384
rect 2313 48378 2379 48381
rect 1534 48376 2379 48378
rect 1534 48320 2318 48376
rect 2374 48320 2379 48376
rect 1534 48318 2379 48320
rect 2313 48315 2379 48318
rect 2957 48376 3023 48381
rect 2957 48320 2962 48376
rect 3018 48320 3023 48376
rect 2957 48315 3023 48320
rect 3877 48378 3943 48381
rect 4654 48378 4660 48380
rect 3877 48376 4660 48378
rect 3877 48320 3882 48376
rect 3938 48320 4660 48376
rect 3877 48318 4660 48320
rect 3877 48315 3943 48318
rect 4654 48316 4660 48318
rect 4724 48316 4730 48380
rect 0 48242 800 48272
rect 3785 48242 3851 48245
rect 0 48240 3851 48242
rect 0 48184 3790 48240
rect 3846 48184 3851 48240
rect 0 48182 3851 48184
rect 0 48152 800 48182
rect 3785 48179 3851 48182
rect 1342 48044 1348 48108
rect 1412 48106 1418 48108
rect 1894 48106 1900 48108
rect 1412 48046 1900 48106
rect 1412 48044 1418 48046
rect 1894 48044 1900 48046
rect 1964 48044 1970 48108
rect 3785 48106 3851 48109
rect 5390 48106 5396 48108
rect 3785 48104 5396 48106
rect 3785 48048 3790 48104
rect 3846 48048 5396 48104
rect 3785 48046 5396 48048
rect 3785 48043 3851 48046
rect 5390 48044 5396 48046
rect 5460 48044 5466 48108
rect 1301 47970 1367 47973
rect 1526 47970 1532 47972
rect 1301 47968 1532 47970
rect 1301 47912 1306 47968
rect 1362 47912 1532 47968
rect 1301 47910 1532 47912
rect 1301 47907 1367 47910
rect 1526 47908 1532 47910
rect 1596 47908 1602 47972
rect 10041 47970 10107 47973
rect 11200 47970 12000 48000
rect 10041 47968 12000 47970
rect 10041 47912 10046 47968
rect 10102 47912 12000 47968
rect 10041 47910 12000 47912
rect 10041 47907 10107 47910
rect 4208 47904 4528 47905
rect 0 47834 800 47864
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 47839 4528 47840
rect 7472 47904 7792 47905
rect 7472 47840 7480 47904
rect 7544 47840 7560 47904
rect 7624 47840 7640 47904
rect 7704 47840 7720 47904
rect 7784 47840 7792 47904
rect 11200 47880 12000 47910
rect 7472 47839 7792 47840
rect 1577 47834 1643 47837
rect 0 47832 1643 47834
rect 0 47776 1582 47832
rect 1638 47776 1643 47832
rect 0 47774 1643 47776
rect 0 47744 800 47774
rect 1577 47771 1643 47774
rect 1393 47562 1459 47565
rect 5390 47562 5396 47564
rect 1393 47560 5396 47562
rect 1393 47504 1398 47560
rect 1454 47504 5396 47560
rect 1393 47502 5396 47504
rect 1393 47499 1459 47502
rect 5390 47500 5396 47502
rect 5460 47500 5466 47564
rect 0 47426 800 47456
rect 1577 47426 1643 47429
rect 0 47424 1643 47426
rect 0 47368 1582 47424
rect 1638 47368 1643 47424
rect 0 47366 1643 47368
rect 0 47336 800 47366
rect 1577 47363 1643 47366
rect 2576 47360 2896 47361
rect 2576 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2576 47295 2896 47296
rect 5840 47360 6160 47361
rect 5840 47296 5848 47360
rect 5912 47296 5928 47360
rect 5992 47296 6008 47360
rect 6072 47296 6088 47360
rect 6152 47296 6160 47360
rect 5840 47295 6160 47296
rect 9104 47360 9424 47361
rect 9104 47296 9112 47360
rect 9176 47296 9192 47360
rect 9256 47296 9272 47360
rect 9336 47296 9352 47360
rect 9416 47296 9424 47360
rect 9104 47295 9424 47296
rect 1761 47154 1827 47157
rect 3182 47154 3188 47156
rect 1761 47152 3188 47154
rect 1761 47096 1766 47152
rect 1822 47096 3188 47152
rect 1761 47094 3188 47096
rect 1761 47091 1827 47094
rect 3182 47092 3188 47094
rect 3252 47092 3258 47156
rect 10041 47154 10107 47157
rect 11200 47154 12000 47184
rect 10041 47152 12000 47154
rect 10041 47096 10046 47152
rect 10102 47096 12000 47152
rect 10041 47094 12000 47096
rect 10041 47091 10107 47094
rect 11200 47064 12000 47094
rect 0 47018 800 47048
rect 3969 47018 4035 47021
rect 0 47016 4035 47018
rect 0 46960 3974 47016
rect 4030 46960 4035 47016
rect 0 46958 4035 46960
rect 0 46928 800 46958
rect 3969 46955 4035 46958
rect 4245 47018 4311 47021
rect 4654 47018 4660 47020
rect 4245 47016 4660 47018
rect 4245 46960 4250 47016
rect 4306 46960 4660 47016
rect 4245 46958 4660 46960
rect 4245 46955 4311 46958
rect 4654 46956 4660 46958
rect 4724 46956 4730 47020
rect 1025 46882 1091 46885
rect 2998 46882 3004 46884
rect 1025 46880 3004 46882
rect 1025 46824 1030 46880
rect 1086 46824 3004 46880
rect 1025 46822 3004 46824
rect 1025 46819 1091 46822
rect 2998 46820 3004 46822
rect 3068 46820 3074 46884
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 7472 46816 7792 46817
rect 7472 46752 7480 46816
rect 7544 46752 7560 46816
rect 7624 46752 7640 46816
rect 7704 46752 7720 46816
rect 7784 46752 7792 46816
rect 7472 46751 7792 46752
rect 422 46684 428 46748
rect 492 46746 498 46748
rect 1526 46746 1532 46748
rect 492 46686 1532 46746
rect 492 46684 498 46686
rect 1526 46684 1532 46686
rect 1596 46684 1602 46748
rect 3182 46684 3188 46748
rect 3252 46746 3258 46748
rect 3550 46746 3556 46748
rect 3252 46686 3556 46746
rect 3252 46684 3258 46686
rect 3550 46684 3556 46686
rect 3620 46684 3626 46748
rect 2313 46610 2379 46613
rect 3550 46610 3556 46612
rect 2313 46608 3556 46610
rect 2313 46552 2318 46608
rect 2374 46552 3556 46608
rect 2313 46550 3556 46552
rect 2313 46547 2379 46550
rect 3550 46548 3556 46550
rect 3620 46548 3626 46612
rect 0 46474 800 46504
rect 2313 46474 2379 46477
rect 0 46472 2379 46474
rect 0 46416 2318 46472
rect 2374 46416 2379 46472
rect 0 46414 2379 46416
rect 0 46384 800 46414
rect 2313 46411 2379 46414
rect 2497 46474 2563 46477
rect 3417 46474 3483 46477
rect 5022 46474 5028 46476
rect 2497 46472 3020 46474
rect 2497 46416 2502 46472
rect 2558 46416 3020 46472
rect 2497 46414 3020 46416
rect 2497 46411 2563 46414
rect 2576 46272 2896 46273
rect 2576 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2576 46207 2896 46208
rect 0 46066 800 46096
rect 2497 46066 2563 46069
rect 2960 46066 3020 46414
rect 3417 46472 5028 46474
rect 3417 46416 3422 46472
rect 3478 46416 5028 46472
rect 3417 46414 5028 46416
rect 3417 46411 3483 46414
rect 5022 46412 5028 46414
rect 5092 46412 5098 46476
rect 10041 46474 10107 46477
rect 11200 46474 12000 46504
rect 10041 46472 12000 46474
rect 10041 46416 10046 46472
rect 10102 46416 12000 46472
rect 10041 46414 12000 46416
rect 10041 46411 10107 46414
rect 11200 46384 12000 46414
rect 5840 46272 6160 46273
rect 5840 46208 5848 46272
rect 5912 46208 5928 46272
rect 5992 46208 6008 46272
rect 6072 46208 6088 46272
rect 6152 46208 6160 46272
rect 5840 46207 6160 46208
rect 9104 46272 9424 46273
rect 9104 46208 9112 46272
rect 9176 46208 9192 46272
rect 9256 46208 9272 46272
rect 9336 46208 9352 46272
rect 9416 46208 9424 46272
rect 9104 46207 9424 46208
rect 0 46064 2563 46066
rect 0 46008 2502 46064
rect 2558 46008 2563 46064
rect 0 46006 2563 46008
rect 0 45976 800 46006
rect 2497 46003 2563 46006
rect 2638 46006 3020 46066
rect 2497 45930 2563 45933
rect 2638 45930 2698 46006
rect 2497 45928 2698 45930
rect 2497 45872 2502 45928
rect 2558 45872 2698 45928
rect 2497 45870 2698 45872
rect 2865 45930 2931 45933
rect 2865 45928 4722 45930
rect 2865 45872 2870 45928
rect 2926 45872 4722 45928
rect 2865 45870 4722 45872
rect 2497 45867 2563 45870
rect 2865 45867 2931 45870
rect 13 45828 79 45831
rect 606 45828 612 45830
rect 13 45826 612 45828
rect 13 45770 18 45826
rect 74 45770 612 45826
rect 13 45768 612 45770
rect 13 45765 79 45768
rect 606 45766 612 45768
rect 676 45766 682 45830
rect 3049 45794 3115 45797
rect 1350 45792 3115 45794
rect 1350 45736 3054 45792
rect 3110 45736 3115 45792
rect 1350 45734 3115 45736
rect 4662 45794 4722 45870
rect 4838 45794 4844 45796
rect 4662 45734 4844 45794
rect 0 45658 800 45688
rect 1350 45658 1410 45734
rect 3049 45731 3115 45734
rect 4838 45732 4844 45734
rect 4908 45732 4914 45796
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 7472 45728 7792 45729
rect 7472 45664 7480 45728
rect 7544 45664 7560 45728
rect 7624 45664 7640 45728
rect 7704 45664 7720 45728
rect 7784 45664 7792 45728
rect 7472 45663 7792 45664
rect 0 45598 1410 45658
rect 3785 45658 3851 45661
rect 3969 45658 4035 45661
rect 3785 45656 4035 45658
rect 3785 45600 3790 45656
rect 3846 45600 3974 45656
rect 4030 45600 4035 45656
rect 3785 45598 4035 45600
rect 0 45568 800 45598
rect 3785 45595 3851 45598
rect 3969 45595 4035 45598
rect 5349 45658 5415 45661
rect 10041 45658 10107 45661
rect 11200 45658 12000 45688
rect 5349 45656 5458 45658
rect 5349 45600 5354 45656
rect 5410 45600 5458 45656
rect 5349 45595 5458 45600
rect 10041 45656 12000 45658
rect 10041 45600 10046 45656
rect 10102 45600 12000 45656
rect 10041 45598 12000 45600
rect 10041 45595 10107 45598
rect 1342 45460 1348 45524
rect 1412 45522 1418 45524
rect 1577 45522 1643 45525
rect 1412 45520 1643 45522
rect 1412 45464 1582 45520
rect 1638 45464 1643 45520
rect 1412 45462 1643 45464
rect 1412 45460 1418 45462
rect 1577 45459 1643 45462
rect 1710 45460 1716 45524
rect 1780 45522 1786 45524
rect 2313 45522 2379 45525
rect 1780 45520 2379 45522
rect 1780 45464 2318 45520
rect 2374 45464 2379 45520
rect 1780 45462 2379 45464
rect 1780 45460 1786 45462
rect 2313 45459 2379 45462
rect 2865 45522 2931 45525
rect 2998 45522 3004 45524
rect 2865 45520 3004 45522
rect 2865 45464 2870 45520
rect 2926 45464 3004 45520
rect 2865 45462 3004 45464
rect 2865 45459 2931 45462
rect 2998 45460 3004 45462
rect 3068 45460 3074 45524
rect 2589 45386 2655 45389
rect 1534 45384 2655 45386
rect 1534 45328 2594 45384
rect 2650 45328 2655 45384
rect 1534 45326 2655 45328
rect 0 45250 800 45280
rect 1534 45250 1594 45326
rect 2589 45323 2655 45326
rect 0 45190 1594 45250
rect 0 45160 800 45190
rect 2576 45184 2896 45185
rect 2576 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2576 45119 2896 45120
rect 5398 44981 5458 45595
rect 11200 45568 12000 45598
rect 5840 45184 6160 45185
rect 5840 45120 5848 45184
rect 5912 45120 5928 45184
rect 5992 45120 6008 45184
rect 6072 45120 6088 45184
rect 6152 45120 6160 45184
rect 5840 45119 6160 45120
rect 9104 45184 9424 45185
rect 9104 45120 9112 45184
rect 9176 45120 9192 45184
rect 9256 45120 9272 45184
rect 9336 45120 9352 45184
rect 9416 45120 9424 45184
rect 9104 45119 9424 45120
rect 3734 44978 3740 44980
rect 3558 44918 3740 44978
rect 0 44842 800 44872
rect 1577 44842 1643 44845
rect 0 44840 1643 44842
rect 0 44784 1582 44840
rect 1638 44784 1643 44840
rect 0 44782 1643 44784
rect 0 44752 800 44782
rect 1577 44779 1643 44782
rect 2313 44842 2379 44845
rect 3366 44842 3372 44844
rect 2313 44840 3372 44842
rect 2313 44784 2318 44840
rect 2374 44784 3372 44840
rect 2313 44782 3372 44784
rect 2313 44779 2379 44782
rect 3366 44780 3372 44782
rect 3436 44780 3442 44844
rect 2957 44706 3023 44709
rect 1350 44704 3023 44706
rect 1350 44648 2962 44704
rect 3018 44648 3023 44704
rect 1350 44646 3023 44648
rect 0 44434 800 44464
rect 1350 44434 1410 44646
rect 2957 44643 3023 44646
rect 1526 44508 1532 44572
rect 1596 44570 1602 44572
rect 3558 44570 3618 44918
rect 3734 44916 3740 44918
rect 3804 44916 3810 44980
rect 5349 44976 5458 44981
rect 5349 44920 5354 44976
rect 5410 44920 5458 44976
rect 5349 44918 5458 44920
rect 5349 44915 5415 44918
rect 3734 44780 3740 44844
rect 3804 44842 3810 44844
rect 4153 44842 4219 44845
rect 3804 44840 4219 44842
rect 3804 44784 4158 44840
rect 4214 44784 4219 44840
rect 3804 44782 4219 44784
rect 3804 44780 3810 44782
rect 4153 44779 4219 44782
rect 10041 44842 10107 44845
rect 11200 44842 12000 44872
rect 10041 44840 12000 44842
rect 10041 44784 10046 44840
rect 10102 44784 12000 44840
rect 10041 44782 12000 44784
rect 10041 44779 10107 44782
rect 11200 44752 12000 44782
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 7472 44640 7792 44641
rect 7472 44576 7480 44640
rect 7544 44576 7560 44640
rect 7624 44576 7640 44640
rect 7704 44576 7720 44640
rect 7784 44576 7792 44640
rect 7472 44575 7792 44576
rect 1596 44510 3618 44570
rect 1596 44508 1602 44510
rect 0 44374 1410 44434
rect 0 44344 800 44374
rect 3141 44300 3207 44301
rect 3141 44296 3188 44300
rect 3252 44298 3258 44300
rect 3141 44240 3146 44296
rect 3141 44236 3188 44240
rect 3252 44238 3298 44298
rect 3252 44236 3258 44238
rect 3141 44235 3207 44236
rect 10041 44162 10107 44165
rect 11200 44162 12000 44192
rect 10041 44160 12000 44162
rect 10041 44104 10046 44160
rect 10102 44104 12000 44160
rect 10041 44102 12000 44104
rect 10041 44099 10107 44102
rect 2576 44096 2896 44097
rect 0 44026 800 44056
rect 2576 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2576 44031 2896 44032
rect 5840 44096 6160 44097
rect 5840 44032 5848 44096
rect 5912 44032 5928 44096
rect 5992 44032 6008 44096
rect 6072 44032 6088 44096
rect 6152 44032 6160 44096
rect 5840 44031 6160 44032
rect 9104 44096 9424 44097
rect 9104 44032 9112 44096
rect 9176 44032 9192 44096
rect 9256 44032 9272 44096
rect 9336 44032 9352 44096
rect 9416 44032 9424 44096
rect 11200 44072 12000 44102
rect 9104 44031 9424 44032
rect 0 43966 1410 44026
rect 0 43936 800 43966
rect 1350 43890 1410 43966
rect 3141 43890 3207 43893
rect 1350 43888 3207 43890
rect 1350 43832 3146 43888
rect 3202 43832 3207 43888
rect 1350 43830 3207 43832
rect 3141 43827 3207 43830
rect 0 43618 800 43648
rect 3969 43618 4035 43621
rect 0 43616 4035 43618
rect 0 43560 3974 43616
rect 4030 43560 4035 43616
rect 0 43558 4035 43560
rect 0 43528 800 43558
rect 3969 43555 4035 43558
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 7472 43552 7792 43553
rect 7472 43488 7480 43552
rect 7544 43488 7560 43552
rect 7624 43488 7640 43552
rect 7704 43488 7720 43552
rect 7784 43488 7792 43552
rect 7472 43487 7792 43488
rect 1710 43420 1716 43484
rect 1780 43482 1786 43484
rect 3049 43482 3115 43485
rect 1780 43480 3115 43482
rect 1780 43424 3054 43480
rect 3110 43424 3115 43480
rect 1780 43422 3115 43424
rect 1780 43420 1786 43422
rect 3049 43419 3115 43422
rect 790 43284 796 43348
rect 860 43346 866 43348
rect 4153 43346 4219 43349
rect 860 43344 4219 43346
rect 860 43288 4158 43344
rect 4214 43288 4219 43344
rect 860 43286 4219 43288
rect 860 43284 866 43286
rect 4153 43283 4219 43286
rect 10041 43346 10107 43349
rect 11200 43346 12000 43376
rect 10041 43344 12000 43346
rect 10041 43288 10046 43344
rect 10102 43288 12000 43344
rect 10041 43286 12000 43288
rect 10041 43283 10107 43286
rect 11200 43256 12000 43286
rect 3969 43210 4035 43213
rect 1350 43208 4035 43210
rect 1350 43152 3974 43208
rect 4030 43152 4035 43208
rect 1350 43150 4035 43152
rect 0 43074 800 43104
rect 1350 43074 1410 43150
rect 3969 43147 4035 43150
rect 0 43014 1410 43074
rect 0 42984 800 43014
rect 3366 43012 3372 43076
rect 3436 43074 3442 43076
rect 3601 43074 3667 43077
rect 3436 43072 3667 43074
rect 3436 43016 3606 43072
rect 3662 43016 3667 43072
rect 3436 43014 3667 43016
rect 3436 43012 3442 43014
rect 3601 43011 3667 43014
rect 2576 43008 2896 43009
rect 2576 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2576 42943 2896 42944
rect 5840 43008 6160 43009
rect 5840 42944 5848 43008
rect 5912 42944 5928 43008
rect 5992 42944 6008 43008
rect 6072 42944 6088 43008
rect 6152 42944 6160 43008
rect 5840 42943 6160 42944
rect 9104 43008 9424 43009
rect 9104 42944 9112 43008
rect 9176 42944 9192 43008
rect 9256 42944 9272 43008
rect 9336 42944 9352 43008
rect 9416 42944 9424 43008
rect 9104 42943 9424 42944
rect 2957 42938 3023 42941
rect 2957 42936 3066 42938
rect 2957 42880 2962 42936
rect 3018 42880 3066 42936
rect 2957 42875 3066 42880
rect 2865 42802 2931 42805
rect 3006 42802 3066 42875
rect 2865 42800 3066 42802
rect 2865 42744 2870 42800
rect 2926 42744 3066 42800
rect 2865 42742 3066 42744
rect 2865 42739 2931 42742
rect 3366 42740 3372 42804
rect 3436 42802 3442 42804
rect 4654 42802 4660 42804
rect 3436 42742 4660 42802
rect 3436 42740 3442 42742
rect 4654 42740 4660 42742
rect 4724 42740 4730 42804
rect 0 42666 800 42696
rect 3969 42666 4035 42669
rect 0 42664 4035 42666
rect 0 42608 3974 42664
rect 4030 42608 4035 42664
rect 0 42606 4035 42608
rect 0 42576 800 42606
rect 3969 42603 4035 42606
rect 1669 42530 1735 42533
rect 1894 42530 1900 42532
rect 1669 42528 1900 42530
rect 1669 42472 1674 42528
rect 1730 42472 1900 42528
rect 1669 42470 1900 42472
rect 1669 42467 1735 42470
rect 1894 42468 1900 42470
rect 1964 42468 1970 42532
rect 10041 42530 10107 42533
rect 11200 42530 12000 42560
rect 10041 42528 12000 42530
rect 10041 42472 10046 42528
rect 10102 42472 12000 42528
rect 10041 42470 12000 42472
rect 10041 42467 10107 42470
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 7472 42464 7792 42465
rect 7472 42400 7480 42464
rect 7544 42400 7560 42464
rect 7624 42400 7640 42464
rect 7704 42400 7720 42464
rect 7784 42400 7792 42464
rect 11200 42440 12000 42470
rect 7472 42399 7792 42400
rect 1761 42394 1827 42397
rect 2262 42394 2268 42396
rect 1761 42392 2268 42394
rect 1761 42336 1766 42392
rect 1822 42336 2268 42392
rect 1761 42334 2268 42336
rect 1761 42331 1827 42334
rect 2262 42332 2268 42334
rect 2332 42332 2338 42396
rect 0 42258 800 42288
rect 2773 42258 2839 42261
rect 0 42256 2839 42258
rect 0 42200 2778 42256
rect 2834 42200 2839 42256
rect 0 42198 2839 42200
rect 0 42168 800 42198
rect 2773 42195 2839 42198
rect 3325 42258 3391 42261
rect 3550 42258 3556 42260
rect 3325 42256 3556 42258
rect 3325 42200 3330 42256
rect 3386 42200 3556 42256
rect 3325 42198 3556 42200
rect 3325 42195 3391 42198
rect 3550 42196 3556 42198
rect 3620 42196 3626 42260
rect 1894 42060 1900 42124
rect 1964 42122 1970 42124
rect 2497 42122 2563 42125
rect 1964 42120 2563 42122
rect 1964 42064 2502 42120
rect 2558 42064 2563 42120
rect 1964 42062 2563 42064
rect 1964 42060 1970 42062
rect 2497 42059 2563 42062
rect 4797 42122 4863 42125
rect 5206 42122 5212 42124
rect 4797 42120 5212 42122
rect 4797 42064 4802 42120
rect 4858 42064 5212 42120
rect 4797 42062 5212 42064
rect 4797 42059 4863 42062
rect 5206 42060 5212 42062
rect 5276 42060 5282 42124
rect 5206 41924 5212 41988
rect 5276 41986 5282 41988
rect 5625 41986 5691 41989
rect 5276 41984 5691 41986
rect 5276 41928 5630 41984
rect 5686 41928 5691 41984
rect 5276 41926 5691 41928
rect 5276 41924 5282 41926
rect 5625 41923 5691 41926
rect 2576 41920 2896 41921
rect 0 41850 800 41880
rect 2576 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2576 41855 2896 41856
rect 5840 41920 6160 41921
rect 5840 41856 5848 41920
rect 5912 41856 5928 41920
rect 5992 41856 6008 41920
rect 6072 41856 6088 41920
rect 6152 41856 6160 41920
rect 5840 41855 6160 41856
rect 9104 41920 9424 41921
rect 9104 41856 9112 41920
rect 9176 41856 9192 41920
rect 9256 41856 9272 41920
rect 9336 41856 9352 41920
rect 9416 41856 9424 41920
rect 9104 41855 9424 41856
rect 10041 41850 10107 41853
rect 11200 41850 12000 41880
rect 0 41790 1410 41850
rect 0 41760 800 41790
rect 1350 41714 1410 41790
rect 10041 41848 12000 41850
rect 10041 41792 10046 41848
rect 10102 41792 12000 41848
rect 10041 41790 12000 41792
rect 10041 41787 10107 41790
rect 11200 41760 12000 41790
rect 3049 41714 3115 41717
rect 1350 41712 3115 41714
rect 1350 41656 3054 41712
rect 3110 41656 3115 41712
rect 1350 41654 3115 41656
rect 3049 41651 3115 41654
rect 3601 41712 3667 41717
rect 3601 41656 3606 41712
rect 3662 41656 3667 41712
rect 3601 41651 3667 41656
rect 2405 41578 2471 41581
rect 2998 41578 3004 41580
rect 2405 41576 3004 41578
rect 2405 41520 2410 41576
rect 2466 41520 3004 41576
rect 2405 41518 3004 41520
rect 2405 41515 2471 41518
rect 2998 41516 3004 41518
rect 3068 41516 3074 41580
rect 0 41442 800 41472
rect 2313 41442 2379 41445
rect 0 41440 2379 41442
rect 0 41384 2318 41440
rect 2374 41384 2379 41440
rect 0 41382 2379 41384
rect 0 41352 800 41382
rect 2313 41379 2379 41382
rect 2221 41306 2287 41309
rect 1534 41304 2287 41306
rect 1534 41248 2226 41304
rect 2282 41248 2287 41304
rect 1534 41246 2287 41248
rect 1534 41173 1594 41246
rect 2221 41243 2287 41246
rect 3604 41173 3664 41651
rect 4429 41578 4495 41581
rect 3972 41576 4495 41578
rect 3972 41520 4434 41576
rect 4490 41520 4495 41576
rect 3972 41518 4495 41520
rect 1485 41168 1594 41173
rect 1485 41112 1490 41168
rect 1546 41112 1594 41168
rect 1485 41110 1594 41112
rect 1485 41107 1551 41110
rect 1894 41108 1900 41172
rect 1964 41170 1970 41172
rect 2221 41170 2287 41173
rect 1964 41168 2287 41170
rect 1964 41112 2226 41168
rect 2282 41112 2287 41168
rect 1964 41110 2287 41112
rect 1964 41108 1970 41110
rect 2221 41107 2287 41110
rect 3601 41168 3667 41173
rect 3601 41112 3606 41168
rect 3662 41112 3667 41168
rect 3601 41107 3667 41112
rect 0 41034 800 41064
rect 2773 41034 2839 41037
rect 3049 41036 3115 41037
rect 0 41000 2376 41034
rect 2638 41032 2839 41034
rect 2638 41000 2778 41032
rect 0 40976 2778 41000
rect 2834 40976 2839 41032
rect 0 40974 2839 40976
rect 0 40944 800 40974
rect 2316 40940 2698 40974
rect 2773 40971 2839 40974
rect 2998 40972 3004 41036
rect 3068 41034 3115 41036
rect 3693 41034 3759 41037
rect 3972 41034 4032 41518
rect 4429 41515 4495 41518
rect 4654 41516 4660 41580
rect 4724 41578 4730 41580
rect 5073 41578 5139 41581
rect 4724 41576 5139 41578
rect 4724 41520 5078 41576
rect 5134 41520 5139 41576
rect 4724 41518 5139 41520
rect 4724 41516 4730 41518
rect 5073 41515 5139 41518
rect 5349 41442 5415 41445
rect 6545 41442 6611 41445
rect 5349 41440 6611 41442
rect 5349 41384 5354 41440
rect 5410 41384 6550 41440
rect 6606 41384 6611 41440
rect 5349 41382 6611 41384
rect 5349 41379 5415 41382
rect 6545 41379 6611 41382
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 7472 41376 7792 41377
rect 7472 41312 7480 41376
rect 7544 41312 7560 41376
rect 7624 41312 7640 41376
rect 7704 41312 7720 41376
rect 7784 41312 7792 41376
rect 7472 41311 7792 41312
rect 3068 41032 3160 41034
rect 3110 40976 3160 41032
rect 3068 40974 3160 40976
rect 3693 41032 4032 41034
rect 3693 40976 3698 41032
rect 3754 40976 4032 41032
rect 3693 40974 4032 40976
rect 10041 41034 10107 41037
rect 11200 41034 12000 41064
rect 10041 41032 12000 41034
rect 10041 40976 10046 41032
rect 10102 40976 12000 41032
rect 10041 40974 12000 40976
rect 3068 40972 3115 40974
rect 3049 40971 3115 40972
rect 3693 40971 3759 40974
rect 10041 40971 10107 40974
rect 11200 40944 12000 40974
rect 1526 40836 1532 40900
rect 1596 40898 1602 40900
rect 1669 40898 1735 40901
rect 1596 40896 1735 40898
rect 1596 40840 1674 40896
rect 1730 40840 1735 40896
rect 1596 40838 1735 40840
rect 1596 40836 1602 40838
rect 1669 40835 1735 40838
rect 2576 40832 2896 40833
rect 2576 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2576 40767 2896 40768
rect 5840 40832 6160 40833
rect 5840 40768 5848 40832
rect 5912 40768 5928 40832
rect 5992 40768 6008 40832
rect 6072 40768 6088 40832
rect 6152 40768 6160 40832
rect 5840 40767 6160 40768
rect 9104 40832 9424 40833
rect 9104 40768 9112 40832
rect 9176 40768 9192 40832
rect 9256 40768 9272 40832
rect 9336 40768 9352 40832
rect 9416 40768 9424 40832
rect 9104 40767 9424 40768
rect 1761 40764 1827 40765
rect 1710 40700 1716 40764
rect 1780 40762 1827 40764
rect 1780 40760 1872 40762
rect 1822 40704 1872 40760
rect 1780 40702 1872 40704
rect 1780 40700 1827 40702
rect 1761 40699 1827 40700
rect 0 40626 800 40656
rect 1577 40626 1643 40629
rect 0 40624 1643 40626
rect 0 40568 1582 40624
rect 1638 40568 1643 40624
rect 0 40566 1643 40568
rect 0 40536 800 40566
rect 1577 40563 1643 40566
rect 10041 40354 10107 40357
rect 11200 40354 12000 40384
rect 10041 40352 12000 40354
rect 10041 40296 10046 40352
rect 10102 40296 12000 40352
rect 10041 40294 12000 40296
rect 10041 40291 10107 40294
rect 4208 40288 4528 40289
rect 0 40218 800 40248
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 7472 40288 7792 40289
rect 7472 40224 7480 40288
rect 7544 40224 7560 40288
rect 7624 40224 7640 40288
rect 7704 40224 7720 40288
rect 7784 40224 7792 40288
rect 11200 40264 12000 40294
rect 7472 40223 7792 40224
rect 3969 40218 4035 40221
rect 0 40216 4035 40218
rect 0 40160 3974 40216
rect 4030 40160 4035 40216
rect 0 40158 4035 40160
rect 0 40128 800 40158
rect 3969 40155 4035 40158
rect 2129 40082 2195 40085
rect 2262 40082 2268 40084
rect 2129 40080 2268 40082
rect 2129 40024 2134 40080
rect 2190 40024 2268 40080
rect 2129 40022 2268 40024
rect 2129 40019 2195 40022
rect 2262 40020 2268 40022
rect 2332 40020 2338 40084
rect 2773 40082 2839 40085
rect 3182 40082 3188 40084
rect 2773 40080 3188 40082
rect 2773 40024 2778 40080
rect 2834 40024 3188 40080
rect 2773 40022 3188 40024
rect 2773 40019 2839 40022
rect 3182 40020 3188 40022
rect 3252 40020 3258 40084
rect 105 39946 171 39949
rect 238 39946 244 39948
rect 105 39944 244 39946
rect 105 39888 110 39944
rect 166 39888 244 39944
rect 105 39886 244 39888
rect 105 39883 171 39886
rect 238 39884 244 39886
rect 308 39884 314 39948
rect 422 39884 428 39948
rect 492 39946 498 39948
rect 657 39946 723 39949
rect 492 39944 723 39946
rect 492 39888 662 39944
rect 718 39888 723 39944
rect 492 39886 723 39888
rect 492 39884 498 39886
rect 657 39883 723 39886
rect 2865 39946 2931 39949
rect 3550 39946 3556 39948
rect 2865 39944 3556 39946
rect 2865 39888 2870 39944
rect 2926 39888 3556 39944
rect 2865 39886 3556 39888
rect 2865 39883 2931 39886
rect 3550 39884 3556 39886
rect 3620 39884 3626 39948
rect 2576 39744 2896 39745
rect 0 39674 800 39704
rect 2576 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2576 39679 2896 39680
rect 5840 39744 6160 39745
rect 5840 39680 5848 39744
rect 5912 39680 5928 39744
rect 5992 39680 6008 39744
rect 6072 39680 6088 39744
rect 6152 39680 6160 39744
rect 5840 39679 6160 39680
rect 9104 39744 9424 39745
rect 9104 39680 9112 39744
rect 9176 39680 9192 39744
rect 9256 39680 9272 39744
rect 9336 39680 9352 39744
rect 9416 39680 9424 39744
rect 9104 39679 9424 39680
rect 0 39614 1410 39674
rect 0 39584 800 39614
rect 1350 39538 1410 39614
rect 3969 39538 4035 39541
rect 1350 39536 4035 39538
rect 1350 39480 3974 39536
rect 4030 39480 4035 39536
rect 1350 39478 4035 39480
rect 3969 39475 4035 39478
rect 10041 39538 10107 39541
rect 11200 39538 12000 39568
rect 10041 39536 12000 39538
rect 10041 39480 10046 39536
rect 10102 39480 12000 39536
rect 10041 39478 12000 39480
rect 10041 39475 10107 39478
rect 11200 39448 12000 39478
rect 0 39266 800 39296
rect 3969 39266 4035 39269
rect 0 39264 4035 39266
rect 0 39208 3974 39264
rect 4030 39208 4035 39264
rect 0 39206 4035 39208
rect 0 39176 800 39206
rect 3969 39203 4035 39206
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 7472 39200 7792 39201
rect 7472 39136 7480 39200
rect 7544 39136 7560 39200
rect 7624 39136 7640 39200
rect 7704 39136 7720 39200
rect 7784 39136 7792 39200
rect 7472 39135 7792 39136
rect 2262 39068 2268 39132
rect 2332 39130 2338 39132
rect 2998 39130 3004 39132
rect 2332 39070 3004 39130
rect 2332 39068 2338 39070
rect 2998 39068 3004 39070
rect 3068 39068 3074 39132
rect 3049 38994 3115 38997
rect 3182 38994 3188 38996
rect 3049 38992 3188 38994
rect 3049 38936 3054 38992
rect 3110 38936 3188 38992
rect 3049 38934 3188 38936
rect 3049 38931 3115 38934
rect 3182 38932 3188 38934
rect 3252 38932 3258 38996
rect 3734 38932 3740 38996
rect 3804 38994 3810 38996
rect 4153 38994 4219 38997
rect 3804 38992 4219 38994
rect 3804 38936 4158 38992
rect 4214 38936 4219 38992
rect 3804 38934 4219 38936
rect 3804 38932 3810 38934
rect 4153 38931 4219 38934
rect 0 38858 800 38888
rect 1577 38858 1643 38861
rect 0 38856 1643 38858
rect 0 38800 1582 38856
rect 1638 38800 1643 38856
rect 0 38798 1643 38800
rect 0 38768 800 38798
rect 1577 38795 1643 38798
rect 2865 38858 2931 38861
rect 2998 38858 3004 38860
rect 2865 38856 3004 38858
rect 2865 38800 2870 38856
rect 2926 38800 3004 38856
rect 2865 38798 3004 38800
rect 2865 38795 2931 38798
rect 2998 38796 3004 38798
rect 3068 38796 3074 38860
rect 3969 38858 4035 38861
rect 5206 38858 5212 38860
rect 3969 38856 5212 38858
rect 3969 38800 3974 38856
rect 4030 38800 5212 38856
rect 3969 38798 5212 38800
rect 3969 38795 4035 38798
rect 5206 38796 5212 38798
rect 5276 38796 5282 38860
rect 10041 38722 10107 38725
rect 11200 38722 12000 38752
rect 10041 38720 12000 38722
rect 10041 38664 10046 38720
rect 10102 38664 12000 38720
rect 10041 38662 12000 38664
rect 10041 38659 10107 38662
rect 2576 38656 2896 38657
rect 2576 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2576 38591 2896 38592
rect 5840 38656 6160 38657
rect 5840 38592 5848 38656
rect 5912 38592 5928 38656
rect 5992 38592 6008 38656
rect 6072 38592 6088 38656
rect 6152 38592 6160 38656
rect 5840 38591 6160 38592
rect 9104 38656 9424 38657
rect 9104 38592 9112 38656
rect 9176 38592 9192 38656
rect 9256 38592 9272 38656
rect 9336 38592 9352 38656
rect 9416 38592 9424 38656
rect 11200 38632 12000 38662
rect 9104 38591 9424 38592
rect 0 38450 800 38480
rect 3693 38450 3759 38453
rect 0 38448 3759 38450
rect 0 38392 3698 38448
rect 3754 38392 3759 38448
rect 0 38390 3759 38392
rect 0 38360 800 38390
rect 3693 38387 3759 38390
rect 2773 38314 2839 38317
rect 4337 38314 4403 38317
rect 5206 38314 5212 38316
rect 2773 38312 5212 38314
rect 2773 38256 2778 38312
rect 2834 38256 4342 38312
rect 4398 38256 5212 38312
rect 2773 38254 5212 38256
rect 2773 38251 2839 38254
rect 4337 38251 4403 38254
rect 5206 38252 5212 38254
rect 5276 38252 5282 38316
rect 1894 38116 1900 38180
rect 1964 38178 1970 38180
rect 2589 38178 2655 38181
rect 1964 38176 2655 38178
rect 1964 38120 2594 38176
rect 2650 38120 2655 38176
rect 1964 38118 2655 38120
rect 1964 38116 1970 38118
rect 2589 38115 2655 38118
rect 4208 38112 4528 38113
rect 0 38042 800 38072
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 7472 38112 7792 38113
rect 7472 38048 7480 38112
rect 7544 38048 7560 38112
rect 7624 38048 7640 38112
rect 7704 38048 7720 38112
rect 7784 38048 7792 38112
rect 7472 38047 7792 38048
rect 2957 38042 3023 38045
rect 0 38040 3023 38042
rect 0 37984 2962 38040
rect 3018 37984 3023 38040
rect 0 37982 3023 37984
rect 0 37952 800 37982
rect 2957 37979 3023 37982
rect 10041 38042 10107 38045
rect 11200 38042 12000 38072
rect 10041 38040 12000 38042
rect 10041 37984 10046 38040
rect 10102 37984 12000 38040
rect 10041 37982 12000 37984
rect 10041 37979 10107 37982
rect 11200 37952 12000 37982
rect 1025 37906 1091 37909
rect 3182 37906 3188 37908
rect 1025 37904 3188 37906
rect 1025 37848 1030 37904
rect 1086 37848 3188 37904
rect 1025 37846 3188 37848
rect 1025 37843 1091 37846
rect 3182 37844 3188 37846
rect 3252 37844 3258 37908
rect 1526 37708 1532 37772
rect 1596 37770 1602 37772
rect 3969 37770 4035 37773
rect 1596 37768 4035 37770
rect 1596 37712 3974 37768
rect 4030 37712 4035 37768
rect 1596 37710 4035 37712
rect 1596 37708 1602 37710
rect 3969 37707 4035 37710
rect 0 37634 800 37664
rect 1393 37634 1459 37637
rect 0 37632 1459 37634
rect 0 37576 1398 37632
rect 1454 37576 1459 37632
rect 0 37574 1459 37576
rect 0 37544 800 37574
rect 1393 37571 1459 37574
rect 2576 37568 2896 37569
rect 2576 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2576 37503 2896 37504
rect 5840 37568 6160 37569
rect 5840 37504 5848 37568
rect 5912 37504 5928 37568
rect 5992 37504 6008 37568
rect 6072 37504 6088 37568
rect 6152 37504 6160 37568
rect 5840 37503 6160 37504
rect 9104 37568 9424 37569
rect 9104 37504 9112 37568
rect 9176 37504 9192 37568
rect 9256 37504 9272 37568
rect 9336 37504 9352 37568
rect 9416 37504 9424 37568
rect 9104 37503 9424 37504
rect 2681 37362 2747 37365
rect 4654 37362 4660 37364
rect 2681 37360 4660 37362
rect 2681 37304 2686 37360
rect 2742 37304 4660 37360
rect 2681 37302 4660 37304
rect 2681 37299 2747 37302
rect 4654 37300 4660 37302
rect 4724 37300 4730 37364
rect 0 37226 800 37256
rect 3969 37226 4035 37229
rect 0 37224 4035 37226
rect 0 37168 3974 37224
rect 4030 37168 4035 37224
rect 0 37166 4035 37168
rect 0 37136 800 37166
rect 3969 37163 4035 37166
rect 10041 37226 10107 37229
rect 11200 37226 12000 37256
rect 10041 37224 12000 37226
rect 10041 37168 10046 37224
rect 10102 37168 12000 37224
rect 10041 37166 12000 37168
rect 10041 37163 10107 37166
rect 11200 37136 12000 37166
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 7472 37024 7792 37025
rect 7472 36960 7480 37024
rect 7544 36960 7560 37024
rect 7624 36960 7640 37024
rect 7704 36960 7720 37024
rect 7784 36960 7792 37024
rect 7472 36959 7792 36960
rect 5349 36954 5415 36957
rect 5349 36952 5642 36954
rect 5349 36896 5354 36952
rect 5410 36896 5642 36952
rect 5349 36894 5642 36896
rect 5349 36891 5415 36894
rect 4654 36756 4660 36820
rect 4724 36818 4730 36820
rect 5390 36818 5396 36820
rect 4724 36758 5396 36818
rect 4724 36756 4730 36758
rect 5390 36756 5396 36758
rect 5460 36756 5466 36820
rect 0 36682 800 36712
rect 3969 36682 4035 36685
rect 5349 36682 5415 36685
rect 0 36680 4035 36682
rect 0 36624 3974 36680
rect 4030 36624 4035 36680
rect 0 36622 4035 36624
rect 0 36592 800 36622
rect 3969 36619 4035 36622
rect 5030 36680 5415 36682
rect 5030 36624 5354 36680
rect 5410 36624 5415 36680
rect 5030 36622 5415 36624
rect 2576 36480 2896 36481
rect 2576 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2576 36415 2896 36416
rect 0 36274 800 36304
rect 5030 36277 5090 36622
rect 5349 36619 5415 36622
rect 5582 36413 5642 36894
rect 5840 36480 6160 36481
rect 5840 36416 5848 36480
rect 5912 36416 5928 36480
rect 5992 36416 6008 36480
rect 6072 36416 6088 36480
rect 6152 36416 6160 36480
rect 5840 36415 6160 36416
rect 9104 36480 9424 36481
rect 9104 36416 9112 36480
rect 9176 36416 9192 36480
rect 9256 36416 9272 36480
rect 9336 36416 9352 36480
rect 9416 36416 9424 36480
rect 9104 36415 9424 36416
rect 5533 36408 5642 36413
rect 5533 36352 5538 36408
rect 5594 36352 5642 36408
rect 5533 36350 5642 36352
rect 10041 36410 10107 36413
rect 11200 36410 12000 36440
rect 10041 36408 12000 36410
rect 10041 36352 10046 36408
rect 10102 36352 12000 36408
rect 10041 36350 12000 36352
rect 5533 36347 5599 36350
rect 10041 36347 10107 36350
rect 11200 36320 12000 36350
rect 3785 36274 3851 36277
rect 0 36272 3851 36274
rect 0 36216 3790 36272
rect 3846 36216 3851 36272
rect 0 36214 3851 36216
rect 0 36184 800 36214
rect 3785 36211 3851 36214
rect 4981 36272 5090 36277
rect 4981 36216 4986 36272
rect 5042 36216 5090 36272
rect 4981 36214 5090 36216
rect 4981 36211 5047 36214
rect 4153 36138 4219 36141
rect 5206 36138 5212 36140
rect 4153 36136 5212 36138
rect 4153 36080 4158 36136
rect 4214 36080 5212 36136
rect 4153 36078 5212 36080
rect 4153 36075 4219 36078
rect 5206 36076 5212 36078
rect 5276 36076 5282 36140
rect 4208 35936 4528 35937
rect 0 35866 800 35896
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 7472 35936 7792 35937
rect 7472 35872 7480 35936
rect 7544 35872 7560 35936
rect 7624 35872 7640 35936
rect 7704 35872 7720 35936
rect 7784 35872 7792 35936
rect 7472 35871 7792 35872
rect 2773 35866 2839 35869
rect 0 35864 2839 35866
rect 0 35808 2778 35864
rect 2834 35808 2839 35864
rect 0 35806 2839 35808
rect 0 35776 800 35806
rect 2773 35803 2839 35806
rect 3693 35866 3759 35869
rect 3969 35866 4035 35869
rect 3693 35864 4035 35866
rect 3693 35808 3698 35864
rect 3754 35808 3974 35864
rect 4030 35808 4035 35864
rect 3693 35806 4035 35808
rect 3693 35803 3759 35806
rect 3969 35803 4035 35806
rect 10041 35730 10107 35733
rect 11200 35730 12000 35760
rect 10041 35728 12000 35730
rect 10041 35672 10046 35728
rect 10102 35672 12000 35728
rect 10041 35670 12000 35672
rect 10041 35667 10107 35670
rect 11200 35640 12000 35670
rect 0 35458 800 35488
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35368 800 35398
rect 1577 35395 1643 35398
rect 2576 35392 2896 35393
rect 2576 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2576 35327 2896 35328
rect 5840 35392 6160 35393
rect 5840 35328 5848 35392
rect 5912 35328 5928 35392
rect 5992 35328 6008 35392
rect 6072 35328 6088 35392
rect 6152 35328 6160 35392
rect 5840 35327 6160 35328
rect 9104 35392 9424 35393
rect 9104 35328 9112 35392
rect 9176 35328 9192 35392
rect 9256 35328 9272 35392
rect 9336 35328 9352 35392
rect 9416 35328 9424 35392
rect 9104 35327 9424 35328
rect 0 35050 800 35080
rect 1485 35050 1551 35053
rect 0 35048 1551 35050
rect 0 34992 1490 35048
rect 1546 34992 1551 35048
rect 0 34990 1551 34992
rect 0 34960 800 34990
rect 1485 34987 1551 34990
rect 1669 34916 1735 34917
rect 1669 34912 1716 34916
rect 1780 34914 1786 34916
rect 10041 34914 10107 34917
rect 11200 34914 12000 34944
rect 1669 34856 1674 34912
rect 1669 34852 1716 34856
rect 1780 34854 1826 34914
rect 10041 34912 12000 34914
rect 10041 34856 10046 34912
rect 10102 34856 12000 34912
rect 10041 34854 12000 34856
rect 1780 34852 1786 34854
rect 1669 34851 1735 34852
rect 10041 34851 10107 34854
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 7472 34848 7792 34849
rect 7472 34784 7480 34848
rect 7544 34784 7560 34848
rect 7624 34784 7640 34848
rect 7704 34784 7720 34848
rect 7784 34784 7792 34848
rect 11200 34824 12000 34854
rect 7472 34783 7792 34784
rect 0 34642 800 34672
rect 1577 34642 1643 34645
rect 0 34640 1643 34642
rect 0 34584 1582 34640
rect 1638 34584 1643 34640
rect 0 34582 1643 34584
rect 0 34552 800 34582
rect 1577 34579 1643 34582
rect 2576 34304 2896 34305
rect 0 34234 800 34264
rect 2576 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2576 34239 2896 34240
rect 5840 34304 6160 34305
rect 5840 34240 5848 34304
rect 5912 34240 5928 34304
rect 5992 34240 6008 34304
rect 6072 34240 6088 34304
rect 6152 34240 6160 34304
rect 5840 34239 6160 34240
rect 9104 34304 9424 34305
rect 9104 34240 9112 34304
rect 9176 34240 9192 34304
rect 9256 34240 9272 34304
rect 9336 34240 9352 34304
rect 9416 34240 9424 34304
rect 9104 34239 9424 34240
rect 2313 34234 2379 34237
rect 0 34232 2379 34234
rect 0 34176 2318 34232
rect 2374 34176 2379 34232
rect 0 34174 2379 34176
rect 0 34144 800 34174
rect 2313 34171 2379 34174
rect 9581 34098 9647 34101
rect 11200 34098 12000 34128
rect 9581 34096 12000 34098
rect 9581 34040 9586 34096
rect 9642 34040 12000 34096
rect 9581 34038 12000 34040
rect 9581 34035 9647 34038
rect 11200 34008 12000 34038
rect 0 33826 800 33856
rect 3049 33826 3115 33829
rect 0 33824 3115 33826
rect 0 33768 3054 33824
rect 3110 33768 3115 33824
rect 0 33766 3115 33768
rect 0 33736 800 33766
rect 3049 33763 3115 33766
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 7472 33760 7792 33761
rect 7472 33696 7480 33760
rect 7544 33696 7560 33760
rect 7624 33696 7640 33760
rect 7704 33696 7720 33760
rect 7784 33696 7792 33760
rect 7472 33695 7792 33696
rect 2405 33554 2471 33557
rect 3049 33554 3115 33557
rect 2405 33552 3115 33554
rect 2405 33496 2410 33552
rect 2466 33496 3054 33552
rect 3110 33496 3115 33552
rect 2405 33494 3115 33496
rect 2405 33491 2471 33494
rect 3049 33491 3115 33494
rect 10041 33418 10107 33421
rect 11200 33418 12000 33448
rect 10041 33416 12000 33418
rect 10041 33360 10046 33416
rect 10102 33360 12000 33416
rect 10041 33358 12000 33360
rect 10041 33355 10107 33358
rect 11200 33328 12000 33358
rect 0 33282 800 33312
rect 2221 33282 2287 33285
rect 0 33280 2287 33282
rect 0 33224 2226 33280
rect 2282 33224 2287 33280
rect 0 33222 2287 33224
rect 0 33192 800 33222
rect 2221 33219 2287 33222
rect 2576 33216 2896 33217
rect 2576 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2576 33151 2896 33152
rect 5840 33216 6160 33217
rect 5840 33152 5848 33216
rect 5912 33152 5928 33216
rect 5992 33152 6008 33216
rect 6072 33152 6088 33216
rect 6152 33152 6160 33216
rect 5840 33151 6160 33152
rect 9104 33216 9424 33217
rect 9104 33152 9112 33216
rect 9176 33152 9192 33216
rect 9256 33152 9272 33216
rect 9336 33152 9352 33216
rect 9416 33152 9424 33216
rect 9104 33151 9424 33152
rect 3550 32948 3556 33012
rect 3620 33010 3626 33012
rect 4521 33010 4587 33013
rect 3620 33008 4587 33010
rect 3620 32952 4526 33008
rect 4582 32952 4587 33008
rect 3620 32950 4587 32952
rect 3620 32948 3626 32950
rect 4521 32947 4587 32950
rect 0 32874 800 32904
rect 3693 32874 3759 32877
rect 0 32872 3759 32874
rect 0 32816 3698 32872
rect 3754 32816 3759 32872
rect 0 32814 3759 32816
rect 0 32784 800 32814
rect 3693 32811 3759 32814
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 7472 32672 7792 32673
rect 7472 32608 7480 32672
rect 7544 32608 7560 32672
rect 7624 32608 7640 32672
rect 7704 32608 7720 32672
rect 7784 32608 7792 32672
rect 7472 32607 7792 32608
rect 10041 32602 10107 32605
rect 11200 32602 12000 32632
rect 10041 32600 12000 32602
rect 10041 32544 10046 32600
rect 10102 32544 12000 32600
rect 10041 32542 12000 32544
rect 10041 32539 10107 32542
rect 11200 32512 12000 32542
rect 0 32466 800 32496
rect 3969 32466 4035 32469
rect 0 32464 4035 32466
rect 0 32408 3974 32464
rect 4030 32408 4035 32464
rect 0 32406 4035 32408
rect 0 32376 800 32406
rect 3969 32403 4035 32406
rect 4521 32466 4587 32469
rect 5206 32466 5212 32468
rect 4521 32464 5212 32466
rect 4521 32408 4526 32464
rect 4582 32408 5212 32464
rect 4521 32406 5212 32408
rect 4521 32403 4587 32406
rect 5206 32404 5212 32406
rect 5276 32404 5282 32468
rect 1393 32330 1459 32333
rect 3509 32330 3575 32333
rect 1393 32328 1594 32330
rect 1393 32272 1398 32328
rect 1454 32272 1594 32328
rect 1393 32270 1594 32272
rect 1393 32267 1459 32270
rect 0 32058 800 32088
rect 1534 32061 1594 32270
rect 3509 32328 3618 32330
rect 3509 32272 3514 32328
rect 3570 32272 3618 32328
rect 3509 32267 3618 32272
rect 1945 32196 2011 32197
rect 1894 32132 1900 32196
rect 1964 32194 2011 32196
rect 1964 32192 2056 32194
rect 2006 32136 2056 32192
rect 1964 32134 2056 32136
rect 1964 32132 2011 32134
rect 3182 32132 3188 32196
rect 3252 32194 3258 32196
rect 3417 32194 3483 32197
rect 3252 32192 3483 32194
rect 3252 32136 3422 32192
rect 3478 32136 3483 32192
rect 3252 32134 3483 32136
rect 3252 32132 3258 32134
rect 1945 32131 2011 32132
rect 3417 32131 3483 32134
rect 2576 32128 2896 32129
rect 2576 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2576 32063 2896 32064
rect 0 31998 1410 32058
rect 1534 32056 1643 32061
rect 1534 32000 1582 32056
rect 1638 32000 1643 32056
rect 1534 31998 1643 32000
rect 0 31968 800 31998
rect 1350 31922 1410 31998
rect 1577 31995 1643 31998
rect 3049 32058 3115 32061
rect 3182 32058 3188 32060
rect 3049 32056 3188 32058
rect 3049 32000 3054 32056
rect 3110 32000 3188 32056
rect 3049 31998 3188 32000
rect 3049 31995 3115 31998
rect 3182 31996 3188 31998
rect 3252 31996 3258 32060
rect 3558 32058 3618 32267
rect 3734 32132 3740 32196
rect 3804 32194 3810 32196
rect 3804 32134 4170 32194
rect 3804 32132 3810 32134
rect 3734 32058 3740 32060
rect 3558 31998 3740 32058
rect 3734 31996 3740 31998
rect 3804 31996 3810 32060
rect 3969 31922 4035 31925
rect 1350 31920 4035 31922
rect 1350 31864 3974 31920
rect 4030 31864 4035 31920
rect 1350 31862 4035 31864
rect 3969 31859 4035 31862
rect 3877 31786 3943 31789
rect 4110 31786 4170 32134
rect 5840 32128 6160 32129
rect 5840 32064 5848 32128
rect 5912 32064 5928 32128
rect 5992 32064 6008 32128
rect 6072 32064 6088 32128
rect 6152 32064 6160 32128
rect 5840 32063 6160 32064
rect 9104 32128 9424 32129
rect 9104 32064 9112 32128
rect 9176 32064 9192 32128
rect 9256 32064 9272 32128
rect 9336 32064 9352 32128
rect 9416 32064 9424 32128
rect 9104 32063 9424 32064
rect 4705 32058 4771 32061
rect 5206 32058 5212 32060
rect 4705 32056 5212 32058
rect 4705 32000 4710 32056
rect 4766 32000 5212 32056
rect 4705 31998 5212 32000
rect 4705 31995 4771 31998
rect 5206 31996 5212 31998
rect 5276 31996 5282 32060
rect 3877 31784 4170 31786
rect 3877 31728 3882 31784
rect 3938 31728 4170 31784
rect 3877 31726 4170 31728
rect 4981 31786 5047 31789
rect 5390 31786 5396 31788
rect 4981 31784 5396 31786
rect 4981 31728 4986 31784
rect 5042 31728 5396 31784
rect 4981 31726 5396 31728
rect 3877 31723 3943 31726
rect 4981 31723 5047 31726
rect 5390 31724 5396 31726
rect 5460 31724 5466 31788
rect 10041 31786 10107 31789
rect 11200 31786 12000 31816
rect 10041 31784 12000 31786
rect 10041 31728 10046 31784
rect 10102 31728 12000 31784
rect 10041 31726 12000 31728
rect 10041 31723 10107 31726
rect 11200 31696 12000 31726
rect 0 31650 800 31680
rect 3325 31650 3391 31653
rect 5257 31650 5323 31653
rect 0 31648 3391 31650
rect 0 31592 3330 31648
rect 3386 31592 3391 31648
rect 0 31590 3391 31592
rect 0 31560 800 31590
rect 3325 31587 3391 31590
rect 4708 31648 5323 31650
rect 4708 31592 5262 31648
rect 5318 31592 5323 31648
rect 4708 31590 5323 31592
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 2998 31452 3004 31516
rect 3068 31514 3074 31516
rect 3325 31514 3391 31517
rect 3068 31512 3391 31514
rect 3068 31456 3330 31512
rect 3386 31456 3391 31512
rect 3068 31454 3391 31456
rect 3068 31452 3074 31454
rect 3325 31451 3391 31454
rect 3734 31452 3740 31516
rect 3804 31514 3810 31516
rect 3877 31514 3943 31517
rect 3804 31512 3943 31514
rect 3804 31456 3882 31512
rect 3938 31456 3943 31512
rect 3804 31454 3943 31456
rect 3804 31452 3810 31454
rect 3877 31451 3943 31454
rect 1894 31316 1900 31380
rect 1964 31378 1970 31380
rect 2129 31378 2195 31381
rect 1964 31376 2195 31378
rect 1964 31320 2134 31376
rect 2190 31320 2195 31376
rect 1964 31318 2195 31320
rect 1964 31316 1970 31318
rect 2129 31315 2195 31318
rect 2773 31378 2839 31381
rect 2998 31378 3004 31380
rect 2773 31376 3004 31378
rect 2773 31320 2778 31376
rect 2834 31320 3004 31376
rect 2773 31318 3004 31320
rect 2773 31315 2839 31318
rect 2998 31316 3004 31318
rect 3068 31316 3074 31380
rect 4153 31378 4219 31381
rect 4708 31378 4768 31590
rect 5257 31587 5323 31590
rect 7472 31584 7792 31585
rect 7472 31520 7480 31584
rect 7544 31520 7560 31584
rect 7624 31520 7640 31584
rect 7704 31520 7720 31584
rect 7784 31520 7792 31584
rect 7472 31519 7792 31520
rect 4153 31376 4768 31378
rect 4153 31320 4158 31376
rect 4214 31320 4768 31376
rect 4153 31318 4768 31320
rect 4153 31315 4219 31318
rect 0 31242 800 31272
rect 3601 31242 3667 31245
rect 0 31240 3667 31242
rect 0 31184 3606 31240
rect 3662 31184 3667 31240
rect 0 31182 3667 31184
rect 0 31152 800 31182
rect 3601 31179 3667 31182
rect 974 31044 980 31108
rect 1044 31106 1050 31108
rect 2313 31106 2379 31109
rect 1044 31104 2379 31106
rect 1044 31048 2318 31104
rect 2374 31048 2379 31104
rect 1044 31046 2379 31048
rect 1044 31044 1050 31046
rect 2313 31043 2379 31046
rect 10041 31106 10107 31109
rect 11200 31106 12000 31136
rect 10041 31104 12000 31106
rect 10041 31048 10046 31104
rect 10102 31048 12000 31104
rect 10041 31046 12000 31048
rect 10041 31043 10107 31046
rect 2576 31040 2896 31041
rect 2576 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2576 30975 2896 30976
rect 5840 31040 6160 31041
rect 5840 30976 5848 31040
rect 5912 30976 5928 31040
rect 5992 30976 6008 31040
rect 6072 30976 6088 31040
rect 6152 30976 6160 31040
rect 5840 30975 6160 30976
rect 9104 31040 9424 31041
rect 9104 30976 9112 31040
rect 9176 30976 9192 31040
rect 9256 30976 9272 31040
rect 9336 30976 9352 31040
rect 9416 30976 9424 31040
rect 11200 31016 12000 31046
rect 9104 30975 9424 30976
rect 3734 30908 3740 30972
rect 3804 30970 3810 30972
rect 3969 30970 4035 30973
rect 3804 30968 4035 30970
rect 3804 30912 3974 30968
rect 4030 30912 4035 30968
rect 3804 30910 4035 30912
rect 3804 30908 3810 30910
rect 3969 30907 4035 30910
rect 0 30834 800 30864
rect 2957 30834 3023 30837
rect 0 30832 3023 30834
rect 0 30776 2962 30832
rect 3018 30776 3023 30832
rect 0 30774 3023 30776
rect 0 30744 800 30774
rect 2957 30771 3023 30774
rect 1526 30636 1532 30700
rect 1596 30698 1602 30700
rect 3601 30698 3667 30701
rect 1596 30696 3667 30698
rect 1596 30640 3606 30696
rect 3662 30640 3667 30696
rect 1596 30638 3667 30640
rect 1596 30636 1602 30638
rect 3601 30635 3667 30638
rect 1342 30500 1348 30564
rect 1412 30562 1418 30564
rect 3141 30562 3207 30565
rect 1412 30560 3207 30562
rect 1412 30504 3146 30560
rect 3202 30504 3207 30560
rect 1412 30502 3207 30504
rect 1412 30500 1418 30502
rect 3141 30499 3207 30502
rect 4208 30496 4528 30497
rect 0 30426 800 30456
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 7472 30496 7792 30497
rect 7472 30432 7480 30496
rect 7544 30432 7560 30496
rect 7624 30432 7640 30496
rect 7704 30432 7720 30496
rect 7784 30432 7792 30496
rect 7472 30431 7792 30432
rect 2773 30426 2839 30429
rect 0 30424 2839 30426
rect 0 30368 2778 30424
rect 2834 30368 2839 30424
rect 0 30366 2839 30368
rect 0 30336 800 30366
rect 2773 30363 2839 30366
rect 3049 30426 3115 30429
rect 3366 30426 3372 30428
rect 3049 30424 3372 30426
rect 3049 30368 3054 30424
rect 3110 30368 3372 30424
rect 3049 30366 3372 30368
rect 3049 30363 3115 30366
rect 3366 30364 3372 30366
rect 3436 30364 3442 30428
rect 1158 30228 1164 30292
rect 1228 30290 1234 30292
rect 2589 30290 2655 30293
rect 1228 30288 2655 30290
rect 1228 30232 2594 30288
rect 2650 30232 2655 30288
rect 1228 30230 2655 30232
rect 1228 30228 1234 30230
rect 2589 30227 2655 30230
rect 10041 30290 10107 30293
rect 11200 30290 12000 30320
rect 10041 30288 12000 30290
rect 10041 30232 10046 30288
rect 10102 30232 12000 30288
rect 10041 30230 12000 30232
rect 10041 30227 10107 30230
rect 11200 30200 12000 30230
rect 1526 29956 1532 30020
rect 1596 30018 1602 30020
rect 2037 30018 2103 30021
rect 1596 30016 2103 30018
rect 1596 29960 2042 30016
rect 2098 29960 2103 30016
rect 1596 29958 2103 29960
rect 1596 29956 1602 29958
rect 2037 29955 2103 29958
rect 2576 29952 2896 29953
rect 0 29882 800 29912
rect 2576 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2576 29887 2896 29888
rect 5840 29952 6160 29953
rect 5840 29888 5848 29952
rect 5912 29888 5928 29952
rect 5992 29888 6008 29952
rect 6072 29888 6088 29952
rect 6152 29888 6160 29952
rect 5840 29887 6160 29888
rect 9104 29952 9424 29953
rect 9104 29888 9112 29952
rect 9176 29888 9192 29952
rect 9256 29888 9272 29952
rect 9336 29888 9352 29952
rect 9416 29888 9424 29952
rect 9104 29887 9424 29888
rect 1485 29882 1551 29885
rect 2037 29884 2103 29885
rect 2037 29882 2084 29884
rect 0 29880 1551 29882
rect 0 29824 1490 29880
rect 1546 29824 1551 29880
rect 0 29822 1551 29824
rect 1992 29880 2084 29882
rect 1992 29824 2042 29880
rect 1992 29822 2084 29824
rect 0 29792 800 29822
rect 1485 29819 1551 29822
rect 2037 29820 2084 29822
rect 2148 29820 2154 29884
rect 2037 29819 2103 29820
rect 0 29474 800 29504
rect 1853 29474 1919 29477
rect 0 29472 1919 29474
rect 0 29416 1858 29472
rect 1914 29416 1919 29472
rect 0 29414 1919 29416
rect 0 29384 800 29414
rect 1853 29411 1919 29414
rect 10133 29474 10199 29477
rect 11200 29474 12000 29504
rect 10133 29472 12000 29474
rect 10133 29416 10138 29472
rect 10194 29416 12000 29472
rect 10133 29414 12000 29416
rect 10133 29411 10199 29414
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 7472 29408 7792 29409
rect 7472 29344 7480 29408
rect 7544 29344 7560 29408
rect 7624 29344 7640 29408
rect 7704 29344 7720 29408
rect 7784 29344 7792 29408
rect 11200 29384 12000 29414
rect 7472 29343 7792 29344
rect 1853 29338 1919 29341
rect 2262 29338 2268 29340
rect 1853 29336 2268 29338
rect 1853 29280 1858 29336
rect 1914 29280 2268 29336
rect 1853 29278 2268 29280
rect 1853 29275 1919 29278
rect 2262 29276 2268 29278
rect 2332 29276 2338 29340
rect 0 29066 800 29096
rect 4061 29066 4127 29069
rect 0 29064 4127 29066
rect 0 29008 4066 29064
rect 4122 29008 4127 29064
rect 0 29006 4127 29008
rect 0 28976 800 29006
rect 4061 29003 4127 29006
rect 1945 28932 2011 28933
rect 2129 28932 2195 28933
rect 1894 28930 1900 28932
rect 1854 28870 1900 28930
rect 1964 28928 2011 28932
rect 2006 28872 2011 28928
rect 1894 28868 1900 28870
rect 1964 28868 2011 28872
rect 2078 28868 2084 28932
rect 2148 28930 2195 28932
rect 2313 28930 2379 28933
rect 2148 28928 2240 28930
rect 2190 28872 2240 28928
rect 2148 28870 2240 28872
rect 2313 28928 2514 28930
rect 2313 28872 2318 28928
rect 2374 28872 2514 28928
rect 2313 28870 2514 28872
rect 2148 28868 2195 28870
rect 1945 28867 2011 28868
rect 2129 28867 2195 28868
rect 2313 28867 2379 28870
rect 933 28794 999 28797
rect 2313 28794 2379 28797
rect 933 28792 2379 28794
rect 933 28736 938 28792
rect 994 28736 2318 28792
rect 2374 28736 2379 28792
rect 933 28734 2379 28736
rect 933 28731 999 28734
rect 2313 28731 2379 28734
rect 0 28658 800 28688
rect 1761 28658 1827 28661
rect 0 28656 1827 28658
rect 0 28600 1766 28656
rect 1822 28600 1827 28656
rect 0 28598 1827 28600
rect 0 28568 800 28598
rect 1761 28595 1827 28598
rect 2129 28522 2195 28525
rect 2262 28522 2268 28524
rect 2129 28520 2268 28522
rect 2129 28464 2134 28520
rect 2190 28464 2268 28520
rect 2129 28462 2268 28464
rect 2129 28459 2195 28462
rect 2262 28460 2268 28462
rect 2332 28460 2338 28524
rect 2221 28386 2287 28389
rect 2454 28386 2514 28870
rect 2576 28864 2896 28865
rect 2576 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2576 28799 2896 28800
rect 5840 28864 6160 28865
rect 5840 28800 5848 28864
rect 5912 28800 5928 28864
rect 5992 28800 6008 28864
rect 6072 28800 6088 28864
rect 6152 28800 6160 28864
rect 5840 28799 6160 28800
rect 9104 28864 9424 28865
rect 9104 28800 9112 28864
rect 9176 28800 9192 28864
rect 9256 28800 9272 28864
rect 9336 28800 9352 28864
rect 9416 28800 9424 28864
rect 9104 28799 9424 28800
rect 10133 28794 10199 28797
rect 11200 28794 12000 28824
rect 10133 28792 12000 28794
rect 10133 28736 10138 28792
rect 10194 28736 12000 28792
rect 10133 28734 12000 28736
rect 10133 28731 10199 28734
rect 11200 28704 12000 28734
rect 2589 28658 2655 28661
rect 2998 28658 3004 28660
rect 2589 28656 3004 28658
rect 2589 28600 2594 28656
rect 2650 28600 3004 28656
rect 2589 28598 3004 28600
rect 2589 28595 2655 28598
rect 2998 28596 3004 28598
rect 3068 28596 3074 28660
rect 2221 28384 2514 28386
rect 2221 28328 2226 28384
rect 2282 28328 2514 28384
rect 2221 28326 2514 28328
rect 2221 28323 2287 28326
rect 4208 28320 4528 28321
rect 0 28250 800 28280
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 7472 28320 7792 28321
rect 7472 28256 7480 28320
rect 7544 28256 7560 28320
rect 7624 28256 7640 28320
rect 7704 28256 7720 28320
rect 7784 28256 7792 28320
rect 7472 28255 7792 28256
rect 1485 28250 1551 28253
rect 0 28248 1551 28250
rect 0 28192 1490 28248
rect 1546 28192 1551 28248
rect 0 28190 1551 28192
rect 0 28160 800 28190
rect 1485 28187 1551 28190
rect 1894 28188 1900 28252
rect 1964 28250 1970 28252
rect 2129 28250 2195 28253
rect 1964 28248 2195 28250
rect 1964 28192 2134 28248
rect 2190 28192 2195 28248
rect 1964 28190 2195 28192
rect 1964 28188 1970 28190
rect 2129 28187 2195 28190
rect 1485 28116 1551 28117
rect 1485 28112 1532 28116
rect 1596 28114 1602 28116
rect 1945 28114 2011 28117
rect 5574 28114 5580 28116
rect 1485 28056 1490 28112
rect 1485 28052 1532 28056
rect 1596 28054 1642 28114
rect 1945 28112 5580 28114
rect 1945 28056 1950 28112
rect 2006 28056 5580 28112
rect 1945 28054 5580 28056
rect 1596 28052 1602 28054
rect 1485 28051 1551 28052
rect 1945 28051 2011 28054
rect 5574 28052 5580 28054
rect 5644 28052 5650 28116
rect 1945 27978 2011 27981
rect 2078 27978 2084 27980
rect 1945 27976 2084 27978
rect 1945 27920 1950 27976
rect 2006 27920 2084 27976
rect 1945 27918 2084 27920
rect 1945 27915 2011 27918
rect 2078 27916 2084 27918
rect 2148 27916 2154 27980
rect 3049 27978 3115 27981
rect 3550 27978 3556 27980
rect 3049 27976 3556 27978
rect 3049 27920 3054 27976
rect 3110 27920 3556 27976
rect 3049 27918 3556 27920
rect 3049 27915 3115 27918
rect 3550 27916 3556 27918
rect 3620 27916 3626 27980
rect 9949 27978 10015 27981
rect 11200 27978 12000 28008
rect 9949 27976 12000 27978
rect 9949 27920 9954 27976
rect 10010 27920 12000 27976
rect 9949 27918 12000 27920
rect 9949 27915 10015 27918
rect 11200 27888 12000 27918
rect 0 27842 800 27872
rect 1393 27842 1459 27845
rect 0 27840 1459 27842
rect 0 27784 1398 27840
rect 1454 27784 1459 27840
rect 0 27782 1459 27784
rect 0 27752 800 27782
rect 1393 27779 1459 27782
rect 2576 27776 2896 27777
rect 2576 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2576 27711 2896 27712
rect 5840 27776 6160 27777
rect 5840 27712 5848 27776
rect 5912 27712 5928 27776
rect 5992 27712 6008 27776
rect 6072 27712 6088 27776
rect 6152 27712 6160 27776
rect 5840 27711 6160 27712
rect 9104 27776 9424 27777
rect 9104 27712 9112 27776
rect 9176 27712 9192 27776
rect 9256 27712 9272 27776
rect 9336 27712 9352 27776
rect 9416 27712 9424 27776
rect 9104 27711 9424 27712
rect 0 27434 800 27464
rect 1393 27434 1459 27437
rect 0 27432 1459 27434
rect 0 27376 1398 27432
rect 1454 27376 1459 27432
rect 0 27374 1459 27376
rect 0 27344 800 27374
rect 1393 27371 1459 27374
rect 3325 27434 3391 27437
rect 3734 27434 3740 27436
rect 3325 27432 3740 27434
rect 3325 27376 3330 27432
rect 3386 27376 3740 27432
rect 3325 27374 3740 27376
rect 3325 27371 3391 27374
rect 3734 27372 3740 27374
rect 3804 27372 3810 27436
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 7472 27232 7792 27233
rect 7472 27168 7480 27232
rect 7544 27168 7560 27232
rect 7624 27168 7640 27232
rect 7704 27168 7720 27232
rect 7784 27168 7792 27232
rect 7472 27167 7792 27168
rect 9949 27162 10015 27165
rect 11200 27162 12000 27192
rect 9949 27160 12000 27162
rect 9949 27104 9954 27160
rect 10010 27104 12000 27160
rect 9949 27102 12000 27104
rect 9949 27099 10015 27102
rect 11200 27072 12000 27102
rect 0 27026 800 27056
rect 2865 27026 2931 27029
rect 0 27024 2931 27026
rect 0 26968 2870 27024
rect 2926 26968 2931 27024
rect 0 26966 2931 26968
rect 0 26936 800 26966
rect 2865 26963 2931 26966
rect 4521 27026 4587 27029
rect 5206 27026 5212 27028
rect 4521 27024 5212 27026
rect 4521 26968 4526 27024
rect 4582 26968 5212 27024
rect 4521 26966 5212 26968
rect 4521 26963 4587 26966
rect 5206 26964 5212 26966
rect 5276 26964 5282 27028
rect 1669 26890 1735 26893
rect 6310 26890 6316 26892
rect 1669 26888 6316 26890
rect 1669 26832 1674 26888
rect 1730 26832 6316 26888
rect 1669 26830 6316 26832
rect 1669 26827 1735 26830
rect 6310 26828 6316 26830
rect 6380 26828 6386 26892
rect 2576 26688 2896 26689
rect 2576 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2576 26623 2896 26624
rect 5840 26688 6160 26689
rect 5840 26624 5848 26688
rect 5912 26624 5928 26688
rect 5992 26624 6008 26688
rect 6072 26624 6088 26688
rect 6152 26624 6160 26688
rect 5840 26623 6160 26624
rect 9104 26688 9424 26689
rect 9104 26624 9112 26688
rect 9176 26624 9192 26688
rect 9256 26624 9272 26688
rect 9336 26624 9352 26688
rect 9416 26624 9424 26688
rect 9104 26623 9424 26624
rect 0 26482 800 26512
rect 3049 26482 3115 26485
rect 0 26480 3115 26482
rect 0 26424 3054 26480
rect 3110 26424 3115 26480
rect 0 26422 3115 26424
rect 0 26392 800 26422
rect 3049 26419 3115 26422
rect 10133 26482 10199 26485
rect 11200 26482 12000 26512
rect 10133 26480 12000 26482
rect 10133 26424 10138 26480
rect 10194 26424 12000 26480
rect 10133 26422 12000 26424
rect 10133 26419 10199 26422
rect 11200 26392 12000 26422
rect 3141 26348 3207 26349
rect 3141 26344 3188 26348
rect 3252 26346 3258 26348
rect 3141 26288 3146 26344
rect 3141 26284 3188 26288
rect 3252 26286 3298 26346
rect 3252 26284 3258 26286
rect 3141 26283 3207 26284
rect 4208 26144 4528 26145
rect 0 26074 800 26104
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 7472 26144 7792 26145
rect 7472 26080 7480 26144
rect 7544 26080 7560 26144
rect 7624 26080 7640 26144
rect 7704 26080 7720 26144
rect 7784 26080 7792 26144
rect 7472 26079 7792 26080
rect 2589 26074 2655 26077
rect 0 26072 2655 26074
rect 0 26016 2594 26072
rect 2650 26016 2655 26072
rect 0 26014 2655 26016
rect 0 25984 800 26014
rect 2589 26011 2655 26014
rect 3325 25802 3391 25805
rect 3601 25804 3667 25805
rect 1396 25800 3391 25802
rect 1396 25744 3330 25800
rect 3386 25744 3391 25800
rect 1396 25742 3391 25744
rect 0 25666 800 25696
rect 1396 25666 1456 25742
rect 3325 25739 3391 25742
rect 3550 25740 3556 25804
rect 3620 25802 3667 25804
rect 3620 25800 3712 25802
rect 3662 25744 3712 25800
rect 3620 25742 3712 25744
rect 3620 25740 3667 25742
rect 3601 25739 3667 25740
rect 0 25606 1456 25666
rect 10133 25666 10199 25669
rect 11200 25666 12000 25696
rect 10133 25664 12000 25666
rect 10133 25608 10138 25664
rect 10194 25608 12000 25664
rect 10133 25606 12000 25608
rect 0 25576 800 25606
rect 10133 25603 10199 25606
rect 2576 25600 2896 25601
rect 2576 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2576 25535 2896 25536
rect 5840 25600 6160 25601
rect 5840 25536 5848 25600
rect 5912 25536 5928 25600
rect 5992 25536 6008 25600
rect 6072 25536 6088 25600
rect 6152 25536 6160 25600
rect 5840 25535 6160 25536
rect 9104 25600 9424 25601
rect 9104 25536 9112 25600
rect 9176 25536 9192 25600
rect 9256 25536 9272 25600
rect 9336 25536 9352 25600
rect 9416 25536 9424 25600
rect 11200 25576 12000 25606
rect 9104 25535 9424 25536
rect 0 25258 800 25288
rect 2957 25258 3023 25261
rect 0 25256 3023 25258
rect 0 25200 2962 25256
rect 3018 25200 3023 25256
rect 0 25198 3023 25200
rect 0 25168 800 25198
rect 2957 25195 3023 25198
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 7472 25056 7792 25057
rect 7472 24992 7480 25056
rect 7544 24992 7560 25056
rect 7624 24992 7640 25056
rect 7704 24992 7720 25056
rect 7784 24992 7792 25056
rect 7472 24991 7792 24992
rect 0 24850 800 24880
rect 3877 24850 3943 24853
rect 0 24848 3943 24850
rect 0 24792 3882 24848
rect 3938 24792 3943 24848
rect 0 24790 3943 24792
rect 0 24760 800 24790
rect 3877 24787 3943 24790
rect 10133 24850 10199 24853
rect 11200 24850 12000 24880
rect 10133 24848 12000 24850
rect 10133 24792 10138 24848
rect 10194 24792 12000 24848
rect 10133 24790 12000 24792
rect 10133 24787 10199 24790
rect 11200 24760 12000 24790
rect 2865 24714 2931 24717
rect 1396 24712 2931 24714
rect 1396 24656 2870 24712
rect 2926 24656 2931 24712
rect 1396 24654 2931 24656
rect 0 24442 800 24472
rect 1396 24442 1456 24654
rect 2865 24651 2931 24654
rect 2576 24512 2896 24513
rect 2576 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2576 24447 2896 24448
rect 5840 24512 6160 24513
rect 5840 24448 5848 24512
rect 5912 24448 5928 24512
rect 5992 24448 6008 24512
rect 6072 24448 6088 24512
rect 6152 24448 6160 24512
rect 5840 24447 6160 24448
rect 9104 24512 9424 24513
rect 9104 24448 9112 24512
rect 9176 24448 9192 24512
rect 9256 24448 9272 24512
rect 9336 24448 9352 24512
rect 9416 24448 9424 24512
rect 9104 24447 9424 24448
rect 0 24382 1456 24442
rect 0 24352 800 24382
rect 2262 24108 2268 24172
rect 2332 24170 2338 24172
rect 2405 24170 2471 24173
rect 2332 24168 2471 24170
rect 2332 24112 2410 24168
rect 2466 24112 2471 24168
rect 2332 24110 2471 24112
rect 2332 24108 2338 24110
rect 2405 24107 2471 24110
rect 10133 24170 10199 24173
rect 11200 24170 12000 24200
rect 10133 24168 12000 24170
rect 10133 24112 10138 24168
rect 10194 24112 12000 24168
rect 10133 24110 12000 24112
rect 10133 24107 10199 24110
rect 11200 24080 12000 24110
rect 0 24034 800 24064
rect 1853 24034 1919 24037
rect 0 24032 1919 24034
rect 0 23976 1858 24032
rect 1914 23976 1919 24032
rect 0 23974 1919 23976
rect 0 23944 800 23974
rect 1853 23971 1919 23974
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 7472 23968 7792 23969
rect 7472 23904 7480 23968
rect 7544 23904 7560 23968
rect 7624 23904 7640 23968
rect 7704 23904 7720 23968
rect 7784 23904 7792 23968
rect 7472 23903 7792 23904
rect 0 23626 800 23656
rect 1117 23626 1183 23629
rect 0 23624 1183 23626
rect 0 23568 1122 23624
rect 1178 23568 1183 23624
rect 0 23566 1183 23568
rect 0 23536 800 23566
rect 1117 23563 1183 23566
rect 2576 23424 2896 23425
rect 2576 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2576 23359 2896 23360
rect 5840 23424 6160 23425
rect 5840 23360 5848 23424
rect 5912 23360 5928 23424
rect 5992 23360 6008 23424
rect 6072 23360 6088 23424
rect 6152 23360 6160 23424
rect 5840 23359 6160 23360
rect 9104 23424 9424 23425
rect 9104 23360 9112 23424
rect 9176 23360 9192 23424
rect 9256 23360 9272 23424
rect 9336 23360 9352 23424
rect 9416 23360 9424 23424
rect 9104 23359 9424 23360
rect 10133 23354 10199 23357
rect 11200 23354 12000 23384
rect 10133 23352 12000 23354
rect 10133 23296 10138 23352
rect 10194 23296 12000 23352
rect 10133 23294 12000 23296
rect 10133 23291 10199 23294
rect 11200 23264 12000 23294
rect 0 23082 800 23112
rect 1393 23082 1459 23085
rect 0 23080 1459 23082
rect 0 23024 1398 23080
rect 1454 23024 1459 23080
rect 0 23022 1459 23024
rect 0 22992 800 23022
rect 1393 23019 1459 23022
rect 4889 22946 4955 22949
rect 4846 22944 4955 22946
rect 4846 22888 4894 22944
rect 4950 22888 4955 22944
rect 4846 22883 4955 22888
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 0 22674 800 22704
rect 4846 22677 4906 22883
rect 7472 22880 7792 22881
rect 7472 22816 7480 22880
rect 7544 22816 7560 22880
rect 7624 22816 7640 22880
rect 7704 22816 7720 22880
rect 7784 22816 7792 22880
rect 7472 22815 7792 22816
rect 3877 22674 3943 22677
rect 0 22672 3943 22674
rect 0 22616 3882 22672
rect 3938 22616 3943 22672
rect 0 22614 3943 22616
rect 4846 22672 4955 22677
rect 4846 22616 4894 22672
rect 4950 22616 4955 22672
rect 4846 22614 4955 22616
rect 0 22584 800 22614
rect 3877 22611 3943 22614
rect 4889 22611 4955 22614
rect 3509 22538 3575 22541
rect 1396 22536 3575 22538
rect 1396 22480 3514 22536
rect 3570 22480 3575 22536
rect 1396 22478 3575 22480
rect 0 22266 800 22296
rect 1396 22266 1456 22478
rect 3509 22475 3575 22478
rect 10133 22538 10199 22541
rect 11200 22538 12000 22568
rect 10133 22536 12000 22538
rect 10133 22480 10138 22536
rect 10194 22480 12000 22536
rect 10133 22478 12000 22480
rect 10133 22475 10199 22478
rect 11200 22448 12000 22478
rect 2576 22336 2896 22337
rect 2576 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2576 22271 2896 22272
rect 5840 22336 6160 22337
rect 5840 22272 5848 22336
rect 5912 22272 5928 22336
rect 5992 22272 6008 22336
rect 6072 22272 6088 22336
rect 6152 22272 6160 22336
rect 5840 22271 6160 22272
rect 9104 22336 9424 22337
rect 9104 22272 9112 22336
rect 9176 22272 9192 22336
rect 9256 22272 9272 22336
rect 9336 22272 9352 22336
rect 9416 22272 9424 22336
rect 9104 22271 9424 22272
rect 0 22206 1456 22266
rect 0 22176 800 22206
rect 0 21858 800 21888
rect 1393 21858 1459 21861
rect 0 21856 1459 21858
rect 0 21800 1398 21856
rect 1454 21800 1459 21856
rect 0 21798 1459 21800
rect 0 21768 800 21798
rect 1393 21795 1459 21798
rect 10133 21858 10199 21861
rect 11200 21858 12000 21888
rect 10133 21856 12000 21858
rect 10133 21800 10138 21856
rect 10194 21800 12000 21856
rect 10133 21798 12000 21800
rect 10133 21795 10199 21798
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 7472 21792 7792 21793
rect 7472 21728 7480 21792
rect 7544 21728 7560 21792
rect 7624 21728 7640 21792
rect 7704 21728 7720 21792
rect 7784 21728 7792 21792
rect 11200 21768 12000 21798
rect 7472 21727 7792 21728
rect 0 21450 800 21480
rect 1209 21450 1275 21453
rect 0 21448 1275 21450
rect 0 21392 1214 21448
rect 1270 21392 1275 21448
rect 0 21390 1275 21392
rect 0 21360 800 21390
rect 1209 21387 1275 21390
rect 2576 21248 2896 21249
rect 2576 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2576 21183 2896 21184
rect 5840 21248 6160 21249
rect 5840 21184 5848 21248
rect 5912 21184 5928 21248
rect 5992 21184 6008 21248
rect 6072 21184 6088 21248
rect 6152 21184 6160 21248
rect 5840 21183 6160 21184
rect 9104 21248 9424 21249
rect 9104 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9272 21248
rect 9336 21184 9352 21248
rect 9416 21184 9424 21248
rect 9104 21183 9424 21184
rect 0 21042 800 21072
rect 1393 21042 1459 21045
rect 0 21040 1459 21042
rect 0 20984 1398 21040
rect 1454 20984 1459 21040
rect 0 20982 1459 20984
rect 0 20952 800 20982
rect 1393 20979 1459 20982
rect 10133 21042 10199 21045
rect 11200 21042 12000 21072
rect 10133 21040 12000 21042
rect 10133 20984 10138 21040
rect 10194 20984 12000 21040
rect 10133 20982 12000 20984
rect 10133 20979 10199 20982
rect 11200 20952 12000 20982
rect 4208 20704 4528 20705
rect 0 20634 800 20664
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 7472 20704 7792 20705
rect 7472 20640 7480 20704
rect 7544 20640 7560 20704
rect 7624 20640 7640 20704
rect 7704 20640 7720 20704
rect 7784 20640 7792 20704
rect 7472 20639 7792 20640
rect 2773 20634 2839 20637
rect 0 20632 2839 20634
rect 0 20576 2778 20632
rect 2834 20576 2839 20632
rect 0 20574 2839 20576
rect 0 20544 800 20574
rect 2773 20571 2839 20574
rect 10041 20362 10107 20365
rect 11200 20362 12000 20392
rect 10041 20360 12000 20362
rect 10041 20304 10046 20360
rect 10102 20304 12000 20360
rect 10041 20302 12000 20304
rect 10041 20299 10107 20302
rect 11200 20272 12000 20302
rect 0 20226 800 20256
rect 1393 20226 1459 20229
rect 0 20224 1459 20226
rect 0 20168 1398 20224
rect 1454 20168 1459 20224
rect 0 20166 1459 20168
rect 0 20136 800 20166
rect 1393 20163 1459 20166
rect 2576 20160 2896 20161
rect 2576 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2576 20095 2896 20096
rect 5840 20160 6160 20161
rect 5840 20096 5848 20160
rect 5912 20096 5928 20160
rect 5992 20096 6008 20160
rect 6072 20096 6088 20160
rect 6152 20096 6160 20160
rect 5840 20095 6160 20096
rect 9104 20160 9424 20161
rect 9104 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9272 20160
rect 9336 20096 9352 20160
rect 9416 20096 9424 20160
rect 9104 20095 9424 20096
rect 0 19682 800 19712
rect 1393 19682 1459 19685
rect 0 19680 1459 19682
rect 0 19624 1398 19680
rect 1454 19624 1459 19680
rect 0 19622 1459 19624
rect 0 19592 800 19622
rect 1393 19619 1459 19622
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 7472 19616 7792 19617
rect 7472 19552 7480 19616
rect 7544 19552 7560 19616
rect 7624 19552 7640 19616
rect 7704 19552 7720 19616
rect 7784 19552 7792 19616
rect 7472 19551 7792 19552
rect 10041 19546 10107 19549
rect 11200 19546 12000 19576
rect 10041 19544 12000 19546
rect 10041 19488 10046 19544
rect 10102 19488 12000 19544
rect 10041 19486 12000 19488
rect 10041 19483 10107 19486
rect 11200 19456 12000 19486
rect 0 19274 800 19304
rect 1209 19274 1275 19277
rect 0 19272 1275 19274
rect 0 19216 1214 19272
rect 1270 19216 1275 19272
rect 0 19214 1275 19216
rect 0 19184 800 19214
rect 1209 19211 1275 19214
rect 2576 19072 2896 19073
rect 2576 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2576 19007 2896 19008
rect 5840 19072 6160 19073
rect 5840 19008 5848 19072
rect 5912 19008 5928 19072
rect 5992 19008 6008 19072
rect 6072 19008 6088 19072
rect 6152 19008 6160 19072
rect 5840 19007 6160 19008
rect 9104 19072 9424 19073
rect 9104 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9272 19072
rect 9336 19008 9352 19072
rect 9416 19008 9424 19072
rect 9104 19007 9424 19008
rect 0 18866 800 18896
rect 1393 18866 1459 18869
rect 0 18864 1459 18866
rect 0 18808 1398 18864
rect 1454 18808 1459 18864
rect 0 18806 1459 18808
rect 0 18776 800 18806
rect 1393 18803 1459 18806
rect 10041 18730 10107 18733
rect 11200 18730 12000 18760
rect 10041 18728 12000 18730
rect 10041 18672 10046 18728
rect 10102 18672 12000 18728
rect 10041 18670 12000 18672
rect 10041 18667 10107 18670
rect 11200 18640 12000 18670
rect 4208 18528 4528 18529
rect 0 18458 800 18488
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 7472 18528 7792 18529
rect 7472 18464 7480 18528
rect 7544 18464 7560 18528
rect 7624 18464 7640 18528
rect 7704 18464 7720 18528
rect 7784 18464 7792 18528
rect 7472 18463 7792 18464
rect 3969 18458 4035 18461
rect 0 18456 4035 18458
rect 0 18400 3974 18456
rect 4030 18400 4035 18456
rect 0 18398 4035 18400
rect 0 18368 800 18398
rect 3969 18395 4035 18398
rect 3693 18186 3759 18189
rect 1350 18184 3759 18186
rect 1350 18128 3698 18184
rect 3754 18128 3759 18184
rect 1350 18126 3759 18128
rect 0 18050 800 18080
rect 1350 18050 1410 18126
rect 3693 18123 3759 18126
rect 0 17990 1410 18050
rect 10041 18050 10107 18053
rect 11200 18050 12000 18080
rect 10041 18048 12000 18050
rect 10041 17992 10046 18048
rect 10102 17992 12000 18048
rect 10041 17990 12000 17992
rect 0 17960 800 17990
rect 10041 17987 10107 17990
rect 2576 17984 2896 17985
rect 2576 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2576 17919 2896 17920
rect 5840 17984 6160 17985
rect 5840 17920 5848 17984
rect 5912 17920 5928 17984
rect 5992 17920 6008 17984
rect 6072 17920 6088 17984
rect 6152 17920 6160 17984
rect 5840 17919 6160 17920
rect 9104 17984 9424 17985
rect 9104 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9272 17984
rect 9336 17920 9352 17984
rect 9416 17920 9424 17984
rect 11200 17960 12000 17990
rect 9104 17919 9424 17920
rect 0 17642 800 17672
rect 3049 17642 3115 17645
rect 0 17640 3115 17642
rect 0 17584 3054 17640
rect 3110 17584 3115 17640
rect 0 17582 3115 17584
rect 0 17552 800 17582
rect 3049 17579 3115 17582
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 7472 17440 7792 17441
rect 7472 17376 7480 17440
rect 7544 17376 7560 17440
rect 7624 17376 7640 17440
rect 7704 17376 7720 17440
rect 7784 17376 7792 17440
rect 7472 17375 7792 17376
rect 0 17234 800 17264
rect 2405 17234 2471 17237
rect 0 17232 2471 17234
rect 0 17176 2410 17232
rect 2466 17176 2471 17232
rect 0 17174 2471 17176
rect 0 17144 800 17174
rect 2405 17171 2471 17174
rect 10041 17234 10107 17237
rect 11200 17234 12000 17264
rect 10041 17232 12000 17234
rect 10041 17176 10046 17232
rect 10102 17176 12000 17232
rect 10041 17174 12000 17176
rect 10041 17171 10107 17174
rect 11200 17144 12000 17174
rect 2998 17036 3004 17100
rect 3068 17098 3074 17100
rect 3233 17098 3299 17101
rect 3068 17096 3299 17098
rect 3068 17040 3238 17096
rect 3294 17040 3299 17096
rect 3068 17038 3299 17040
rect 3068 17036 3074 17038
rect 3233 17035 3299 17038
rect 2576 16896 2896 16897
rect 2576 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2576 16831 2896 16832
rect 5840 16896 6160 16897
rect 5840 16832 5848 16896
rect 5912 16832 5928 16896
rect 5992 16832 6008 16896
rect 6072 16832 6088 16896
rect 6152 16832 6160 16896
rect 5840 16831 6160 16832
rect 9104 16896 9424 16897
rect 9104 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9272 16896
rect 9336 16832 9352 16896
rect 9416 16832 9424 16896
rect 9104 16831 9424 16832
rect 0 16690 800 16720
rect 1577 16690 1643 16693
rect 0 16688 1643 16690
rect 0 16632 1582 16688
rect 1638 16632 1643 16688
rect 0 16630 1643 16632
rect 0 16600 800 16630
rect 1577 16627 1643 16630
rect 10041 16418 10107 16421
rect 11200 16418 12000 16448
rect 10041 16416 12000 16418
rect 10041 16360 10046 16416
rect 10102 16360 12000 16416
rect 10041 16358 12000 16360
rect 10041 16355 10107 16358
rect 4208 16352 4528 16353
rect 0 16282 800 16312
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 7472 16352 7792 16353
rect 7472 16288 7480 16352
rect 7544 16288 7560 16352
rect 7624 16288 7640 16352
rect 7704 16288 7720 16352
rect 7784 16288 7792 16352
rect 11200 16328 12000 16358
rect 7472 16287 7792 16288
rect 3969 16282 4035 16285
rect 0 16280 4035 16282
rect 0 16224 3974 16280
rect 4030 16224 4035 16280
rect 0 16222 4035 16224
rect 0 16192 800 16222
rect 3969 16219 4035 16222
rect 2865 16010 2931 16013
rect 1350 16008 2931 16010
rect 1350 15952 2870 16008
rect 2926 15952 2931 16008
rect 1350 15950 2931 15952
rect 0 15874 800 15904
rect 1350 15874 1410 15950
rect 2865 15947 2931 15950
rect 0 15814 1410 15874
rect 0 15784 800 15814
rect 2576 15808 2896 15809
rect 2576 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2576 15743 2896 15744
rect 5840 15808 6160 15809
rect 5840 15744 5848 15808
rect 5912 15744 5928 15808
rect 5992 15744 6008 15808
rect 6072 15744 6088 15808
rect 6152 15744 6160 15808
rect 5840 15743 6160 15744
rect 9104 15808 9424 15809
rect 9104 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9272 15808
rect 9336 15744 9352 15808
rect 9416 15744 9424 15808
rect 9104 15743 9424 15744
rect 3417 15740 3483 15741
rect 3366 15738 3372 15740
rect 3326 15678 3372 15738
rect 3436 15736 3483 15740
rect 3478 15680 3483 15736
rect 3366 15676 3372 15678
rect 3436 15676 3483 15680
rect 3417 15675 3483 15676
rect 10041 15738 10107 15741
rect 11200 15738 12000 15768
rect 10041 15736 12000 15738
rect 10041 15680 10046 15736
rect 10102 15680 12000 15736
rect 10041 15678 12000 15680
rect 10041 15675 10107 15678
rect 11200 15648 12000 15678
rect 0 15466 800 15496
rect 2221 15466 2287 15469
rect 0 15464 2287 15466
rect 0 15408 2226 15464
rect 2282 15408 2287 15464
rect 0 15406 2287 15408
rect 0 15376 800 15406
rect 2221 15403 2287 15406
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 7472 15264 7792 15265
rect 7472 15200 7480 15264
rect 7544 15200 7560 15264
rect 7624 15200 7640 15264
rect 7704 15200 7720 15264
rect 7784 15200 7792 15264
rect 7472 15199 7792 15200
rect 0 15058 800 15088
rect 1209 15058 1275 15061
rect 0 15056 1275 15058
rect 0 15000 1214 15056
rect 1270 15000 1275 15056
rect 0 14998 1275 15000
rect 0 14968 800 14998
rect 1209 14995 1275 14998
rect 10041 14922 10107 14925
rect 11200 14922 12000 14952
rect 10041 14920 12000 14922
rect 10041 14864 10046 14920
rect 10102 14864 12000 14920
rect 10041 14862 12000 14864
rect 10041 14859 10107 14862
rect 11200 14832 12000 14862
rect 2576 14720 2896 14721
rect 0 14650 800 14680
rect 2576 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2576 14655 2896 14656
rect 5840 14720 6160 14721
rect 5840 14656 5848 14720
rect 5912 14656 5928 14720
rect 5992 14656 6008 14720
rect 6072 14656 6088 14720
rect 6152 14656 6160 14720
rect 5840 14655 6160 14656
rect 9104 14720 9424 14721
rect 9104 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9272 14720
rect 9336 14656 9352 14720
rect 9416 14656 9424 14720
rect 9104 14655 9424 14656
rect 1393 14650 1459 14653
rect 0 14648 1459 14650
rect 0 14592 1398 14648
rect 1454 14592 1459 14648
rect 0 14590 1459 14592
rect 0 14560 800 14590
rect 1393 14587 1459 14590
rect 0 14242 800 14272
rect 3969 14242 4035 14245
rect 0 14240 4035 14242
rect 0 14184 3974 14240
rect 4030 14184 4035 14240
rect 0 14182 4035 14184
rect 0 14152 800 14182
rect 3969 14179 4035 14182
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 7472 14176 7792 14177
rect 7472 14112 7480 14176
rect 7544 14112 7560 14176
rect 7624 14112 7640 14176
rect 7704 14112 7720 14176
rect 7784 14112 7792 14176
rect 7472 14111 7792 14112
rect 3601 14108 3667 14109
rect 3550 14106 3556 14108
rect 3510 14046 3556 14106
rect 3620 14104 3667 14108
rect 3662 14048 3667 14104
rect 3550 14044 3556 14046
rect 3620 14044 3667 14048
rect 3601 14043 3667 14044
rect 10041 14106 10107 14109
rect 11200 14106 12000 14136
rect 10041 14104 12000 14106
rect 10041 14048 10046 14104
rect 10102 14048 12000 14104
rect 10041 14046 12000 14048
rect 10041 14043 10107 14046
rect 11200 14016 12000 14046
rect 0 13834 800 13864
rect 2957 13834 3023 13837
rect 0 13832 3023 13834
rect 0 13776 2962 13832
rect 3018 13776 3023 13832
rect 0 13774 3023 13776
rect 0 13744 800 13774
rect 2957 13771 3023 13774
rect 2576 13632 2896 13633
rect 2576 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2576 13567 2896 13568
rect 5840 13632 6160 13633
rect 5840 13568 5848 13632
rect 5912 13568 5928 13632
rect 5992 13568 6008 13632
rect 6072 13568 6088 13632
rect 6152 13568 6160 13632
rect 5840 13567 6160 13568
rect 9104 13632 9424 13633
rect 9104 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9272 13632
rect 9336 13568 9352 13632
rect 9416 13568 9424 13632
rect 9104 13567 9424 13568
rect 3877 13426 3943 13429
rect 3742 13424 3943 13426
rect 3742 13368 3882 13424
rect 3938 13368 3943 13424
rect 3742 13366 3943 13368
rect 0 13290 800 13320
rect 3417 13290 3483 13293
rect 0 13288 3483 13290
rect 0 13232 3422 13288
rect 3478 13232 3483 13288
rect 0 13230 3483 13232
rect 0 13200 800 13230
rect 3417 13227 3483 13230
rect 3509 13018 3575 13021
rect 3742 13018 3802 13366
rect 3877 13363 3943 13366
rect 9581 13426 9647 13429
rect 11200 13426 12000 13456
rect 9581 13424 12000 13426
rect 9581 13368 9586 13424
rect 9642 13368 12000 13424
rect 9581 13366 12000 13368
rect 9581 13363 9647 13366
rect 11200 13336 12000 13366
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 7472 13088 7792 13089
rect 7472 13024 7480 13088
rect 7544 13024 7560 13088
rect 7624 13024 7640 13088
rect 7704 13024 7720 13088
rect 7784 13024 7792 13088
rect 7472 13023 7792 13024
rect 3509 13016 3802 13018
rect 3509 12960 3514 13016
rect 3570 12960 3802 13016
rect 3509 12958 3802 12960
rect 3509 12955 3575 12958
rect 0 12882 800 12912
rect 3969 12882 4035 12885
rect 0 12880 4035 12882
rect 0 12824 3974 12880
rect 4030 12824 4035 12880
rect 0 12822 4035 12824
rect 0 12792 800 12822
rect 3969 12819 4035 12822
rect 10041 12610 10107 12613
rect 11200 12610 12000 12640
rect 10041 12608 12000 12610
rect 10041 12552 10046 12608
rect 10102 12552 12000 12608
rect 10041 12550 12000 12552
rect 10041 12547 10107 12550
rect 2576 12544 2896 12545
rect 0 12474 800 12504
rect 2576 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2576 12479 2896 12480
rect 5840 12544 6160 12545
rect 5840 12480 5848 12544
rect 5912 12480 5928 12544
rect 5992 12480 6008 12544
rect 6072 12480 6088 12544
rect 6152 12480 6160 12544
rect 5840 12479 6160 12480
rect 9104 12544 9424 12545
rect 9104 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9272 12544
rect 9336 12480 9352 12544
rect 9416 12480 9424 12544
rect 11200 12520 12000 12550
rect 9104 12479 9424 12480
rect 1485 12474 1551 12477
rect 0 12472 1551 12474
rect 0 12416 1490 12472
rect 1546 12416 1551 12472
rect 0 12414 1551 12416
rect 0 12384 800 12414
rect 1485 12411 1551 12414
rect 3417 12474 3483 12477
rect 3550 12474 3556 12476
rect 3417 12472 3556 12474
rect 3417 12416 3422 12472
rect 3478 12416 3556 12472
rect 3417 12414 3556 12416
rect 3417 12411 3483 12414
rect 3550 12412 3556 12414
rect 3620 12412 3626 12476
rect 0 12066 800 12096
rect 1577 12066 1643 12069
rect 0 12064 1643 12066
rect 0 12008 1582 12064
rect 1638 12008 1643 12064
rect 0 12006 1643 12008
rect 0 11976 800 12006
rect 1577 12003 1643 12006
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 7472 12000 7792 12001
rect 7472 11936 7480 12000
rect 7544 11936 7560 12000
rect 7624 11936 7640 12000
rect 7704 11936 7720 12000
rect 7784 11936 7792 12000
rect 7472 11935 7792 11936
rect 3049 11796 3115 11797
rect 2998 11794 3004 11796
rect 2958 11734 3004 11794
rect 3068 11792 3115 11796
rect 3110 11736 3115 11792
rect 2998 11732 3004 11734
rect 3068 11732 3115 11736
rect 3049 11731 3115 11732
rect 10041 11794 10107 11797
rect 11200 11794 12000 11824
rect 10041 11792 12000 11794
rect 10041 11736 10046 11792
rect 10102 11736 12000 11792
rect 10041 11734 12000 11736
rect 10041 11731 10107 11734
rect 11200 11704 12000 11734
rect 0 11658 800 11688
rect 3693 11658 3759 11661
rect 0 11656 3759 11658
rect 0 11600 3698 11656
rect 3754 11600 3759 11656
rect 0 11598 3759 11600
rect 0 11568 800 11598
rect 3693 11595 3759 11598
rect 2957 11522 3023 11525
rect 3366 11522 3372 11524
rect 2957 11520 3372 11522
rect 2957 11464 2962 11520
rect 3018 11464 3372 11520
rect 2957 11462 3372 11464
rect 2957 11459 3023 11462
rect 3366 11460 3372 11462
rect 3436 11460 3442 11524
rect 2576 11456 2896 11457
rect 2576 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2576 11391 2896 11392
rect 5840 11456 6160 11457
rect 5840 11392 5848 11456
rect 5912 11392 5928 11456
rect 5992 11392 6008 11456
rect 6072 11392 6088 11456
rect 6152 11392 6160 11456
rect 5840 11391 6160 11392
rect 9104 11456 9424 11457
rect 9104 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9272 11456
rect 9336 11392 9352 11456
rect 9416 11392 9424 11456
rect 9104 11391 9424 11392
rect 0 11250 800 11280
rect 1209 11250 1275 11253
rect 0 11248 1275 11250
rect 0 11192 1214 11248
rect 1270 11192 1275 11248
rect 0 11190 1275 11192
rect 0 11160 800 11190
rect 1209 11187 1275 11190
rect 10041 11114 10107 11117
rect 11200 11114 12000 11144
rect 10041 11112 12000 11114
rect 10041 11056 10046 11112
rect 10102 11056 12000 11112
rect 10041 11054 12000 11056
rect 10041 11051 10107 11054
rect 11200 11024 12000 11054
rect 4208 10912 4528 10913
rect 0 10842 800 10872
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 7472 10912 7792 10913
rect 7472 10848 7480 10912
rect 7544 10848 7560 10912
rect 7624 10848 7640 10912
rect 7704 10848 7720 10912
rect 7784 10848 7792 10912
rect 7472 10847 7792 10848
rect 1393 10842 1459 10845
rect 0 10840 1459 10842
rect 0 10784 1398 10840
rect 1454 10784 1459 10840
rect 0 10782 1459 10784
rect 0 10752 800 10782
rect 1393 10779 1459 10782
rect 0 10434 800 10464
rect 1485 10434 1551 10437
rect 0 10432 1551 10434
rect 0 10376 1490 10432
rect 1546 10376 1551 10432
rect 0 10374 1551 10376
rect 0 10344 800 10374
rect 1485 10371 1551 10374
rect 2576 10368 2896 10369
rect 2576 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2576 10303 2896 10304
rect 5840 10368 6160 10369
rect 5840 10304 5848 10368
rect 5912 10304 5928 10368
rect 5992 10304 6008 10368
rect 6072 10304 6088 10368
rect 6152 10304 6160 10368
rect 5840 10303 6160 10304
rect 9104 10368 9424 10369
rect 9104 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9272 10368
rect 9336 10304 9352 10368
rect 9416 10304 9424 10368
rect 9104 10303 9424 10304
rect 3969 10300 4035 10301
rect 3918 10236 3924 10300
rect 3988 10298 4035 10300
rect 10041 10298 10107 10301
rect 11200 10298 12000 10328
rect 3988 10296 4080 10298
rect 4030 10240 4080 10296
rect 3988 10238 4080 10240
rect 10041 10296 12000 10298
rect 10041 10240 10046 10296
rect 10102 10240 12000 10296
rect 10041 10238 12000 10240
rect 3988 10236 4035 10238
rect 3969 10235 4035 10236
rect 10041 10235 10107 10238
rect 11200 10208 12000 10238
rect 0 9890 800 9920
rect 1393 9890 1459 9893
rect 0 9888 1459 9890
rect 0 9832 1398 9888
rect 1454 9832 1459 9888
rect 0 9830 1459 9832
rect 0 9800 800 9830
rect 1393 9827 1459 9830
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 7472 9824 7792 9825
rect 7472 9760 7480 9824
rect 7544 9760 7560 9824
rect 7624 9760 7640 9824
rect 7704 9760 7720 9824
rect 7784 9760 7792 9824
rect 7472 9759 7792 9760
rect 0 9482 800 9512
rect 1485 9482 1551 9485
rect 0 9480 1551 9482
rect 0 9424 1490 9480
rect 1546 9424 1551 9480
rect 0 9422 1551 9424
rect 0 9392 800 9422
rect 1485 9419 1551 9422
rect 10041 9482 10107 9485
rect 11200 9482 12000 9512
rect 10041 9480 12000 9482
rect 10041 9424 10046 9480
rect 10102 9424 12000 9480
rect 10041 9422 12000 9424
rect 10041 9419 10107 9422
rect 11200 9392 12000 9422
rect 2576 9280 2896 9281
rect 2576 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2576 9215 2896 9216
rect 5840 9280 6160 9281
rect 5840 9216 5848 9280
rect 5912 9216 5928 9280
rect 5992 9216 6008 9280
rect 6072 9216 6088 9280
rect 6152 9216 6160 9280
rect 5840 9215 6160 9216
rect 9104 9280 9424 9281
rect 9104 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9272 9280
rect 9336 9216 9352 9280
rect 9416 9216 9424 9280
rect 9104 9215 9424 9216
rect 0 9074 800 9104
rect 1393 9074 1459 9077
rect 0 9072 1459 9074
rect 0 9016 1398 9072
rect 1454 9016 1459 9072
rect 0 9014 1459 9016
rect 0 8984 800 9014
rect 1393 9011 1459 9014
rect 10041 8802 10107 8805
rect 11200 8802 12000 8832
rect 10041 8800 12000 8802
rect 10041 8744 10046 8800
rect 10102 8744 12000 8800
rect 10041 8742 12000 8744
rect 10041 8739 10107 8742
rect 4208 8736 4528 8737
rect 0 8666 800 8696
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 7472 8736 7792 8737
rect 7472 8672 7480 8736
rect 7544 8672 7560 8736
rect 7624 8672 7640 8736
rect 7704 8672 7720 8736
rect 7784 8672 7792 8736
rect 11200 8712 12000 8742
rect 7472 8671 7792 8672
rect 1393 8666 1459 8669
rect 0 8664 1459 8666
rect 0 8608 1398 8664
rect 1454 8608 1459 8664
rect 0 8606 1459 8608
rect 0 8576 800 8606
rect 1393 8603 1459 8606
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 2576 8192 2896 8193
rect 2576 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2576 8127 2896 8128
rect 5840 8192 6160 8193
rect 5840 8128 5848 8192
rect 5912 8128 5928 8192
rect 5992 8128 6008 8192
rect 6072 8128 6088 8192
rect 6152 8128 6160 8192
rect 5840 8127 6160 8128
rect 9104 8192 9424 8193
rect 9104 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9272 8192
rect 9336 8128 9352 8192
rect 9416 8128 9424 8192
rect 9104 8127 9424 8128
rect 10041 7986 10107 7989
rect 11200 7986 12000 8016
rect 10041 7984 12000 7986
rect 10041 7928 10046 7984
rect 10102 7928 12000 7984
rect 10041 7926 12000 7928
rect 10041 7923 10107 7926
rect 11200 7896 12000 7926
rect 0 7850 800 7880
rect 1393 7850 1459 7853
rect 0 7848 1459 7850
rect 0 7792 1398 7848
rect 1454 7792 1459 7848
rect 0 7790 1459 7792
rect 0 7760 800 7790
rect 1393 7787 1459 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 7472 7648 7792 7649
rect 7472 7584 7480 7648
rect 7544 7584 7560 7648
rect 7624 7584 7640 7648
rect 7704 7584 7720 7648
rect 7784 7584 7792 7648
rect 7472 7583 7792 7584
rect 0 7442 800 7472
rect 2957 7442 3023 7445
rect 0 7440 3023 7442
rect 0 7384 2962 7440
rect 3018 7384 3023 7440
rect 0 7382 3023 7384
rect 0 7352 800 7382
rect 2957 7379 3023 7382
rect 3601 7306 3667 7309
rect 1902 7304 3667 7306
rect 1902 7248 3606 7304
rect 3662 7248 3667 7304
rect 1902 7246 3667 7248
rect 0 7034 800 7064
rect 1902 7034 1962 7246
rect 3601 7243 3667 7246
rect 10041 7170 10107 7173
rect 11200 7170 12000 7200
rect 10041 7168 12000 7170
rect 10041 7112 10046 7168
rect 10102 7112 12000 7168
rect 10041 7110 12000 7112
rect 10041 7107 10107 7110
rect 2576 7104 2896 7105
rect 2576 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2576 7039 2896 7040
rect 5840 7104 6160 7105
rect 5840 7040 5848 7104
rect 5912 7040 5928 7104
rect 5992 7040 6008 7104
rect 6072 7040 6088 7104
rect 6152 7040 6160 7104
rect 5840 7039 6160 7040
rect 9104 7104 9424 7105
rect 9104 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9272 7104
rect 9336 7040 9352 7104
rect 9416 7040 9424 7104
rect 11200 7080 12000 7110
rect 9104 7039 9424 7040
rect 0 6974 1962 7034
rect 0 6944 800 6974
rect 2589 6762 2655 6765
rect 5022 6762 5028 6764
rect 2589 6760 5028 6762
rect 2589 6704 2594 6760
rect 2650 6704 5028 6760
rect 2589 6702 5028 6704
rect 2589 6699 2655 6702
rect 5022 6700 5028 6702
rect 5092 6700 5098 6764
rect 4208 6560 4528 6561
rect 0 6490 800 6520
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 7472 6560 7792 6561
rect 7472 6496 7480 6560
rect 7544 6496 7560 6560
rect 7624 6496 7640 6560
rect 7704 6496 7720 6560
rect 7784 6496 7792 6560
rect 7472 6495 7792 6496
rect 3141 6490 3207 6493
rect 0 6488 3207 6490
rect 0 6432 3146 6488
rect 3202 6432 3207 6488
rect 0 6430 3207 6432
rect 0 6400 800 6430
rect 3141 6427 3207 6430
rect 10041 6490 10107 6493
rect 11200 6490 12000 6520
rect 10041 6488 12000 6490
rect 10041 6432 10046 6488
rect 10102 6432 12000 6488
rect 10041 6430 12000 6432
rect 10041 6427 10107 6430
rect 11200 6400 12000 6430
rect 2957 6218 3023 6221
rect 1534 6216 3023 6218
rect 1534 6160 2962 6216
rect 3018 6160 3023 6216
rect 1534 6158 3023 6160
rect 0 6082 800 6112
rect 1534 6082 1594 6158
rect 2957 6155 3023 6158
rect 0 6022 1594 6082
rect 0 5992 800 6022
rect 2576 6016 2896 6017
rect 2576 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2576 5951 2896 5952
rect 5840 6016 6160 6017
rect 5840 5952 5848 6016
rect 5912 5952 5928 6016
rect 5992 5952 6008 6016
rect 6072 5952 6088 6016
rect 6152 5952 6160 6016
rect 5840 5951 6160 5952
rect 9104 6016 9424 6017
rect 9104 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9272 6016
rect 9336 5952 9352 6016
rect 9416 5952 9424 6016
rect 9104 5951 9424 5952
rect 2957 5946 3023 5949
rect 4654 5946 4660 5948
rect 2957 5944 4660 5946
rect 2957 5888 2962 5944
rect 3018 5888 4660 5944
rect 2957 5886 4660 5888
rect 2957 5883 3023 5886
rect 4654 5884 4660 5886
rect 4724 5884 4730 5948
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 10041 5674 10107 5677
rect 11200 5674 12000 5704
rect 10041 5672 12000 5674
rect 10041 5616 10046 5672
rect 10102 5616 12000 5672
rect 10041 5614 12000 5616
rect 10041 5611 10107 5614
rect 11200 5584 12000 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 7472 5472 7792 5473
rect 7472 5408 7480 5472
rect 7544 5408 7560 5472
rect 7624 5408 7640 5472
rect 7704 5408 7720 5472
rect 7784 5408 7792 5472
rect 7472 5407 7792 5408
rect 0 5266 800 5296
rect 1393 5266 1459 5269
rect 0 5264 1459 5266
rect 0 5208 1398 5264
rect 1454 5208 1459 5264
rect 0 5206 1459 5208
rect 0 5176 800 5206
rect 1393 5203 1459 5206
rect 2865 5266 2931 5269
rect 4838 5266 4844 5268
rect 2865 5264 4844 5266
rect 2865 5208 2870 5264
rect 2926 5208 4844 5264
rect 2865 5206 4844 5208
rect 2865 5203 2931 5206
rect 4838 5204 4844 5206
rect 4908 5204 4914 5268
rect 2576 4928 2896 4929
rect 0 4858 800 4888
rect 2576 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2576 4863 2896 4864
rect 5840 4928 6160 4929
rect 5840 4864 5848 4928
rect 5912 4864 5928 4928
rect 5992 4864 6008 4928
rect 6072 4864 6088 4928
rect 6152 4864 6160 4928
rect 5840 4863 6160 4864
rect 9104 4928 9424 4929
rect 9104 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9272 4928
rect 9336 4864 9352 4928
rect 9416 4864 9424 4928
rect 9104 4863 9424 4864
rect 10041 4858 10107 4861
rect 11200 4858 12000 4888
rect 0 4798 2330 4858
rect 0 4768 800 4798
rect 2270 4722 2330 4798
rect 10041 4856 12000 4858
rect 10041 4800 10046 4856
rect 10102 4800 12000 4856
rect 10041 4798 12000 4800
rect 10041 4795 10107 4798
rect 11200 4768 12000 4798
rect 4061 4722 4127 4725
rect 2270 4720 4127 4722
rect 2270 4664 4066 4720
rect 4122 4664 4127 4720
rect 2270 4662 4127 4664
rect 4061 4659 4127 4662
rect 0 4450 800 4480
rect 3601 4450 3667 4453
rect 0 4448 3667 4450
rect 0 4392 3606 4448
rect 3662 4392 3667 4448
rect 0 4390 3667 4392
rect 0 4360 800 4390
rect 3601 4387 3667 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 7472 4384 7792 4385
rect 7472 4320 7480 4384
rect 7544 4320 7560 4384
rect 7624 4320 7640 4384
rect 7704 4320 7720 4384
rect 7784 4320 7792 4384
rect 7472 4319 7792 4320
rect 10041 4178 10107 4181
rect 11200 4178 12000 4208
rect 10041 4176 12000 4178
rect 10041 4120 10046 4176
rect 10102 4120 12000 4176
rect 10041 4118 12000 4120
rect 10041 4115 10107 4118
rect 11200 4088 12000 4118
rect 0 4042 800 4072
rect 1485 4042 1551 4045
rect 0 4040 1551 4042
rect 0 3984 1490 4040
rect 1546 3984 1551 4040
rect 0 3982 1551 3984
rect 0 3952 800 3982
rect 1485 3979 1551 3982
rect 2576 3840 2896 3841
rect 2576 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2576 3775 2896 3776
rect 5840 3840 6160 3841
rect 5840 3776 5848 3840
rect 5912 3776 5928 3840
rect 5992 3776 6008 3840
rect 6072 3776 6088 3840
rect 6152 3776 6160 3840
rect 5840 3775 6160 3776
rect 9104 3840 9424 3841
rect 9104 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9272 3840
rect 9336 3776 9352 3840
rect 9416 3776 9424 3840
rect 9104 3775 9424 3776
rect 0 3634 800 3664
rect 1393 3634 1459 3637
rect 0 3632 1459 3634
rect 0 3576 1398 3632
rect 1454 3576 1459 3632
rect 0 3574 1459 3576
rect 0 3544 800 3574
rect 1393 3571 1459 3574
rect 10041 3362 10107 3365
rect 11200 3362 12000 3392
rect 10041 3360 12000 3362
rect 10041 3304 10046 3360
rect 10102 3304 12000 3360
rect 10041 3302 12000 3304
rect 10041 3299 10107 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 7472 3296 7792 3297
rect 7472 3232 7480 3296
rect 7544 3232 7560 3296
rect 7624 3232 7640 3296
rect 7704 3232 7720 3296
rect 7784 3232 7792 3296
rect 11200 3272 12000 3302
rect 7472 3231 7792 3232
rect 0 3090 800 3120
rect 1577 3090 1643 3093
rect 0 3088 1643 3090
rect 0 3032 1582 3088
rect 1638 3032 1643 3088
rect 0 3030 1643 3032
rect 0 3000 800 3030
rect 1577 3027 1643 3030
rect 2576 2752 2896 2753
rect 0 2682 800 2712
rect 2576 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2576 2687 2896 2688
rect 5840 2752 6160 2753
rect 5840 2688 5848 2752
rect 5912 2688 5928 2752
rect 5992 2688 6008 2752
rect 6072 2688 6088 2752
rect 6152 2688 6160 2752
rect 5840 2687 6160 2688
rect 9104 2752 9424 2753
rect 9104 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9272 2752
rect 9336 2688 9352 2752
rect 9416 2688 9424 2752
rect 9104 2687 9424 2688
rect 0 2622 1778 2682
rect 0 2592 800 2622
rect 1718 2546 1778 2622
rect 3509 2546 3575 2549
rect 1718 2544 3575 2546
rect 1718 2488 3514 2544
rect 3570 2488 3575 2544
rect 1718 2486 3575 2488
rect 3509 2483 3575 2486
rect 10041 2546 10107 2549
rect 11200 2546 12000 2576
rect 10041 2544 12000 2546
rect 10041 2488 10046 2544
rect 10102 2488 12000 2544
rect 10041 2486 12000 2488
rect 10041 2483 10107 2486
rect 11200 2456 12000 2486
rect 0 2274 800 2304
rect 2957 2274 3023 2277
rect 0 2272 3023 2274
rect 0 2216 2962 2272
rect 3018 2216 3023 2272
rect 0 2214 3023 2216
rect 0 2184 800 2214
rect 2957 2211 3023 2214
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 7472 2208 7792 2209
rect 7472 2144 7480 2208
rect 7544 2144 7560 2208
rect 7624 2144 7640 2208
rect 7704 2144 7720 2208
rect 7784 2144 7792 2208
rect 7472 2143 7792 2144
rect 0 1866 800 1896
rect 2221 1866 2287 1869
rect 0 1864 2287 1866
rect 0 1808 2226 1864
rect 2282 1808 2287 1864
rect 0 1806 2287 1808
rect 0 1776 800 1806
rect 2221 1803 2287 1806
rect 9489 1866 9555 1869
rect 11200 1866 12000 1896
rect 9489 1864 12000 1866
rect 9489 1808 9494 1864
rect 9550 1808 12000 1864
rect 9489 1806 12000 1808
rect 9489 1803 9555 1806
rect 11200 1776 12000 1806
rect 0 1458 800 1488
rect 2865 1458 2931 1461
rect 0 1456 2931 1458
rect 0 1400 2870 1456
rect 2926 1400 2931 1456
rect 0 1398 2931 1400
rect 0 1368 800 1398
rect 2865 1395 2931 1398
rect 0 1050 800 1080
rect 2865 1050 2931 1053
rect 0 1048 2931 1050
rect 0 992 2870 1048
rect 2926 992 2931 1048
rect 0 990 2931 992
rect 0 960 800 990
rect 2865 987 2931 990
rect 9581 1050 9647 1053
rect 11200 1050 12000 1080
rect 9581 1048 12000 1050
rect 9581 992 9586 1048
rect 9642 992 12000 1048
rect 9581 990 12000 992
rect 9581 987 9647 990
rect 11200 960 12000 990
rect 0 642 800 672
rect 2773 642 2839 645
rect 0 640 2839 642
rect 0 584 2778 640
rect 2834 584 2839 640
rect 0 582 2839 584
rect 0 552 800 582
rect 2773 579 2839 582
rect 9305 370 9371 373
rect 11200 370 12000 400
rect 9305 368 12000 370
rect 9305 312 9310 368
rect 9366 312 12000 368
rect 9305 310 12000 312
rect 9305 307 9371 310
rect 11200 280 12000 310
rect 0 234 800 264
rect 3969 234 4035 237
rect 0 232 4035 234
rect 0 176 3974 232
rect 4030 176 4035 232
rect 0 174 4035 176
rect 0 144 800 174
rect 3969 171 4035 174
<< via3 >>
rect 2584 77820 2648 77824
rect 2584 77764 2588 77820
rect 2588 77764 2644 77820
rect 2644 77764 2648 77820
rect 2584 77760 2648 77764
rect 2664 77820 2728 77824
rect 2664 77764 2668 77820
rect 2668 77764 2724 77820
rect 2724 77764 2728 77820
rect 2664 77760 2728 77764
rect 2744 77820 2808 77824
rect 2744 77764 2748 77820
rect 2748 77764 2804 77820
rect 2804 77764 2808 77820
rect 2744 77760 2808 77764
rect 2824 77820 2888 77824
rect 2824 77764 2828 77820
rect 2828 77764 2884 77820
rect 2884 77764 2888 77820
rect 2824 77760 2888 77764
rect 5848 77820 5912 77824
rect 5848 77764 5852 77820
rect 5852 77764 5908 77820
rect 5908 77764 5912 77820
rect 5848 77760 5912 77764
rect 5928 77820 5992 77824
rect 5928 77764 5932 77820
rect 5932 77764 5988 77820
rect 5988 77764 5992 77820
rect 5928 77760 5992 77764
rect 6008 77820 6072 77824
rect 6008 77764 6012 77820
rect 6012 77764 6068 77820
rect 6068 77764 6072 77820
rect 6008 77760 6072 77764
rect 6088 77820 6152 77824
rect 6088 77764 6092 77820
rect 6092 77764 6148 77820
rect 6148 77764 6152 77820
rect 6088 77760 6152 77764
rect 9112 77820 9176 77824
rect 9112 77764 9116 77820
rect 9116 77764 9172 77820
rect 9172 77764 9176 77820
rect 9112 77760 9176 77764
rect 9192 77820 9256 77824
rect 9192 77764 9196 77820
rect 9196 77764 9252 77820
rect 9252 77764 9256 77820
rect 9192 77760 9256 77764
rect 9272 77820 9336 77824
rect 9272 77764 9276 77820
rect 9276 77764 9332 77820
rect 9332 77764 9336 77820
rect 9272 77760 9336 77764
rect 9352 77820 9416 77824
rect 9352 77764 9356 77820
rect 9356 77764 9412 77820
rect 9412 77764 9416 77820
rect 9352 77760 9416 77764
rect 4216 77276 4280 77280
rect 4216 77220 4220 77276
rect 4220 77220 4276 77276
rect 4276 77220 4280 77276
rect 4216 77216 4280 77220
rect 4296 77276 4360 77280
rect 4296 77220 4300 77276
rect 4300 77220 4356 77276
rect 4356 77220 4360 77276
rect 4296 77216 4360 77220
rect 4376 77276 4440 77280
rect 4376 77220 4380 77276
rect 4380 77220 4436 77276
rect 4436 77220 4440 77276
rect 4376 77216 4440 77220
rect 4456 77276 4520 77280
rect 4456 77220 4460 77276
rect 4460 77220 4516 77276
rect 4516 77220 4520 77276
rect 4456 77216 4520 77220
rect 7480 77276 7544 77280
rect 7480 77220 7484 77276
rect 7484 77220 7540 77276
rect 7540 77220 7544 77276
rect 7480 77216 7544 77220
rect 7560 77276 7624 77280
rect 7560 77220 7564 77276
rect 7564 77220 7620 77276
rect 7620 77220 7624 77276
rect 7560 77216 7624 77220
rect 7640 77276 7704 77280
rect 7640 77220 7644 77276
rect 7644 77220 7700 77276
rect 7700 77220 7704 77276
rect 7640 77216 7704 77220
rect 7720 77276 7784 77280
rect 7720 77220 7724 77276
rect 7724 77220 7780 77276
rect 7780 77220 7784 77276
rect 7720 77216 7784 77220
rect 2584 76732 2648 76736
rect 2584 76676 2588 76732
rect 2588 76676 2644 76732
rect 2644 76676 2648 76732
rect 2584 76672 2648 76676
rect 2664 76732 2728 76736
rect 2664 76676 2668 76732
rect 2668 76676 2724 76732
rect 2724 76676 2728 76732
rect 2664 76672 2728 76676
rect 2744 76732 2808 76736
rect 2744 76676 2748 76732
rect 2748 76676 2804 76732
rect 2804 76676 2808 76732
rect 2744 76672 2808 76676
rect 2824 76732 2888 76736
rect 2824 76676 2828 76732
rect 2828 76676 2884 76732
rect 2884 76676 2888 76732
rect 2824 76672 2888 76676
rect 5848 76732 5912 76736
rect 5848 76676 5852 76732
rect 5852 76676 5908 76732
rect 5908 76676 5912 76732
rect 5848 76672 5912 76676
rect 5928 76732 5992 76736
rect 5928 76676 5932 76732
rect 5932 76676 5988 76732
rect 5988 76676 5992 76732
rect 5928 76672 5992 76676
rect 6008 76732 6072 76736
rect 6008 76676 6012 76732
rect 6012 76676 6068 76732
rect 6068 76676 6072 76732
rect 6008 76672 6072 76676
rect 6088 76732 6152 76736
rect 6088 76676 6092 76732
rect 6092 76676 6148 76732
rect 6148 76676 6152 76732
rect 6088 76672 6152 76676
rect 9112 76732 9176 76736
rect 9112 76676 9116 76732
rect 9116 76676 9172 76732
rect 9172 76676 9176 76732
rect 9112 76672 9176 76676
rect 9192 76732 9256 76736
rect 9192 76676 9196 76732
rect 9196 76676 9252 76732
rect 9252 76676 9256 76732
rect 9192 76672 9256 76676
rect 9272 76732 9336 76736
rect 9272 76676 9276 76732
rect 9276 76676 9332 76732
rect 9332 76676 9336 76732
rect 9272 76672 9336 76676
rect 9352 76732 9416 76736
rect 9352 76676 9356 76732
rect 9356 76676 9412 76732
rect 9412 76676 9416 76732
rect 9352 76672 9416 76676
rect 4216 76188 4280 76192
rect 4216 76132 4220 76188
rect 4220 76132 4276 76188
rect 4276 76132 4280 76188
rect 4216 76128 4280 76132
rect 4296 76188 4360 76192
rect 4296 76132 4300 76188
rect 4300 76132 4356 76188
rect 4356 76132 4360 76188
rect 4296 76128 4360 76132
rect 4376 76188 4440 76192
rect 4376 76132 4380 76188
rect 4380 76132 4436 76188
rect 4436 76132 4440 76188
rect 4376 76128 4440 76132
rect 4456 76188 4520 76192
rect 4456 76132 4460 76188
rect 4460 76132 4516 76188
rect 4516 76132 4520 76188
rect 4456 76128 4520 76132
rect 7480 76188 7544 76192
rect 7480 76132 7484 76188
rect 7484 76132 7540 76188
rect 7540 76132 7544 76188
rect 7480 76128 7544 76132
rect 7560 76188 7624 76192
rect 7560 76132 7564 76188
rect 7564 76132 7620 76188
rect 7620 76132 7624 76188
rect 7560 76128 7624 76132
rect 7640 76188 7704 76192
rect 7640 76132 7644 76188
rect 7644 76132 7700 76188
rect 7700 76132 7704 76188
rect 7640 76128 7704 76132
rect 7720 76188 7784 76192
rect 7720 76132 7724 76188
rect 7724 76132 7780 76188
rect 7780 76132 7784 76188
rect 7720 76128 7784 76132
rect 2584 75644 2648 75648
rect 2584 75588 2588 75644
rect 2588 75588 2644 75644
rect 2644 75588 2648 75644
rect 2584 75584 2648 75588
rect 2664 75644 2728 75648
rect 2664 75588 2668 75644
rect 2668 75588 2724 75644
rect 2724 75588 2728 75644
rect 2664 75584 2728 75588
rect 2744 75644 2808 75648
rect 2744 75588 2748 75644
rect 2748 75588 2804 75644
rect 2804 75588 2808 75644
rect 2744 75584 2808 75588
rect 2824 75644 2888 75648
rect 2824 75588 2828 75644
rect 2828 75588 2884 75644
rect 2884 75588 2888 75644
rect 2824 75584 2888 75588
rect 5848 75644 5912 75648
rect 5848 75588 5852 75644
rect 5852 75588 5908 75644
rect 5908 75588 5912 75644
rect 5848 75584 5912 75588
rect 5928 75644 5992 75648
rect 5928 75588 5932 75644
rect 5932 75588 5988 75644
rect 5988 75588 5992 75644
rect 5928 75584 5992 75588
rect 6008 75644 6072 75648
rect 6008 75588 6012 75644
rect 6012 75588 6068 75644
rect 6068 75588 6072 75644
rect 6008 75584 6072 75588
rect 6088 75644 6152 75648
rect 6088 75588 6092 75644
rect 6092 75588 6148 75644
rect 6148 75588 6152 75644
rect 6088 75584 6152 75588
rect 9112 75644 9176 75648
rect 9112 75588 9116 75644
rect 9116 75588 9172 75644
rect 9172 75588 9176 75644
rect 9112 75584 9176 75588
rect 9192 75644 9256 75648
rect 9192 75588 9196 75644
rect 9196 75588 9252 75644
rect 9252 75588 9256 75644
rect 9192 75584 9256 75588
rect 9272 75644 9336 75648
rect 9272 75588 9276 75644
rect 9276 75588 9332 75644
rect 9332 75588 9336 75644
rect 9272 75584 9336 75588
rect 9352 75644 9416 75648
rect 9352 75588 9356 75644
rect 9356 75588 9412 75644
rect 9412 75588 9416 75644
rect 9352 75584 9416 75588
rect 4216 75100 4280 75104
rect 4216 75044 4220 75100
rect 4220 75044 4276 75100
rect 4276 75044 4280 75100
rect 4216 75040 4280 75044
rect 4296 75100 4360 75104
rect 4296 75044 4300 75100
rect 4300 75044 4356 75100
rect 4356 75044 4360 75100
rect 4296 75040 4360 75044
rect 4376 75100 4440 75104
rect 4376 75044 4380 75100
rect 4380 75044 4436 75100
rect 4436 75044 4440 75100
rect 4376 75040 4440 75044
rect 4456 75100 4520 75104
rect 4456 75044 4460 75100
rect 4460 75044 4516 75100
rect 4516 75044 4520 75100
rect 4456 75040 4520 75044
rect 7480 75100 7544 75104
rect 7480 75044 7484 75100
rect 7484 75044 7540 75100
rect 7540 75044 7544 75100
rect 7480 75040 7544 75044
rect 7560 75100 7624 75104
rect 7560 75044 7564 75100
rect 7564 75044 7620 75100
rect 7620 75044 7624 75100
rect 7560 75040 7624 75044
rect 7640 75100 7704 75104
rect 7640 75044 7644 75100
rect 7644 75044 7700 75100
rect 7700 75044 7704 75100
rect 7640 75040 7704 75044
rect 7720 75100 7784 75104
rect 7720 75044 7724 75100
rect 7724 75044 7780 75100
rect 7780 75044 7784 75100
rect 7720 75040 7784 75044
rect 2084 74700 2148 74764
rect 2584 74556 2648 74560
rect 2584 74500 2588 74556
rect 2588 74500 2644 74556
rect 2644 74500 2648 74556
rect 2584 74496 2648 74500
rect 2664 74556 2728 74560
rect 2664 74500 2668 74556
rect 2668 74500 2724 74556
rect 2724 74500 2728 74556
rect 2664 74496 2728 74500
rect 2744 74556 2808 74560
rect 2744 74500 2748 74556
rect 2748 74500 2804 74556
rect 2804 74500 2808 74556
rect 2744 74496 2808 74500
rect 2824 74556 2888 74560
rect 2824 74500 2828 74556
rect 2828 74500 2884 74556
rect 2884 74500 2888 74556
rect 2824 74496 2888 74500
rect 5848 74556 5912 74560
rect 5848 74500 5852 74556
rect 5852 74500 5908 74556
rect 5908 74500 5912 74556
rect 5848 74496 5912 74500
rect 5928 74556 5992 74560
rect 5928 74500 5932 74556
rect 5932 74500 5988 74556
rect 5988 74500 5992 74556
rect 5928 74496 5992 74500
rect 6008 74556 6072 74560
rect 6008 74500 6012 74556
rect 6012 74500 6068 74556
rect 6068 74500 6072 74556
rect 6008 74496 6072 74500
rect 6088 74556 6152 74560
rect 6088 74500 6092 74556
rect 6092 74500 6148 74556
rect 6148 74500 6152 74556
rect 6088 74496 6152 74500
rect 9112 74556 9176 74560
rect 9112 74500 9116 74556
rect 9116 74500 9172 74556
rect 9172 74500 9176 74556
rect 9112 74496 9176 74500
rect 9192 74556 9256 74560
rect 9192 74500 9196 74556
rect 9196 74500 9252 74556
rect 9252 74500 9256 74556
rect 9192 74496 9256 74500
rect 9272 74556 9336 74560
rect 9272 74500 9276 74556
rect 9276 74500 9332 74556
rect 9332 74500 9336 74556
rect 9272 74496 9336 74500
rect 9352 74556 9416 74560
rect 9352 74500 9356 74556
rect 9356 74500 9412 74556
rect 9412 74500 9416 74556
rect 9352 74496 9416 74500
rect 4216 74012 4280 74016
rect 4216 73956 4220 74012
rect 4220 73956 4276 74012
rect 4276 73956 4280 74012
rect 4216 73952 4280 73956
rect 4296 74012 4360 74016
rect 4296 73956 4300 74012
rect 4300 73956 4356 74012
rect 4356 73956 4360 74012
rect 4296 73952 4360 73956
rect 4376 74012 4440 74016
rect 4376 73956 4380 74012
rect 4380 73956 4436 74012
rect 4436 73956 4440 74012
rect 4376 73952 4440 73956
rect 4456 74012 4520 74016
rect 4456 73956 4460 74012
rect 4460 73956 4516 74012
rect 4516 73956 4520 74012
rect 4456 73952 4520 73956
rect 7480 74012 7544 74016
rect 7480 73956 7484 74012
rect 7484 73956 7540 74012
rect 7540 73956 7544 74012
rect 7480 73952 7544 73956
rect 7560 74012 7624 74016
rect 7560 73956 7564 74012
rect 7564 73956 7620 74012
rect 7620 73956 7624 74012
rect 7560 73952 7624 73956
rect 7640 74012 7704 74016
rect 7640 73956 7644 74012
rect 7644 73956 7700 74012
rect 7700 73956 7704 74012
rect 7640 73952 7704 73956
rect 7720 74012 7784 74016
rect 7720 73956 7724 74012
rect 7724 73956 7780 74012
rect 7780 73956 7784 74012
rect 7720 73952 7784 73956
rect 2584 73468 2648 73472
rect 2584 73412 2588 73468
rect 2588 73412 2644 73468
rect 2644 73412 2648 73468
rect 2584 73408 2648 73412
rect 2664 73468 2728 73472
rect 2664 73412 2668 73468
rect 2668 73412 2724 73468
rect 2724 73412 2728 73468
rect 2664 73408 2728 73412
rect 2744 73468 2808 73472
rect 2744 73412 2748 73468
rect 2748 73412 2804 73468
rect 2804 73412 2808 73468
rect 2744 73408 2808 73412
rect 2824 73468 2888 73472
rect 2824 73412 2828 73468
rect 2828 73412 2884 73468
rect 2884 73412 2888 73468
rect 2824 73408 2888 73412
rect 5848 73468 5912 73472
rect 5848 73412 5852 73468
rect 5852 73412 5908 73468
rect 5908 73412 5912 73468
rect 5848 73408 5912 73412
rect 5928 73468 5992 73472
rect 5928 73412 5932 73468
rect 5932 73412 5988 73468
rect 5988 73412 5992 73468
rect 5928 73408 5992 73412
rect 6008 73468 6072 73472
rect 6008 73412 6012 73468
rect 6012 73412 6068 73468
rect 6068 73412 6072 73468
rect 6008 73408 6072 73412
rect 6088 73468 6152 73472
rect 6088 73412 6092 73468
rect 6092 73412 6148 73468
rect 6148 73412 6152 73468
rect 6088 73408 6152 73412
rect 9112 73468 9176 73472
rect 9112 73412 9116 73468
rect 9116 73412 9172 73468
rect 9172 73412 9176 73468
rect 9112 73408 9176 73412
rect 9192 73468 9256 73472
rect 9192 73412 9196 73468
rect 9196 73412 9252 73468
rect 9252 73412 9256 73468
rect 9192 73408 9256 73412
rect 9272 73468 9336 73472
rect 9272 73412 9276 73468
rect 9276 73412 9332 73468
rect 9332 73412 9336 73468
rect 9272 73408 9336 73412
rect 9352 73468 9416 73472
rect 9352 73412 9356 73468
rect 9356 73412 9412 73468
rect 9412 73412 9416 73468
rect 9352 73408 9416 73412
rect 4216 72924 4280 72928
rect 4216 72868 4220 72924
rect 4220 72868 4276 72924
rect 4276 72868 4280 72924
rect 4216 72864 4280 72868
rect 4296 72924 4360 72928
rect 4296 72868 4300 72924
rect 4300 72868 4356 72924
rect 4356 72868 4360 72924
rect 4296 72864 4360 72868
rect 4376 72924 4440 72928
rect 4376 72868 4380 72924
rect 4380 72868 4436 72924
rect 4436 72868 4440 72924
rect 4376 72864 4440 72868
rect 4456 72924 4520 72928
rect 4456 72868 4460 72924
rect 4460 72868 4516 72924
rect 4516 72868 4520 72924
rect 4456 72864 4520 72868
rect 7480 72924 7544 72928
rect 7480 72868 7484 72924
rect 7484 72868 7540 72924
rect 7540 72868 7544 72924
rect 7480 72864 7544 72868
rect 7560 72924 7624 72928
rect 7560 72868 7564 72924
rect 7564 72868 7620 72924
rect 7620 72868 7624 72924
rect 7560 72864 7624 72868
rect 7640 72924 7704 72928
rect 7640 72868 7644 72924
rect 7644 72868 7700 72924
rect 7700 72868 7704 72924
rect 7640 72864 7704 72868
rect 7720 72924 7784 72928
rect 7720 72868 7724 72924
rect 7724 72868 7780 72924
rect 7780 72868 7784 72924
rect 7720 72864 7784 72868
rect 1900 72660 1964 72724
rect 2584 72380 2648 72384
rect 2584 72324 2588 72380
rect 2588 72324 2644 72380
rect 2644 72324 2648 72380
rect 2584 72320 2648 72324
rect 2664 72380 2728 72384
rect 2664 72324 2668 72380
rect 2668 72324 2724 72380
rect 2724 72324 2728 72380
rect 2664 72320 2728 72324
rect 2744 72380 2808 72384
rect 2744 72324 2748 72380
rect 2748 72324 2804 72380
rect 2804 72324 2808 72380
rect 2744 72320 2808 72324
rect 2824 72380 2888 72384
rect 2824 72324 2828 72380
rect 2828 72324 2884 72380
rect 2884 72324 2888 72380
rect 2824 72320 2888 72324
rect 5848 72380 5912 72384
rect 5848 72324 5852 72380
rect 5852 72324 5908 72380
rect 5908 72324 5912 72380
rect 5848 72320 5912 72324
rect 5928 72380 5992 72384
rect 5928 72324 5932 72380
rect 5932 72324 5988 72380
rect 5988 72324 5992 72380
rect 5928 72320 5992 72324
rect 6008 72380 6072 72384
rect 6008 72324 6012 72380
rect 6012 72324 6068 72380
rect 6068 72324 6072 72380
rect 6008 72320 6072 72324
rect 6088 72380 6152 72384
rect 6088 72324 6092 72380
rect 6092 72324 6148 72380
rect 6148 72324 6152 72380
rect 6088 72320 6152 72324
rect 9112 72380 9176 72384
rect 9112 72324 9116 72380
rect 9116 72324 9172 72380
rect 9172 72324 9176 72380
rect 9112 72320 9176 72324
rect 9192 72380 9256 72384
rect 9192 72324 9196 72380
rect 9196 72324 9252 72380
rect 9252 72324 9256 72380
rect 9192 72320 9256 72324
rect 9272 72380 9336 72384
rect 9272 72324 9276 72380
rect 9276 72324 9332 72380
rect 9332 72324 9336 72380
rect 9272 72320 9336 72324
rect 9352 72380 9416 72384
rect 9352 72324 9356 72380
rect 9356 72324 9412 72380
rect 9412 72324 9416 72380
rect 9352 72320 9416 72324
rect 1532 72176 1596 72180
rect 1532 72120 1582 72176
rect 1582 72120 1596 72176
rect 1532 72116 1596 72120
rect 4216 71836 4280 71840
rect 4216 71780 4220 71836
rect 4220 71780 4276 71836
rect 4276 71780 4280 71836
rect 4216 71776 4280 71780
rect 4296 71836 4360 71840
rect 4296 71780 4300 71836
rect 4300 71780 4356 71836
rect 4356 71780 4360 71836
rect 4296 71776 4360 71780
rect 4376 71836 4440 71840
rect 4376 71780 4380 71836
rect 4380 71780 4436 71836
rect 4436 71780 4440 71836
rect 4376 71776 4440 71780
rect 4456 71836 4520 71840
rect 4456 71780 4460 71836
rect 4460 71780 4516 71836
rect 4516 71780 4520 71836
rect 4456 71776 4520 71780
rect 7480 71836 7544 71840
rect 7480 71780 7484 71836
rect 7484 71780 7540 71836
rect 7540 71780 7544 71836
rect 7480 71776 7544 71780
rect 7560 71836 7624 71840
rect 7560 71780 7564 71836
rect 7564 71780 7620 71836
rect 7620 71780 7624 71836
rect 7560 71776 7624 71780
rect 7640 71836 7704 71840
rect 7640 71780 7644 71836
rect 7644 71780 7700 71836
rect 7700 71780 7704 71836
rect 7640 71776 7704 71780
rect 7720 71836 7784 71840
rect 7720 71780 7724 71836
rect 7724 71780 7780 71836
rect 7780 71780 7784 71836
rect 7720 71776 7784 71780
rect 2584 71292 2648 71296
rect 2584 71236 2588 71292
rect 2588 71236 2644 71292
rect 2644 71236 2648 71292
rect 2584 71232 2648 71236
rect 2664 71292 2728 71296
rect 2664 71236 2668 71292
rect 2668 71236 2724 71292
rect 2724 71236 2728 71292
rect 2664 71232 2728 71236
rect 2744 71292 2808 71296
rect 2744 71236 2748 71292
rect 2748 71236 2804 71292
rect 2804 71236 2808 71292
rect 2744 71232 2808 71236
rect 2824 71292 2888 71296
rect 2824 71236 2828 71292
rect 2828 71236 2884 71292
rect 2884 71236 2888 71292
rect 2824 71232 2888 71236
rect 5848 71292 5912 71296
rect 5848 71236 5852 71292
rect 5852 71236 5908 71292
rect 5908 71236 5912 71292
rect 5848 71232 5912 71236
rect 5928 71292 5992 71296
rect 5928 71236 5932 71292
rect 5932 71236 5988 71292
rect 5988 71236 5992 71292
rect 5928 71232 5992 71236
rect 6008 71292 6072 71296
rect 6008 71236 6012 71292
rect 6012 71236 6068 71292
rect 6068 71236 6072 71292
rect 6008 71232 6072 71236
rect 6088 71292 6152 71296
rect 6088 71236 6092 71292
rect 6092 71236 6148 71292
rect 6148 71236 6152 71292
rect 6088 71232 6152 71236
rect 9112 71292 9176 71296
rect 9112 71236 9116 71292
rect 9116 71236 9172 71292
rect 9172 71236 9176 71292
rect 9112 71232 9176 71236
rect 9192 71292 9256 71296
rect 9192 71236 9196 71292
rect 9196 71236 9252 71292
rect 9252 71236 9256 71292
rect 9192 71232 9256 71236
rect 9272 71292 9336 71296
rect 9272 71236 9276 71292
rect 9276 71236 9332 71292
rect 9332 71236 9336 71292
rect 9272 71232 9336 71236
rect 9352 71292 9416 71296
rect 9352 71236 9356 71292
rect 9356 71236 9412 71292
rect 9412 71236 9416 71292
rect 9352 71232 9416 71236
rect 4216 70748 4280 70752
rect 4216 70692 4220 70748
rect 4220 70692 4276 70748
rect 4276 70692 4280 70748
rect 4216 70688 4280 70692
rect 4296 70748 4360 70752
rect 4296 70692 4300 70748
rect 4300 70692 4356 70748
rect 4356 70692 4360 70748
rect 4296 70688 4360 70692
rect 4376 70748 4440 70752
rect 4376 70692 4380 70748
rect 4380 70692 4436 70748
rect 4436 70692 4440 70748
rect 4376 70688 4440 70692
rect 4456 70748 4520 70752
rect 4456 70692 4460 70748
rect 4460 70692 4516 70748
rect 4516 70692 4520 70748
rect 4456 70688 4520 70692
rect 7480 70748 7544 70752
rect 7480 70692 7484 70748
rect 7484 70692 7540 70748
rect 7540 70692 7544 70748
rect 7480 70688 7544 70692
rect 7560 70748 7624 70752
rect 7560 70692 7564 70748
rect 7564 70692 7620 70748
rect 7620 70692 7624 70748
rect 7560 70688 7624 70692
rect 7640 70748 7704 70752
rect 7640 70692 7644 70748
rect 7644 70692 7700 70748
rect 7700 70692 7704 70748
rect 7640 70688 7704 70692
rect 7720 70748 7784 70752
rect 7720 70692 7724 70748
rect 7724 70692 7780 70748
rect 7780 70692 7784 70748
rect 7720 70688 7784 70692
rect 2268 70620 2332 70684
rect 1532 70408 1596 70412
rect 1532 70352 1546 70408
rect 1546 70352 1596 70408
rect 1532 70348 1596 70352
rect 1900 70272 1964 70276
rect 1900 70216 1950 70272
rect 1950 70216 1964 70272
rect 1900 70212 1964 70216
rect 2268 70272 2332 70276
rect 2268 70216 2318 70272
rect 2318 70216 2332 70272
rect 2268 70212 2332 70216
rect 2584 70204 2648 70208
rect 2584 70148 2588 70204
rect 2588 70148 2644 70204
rect 2644 70148 2648 70204
rect 2584 70144 2648 70148
rect 2664 70204 2728 70208
rect 2664 70148 2668 70204
rect 2668 70148 2724 70204
rect 2724 70148 2728 70204
rect 2664 70144 2728 70148
rect 2744 70204 2808 70208
rect 2744 70148 2748 70204
rect 2748 70148 2804 70204
rect 2804 70148 2808 70204
rect 2744 70144 2808 70148
rect 2824 70204 2888 70208
rect 2824 70148 2828 70204
rect 2828 70148 2884 70204
rect 2884 70148 2888 70204
rect 2824 70144 2888 70148
rect 5848 70204 5912 70208
rect 5848 70148 5852 70204
rect 5852 70148 5908 70204
rect 5908 70148 5912 70204
rect 5848 70144 5912 70148
rect 5928 70204 5992 70208
rect 5928 70148 5932 70204
rect 5932 70148 5988 70204
rect 5988 70148 5992 70204
rect 5928 70144 5992 70148
rect 6008 70204 6072 70208
rect 6008 70148 6012 70204
rect 6012 70148 6068 70204
rect 6068 70148 6072 70204
rect 6008 70144 6072 70148
rect 6088 70204 6152 70208
rect 6088 70148 6092 70204
rect 6092 70148 6148 70204
rect 6148 70148 6152 70204
rect 6088 70144 6152 70148
rect 9112 70204 9176 70208
rect 9112 70148 9116 70204
rect 9116 70148 9172 70204
rect 9172 70148 9176 70204
rect 9112 70144 9176 70148
rect 9192 70204 9256 70208
rect 9192 70148 9196 70204
rect 9196 70148 9252 70204
rect 9252 70148 9256 70204
rect 9192 70144 9256 70148
rect 9272 70204 9336 70208
rect 9272 70148 9276 70204
rect 9276 70148 9332 70204
rect 9332 70148 9336 70204
rect 9272 70144 9336 70148
rect 9352 70204 9416 70208
rect 9352 70148 9356 70204
rect 9356 70148 9412 70204
rect 9412 70148 9416 70204
rect 9352 70144 9416 70148
rect 2268 70076 2332 70140
rect 1348 70000 1412 70004
rect 1348 69944 1398 70000
rect 1398 69944 1412 70000
rect 1348 69940 1412 69944
rect 4216 69660 4280 69664
rect 4216 69604 4220 69660
rect 4220 69604 4276 69660
rect 4276 69604 4280 69660
rect 4216 69600 4280 69604
rect 4296 69660 4360 69664
rect 4296 69604 4300 69660
rect 4300 69604 4356 69660
rect 4356 69604 4360 69660
rect 4296 69600 4360 69604
rect 4376 69660 4440 69664
rect 4376 69604 4380 69660
rect 4380 69604 4436 69660
rect 4436 69604 4440 69660
rect 4376 69600 4440 69604
rect 4456 69660 4520 69664
rect 4456 69604 4460 69660
rect 4460 69604 4516 69660
rect 4516 69604 4520 69660
rect 4456 69600 4520 69604
rect 7480 69660 7544 69664
rect 7480 69604 7484 69660
rect 7484 69604 7540 69660
rect 7540 69604 7544 69660
rect 7480 69600 7544 69604
rect 7560 69660 7624 69664
rect 7560 69604 7564 69660
rect 7564 69604 7620 69660
rect 7620 69604 7624 69660
rect 7560 69600 7624 69604
rect 7640 69660 7704 69664
rect 7640 69604 7644 69660
rect 7644 69604 7700 69660
rect 7700 69604 7704 69660
rect 7640 69600 7704 69604
rect 7720 69660 7784 69664
rect 7720 69604 7724 69660
rect 7724 69604 7780 69660
rect 7780 69604 7784 69660
rect 7720 69600 7784 69604
rect 2584 69116 2648 69120
rect 2584 69060 2588 69116
rect 2588 69060 2644 69116
rect 2644 69060 2648 69116
rect 2584 69056 2648 69060
rect 2664 69116 2728 69120
rect 2664 69060 2668 69116
rect 2668 69060 2724 69116
rect 2724 69060 2728 69116
rect 2664 69056 2728 69060
rect 2744 69116 2808 69120
rect 2744 69060 2748 69116
rect 2748 69060 2804 69116
rect 2804 69060 2808 69116
rect 2744 69056 2808 69060
rect 2824 69116 2888 69120
rect 2824 69060 2828 69116
rect 2828 69060 2884 69116
rect 2884 69060 2888 69116
rect 2824 69056 2888 69060
rect 5848 69116 5912 69120
rect 5848 69060 5852 69116
rect 5852 69060 5908 69116
rect 5908 69060 5912 69116
rect 5848 69056 5912 69060
rect 5928 69116 5992 69120
rect 5928 69060 5932 69116
rect 5932 69060 5988 69116
rect 5988 69060 5992 69116
rect 5928 69056 5992 69060
rect 6008 69116 6072 69120
rect 6008 69060 6012 69116
rect 6012 69060 6068 69116
rect 6068 69060 6072 69116
rect 6008 69056 6072 69060
rect 6088 69116 6152 69120
rect 6088 69060 6092 69116
rect 6092 69060 6148 69116
rect 6148 69060 6152 69116
rect 6088 69056 6152 69060
rect 9112 69116 9176 69120
rect 9112 69060 9116 69116
rect 9116 69060 9172 69116
rect 9172 69060 9176 69116
rect 9112 69056 9176 69060
rect 9192 69116 9256 69120
rect 9192 69060 9196 69116
rect 9196 69060 9252 69116
rect 9252 69060 9256 69116
rect 9192 69056 9256 69060
rect 9272 69116 9336 69120
rect 9272 69060 9276 69116
rect 9276 69060 9332 69116
rect 9332 69060 9336 69116
rect 9272 69056 9336 69060
rect 9352 69116 9416 69120
rect 9352 69060 9356 69116
rect 9356 69060 9412 69116
rect 9412 69060 9416 69116
rect 9352 69056 9416 69060
rect 4216 68572 4280 68576
rect 4216 68516 4220 68572
rect 4220 68516 4276 68572
rect 4276 68516 4280 68572
rect 4216 68512 4280 68516
rect 4296 68572 4360 68576
rect 4296 68516 4300 68572
rect 4300 68516 4356 68572
rect 4356 68516 4360 68572
rect 4296 68512 4360 68516
rect 4376 68572 4440 68576
rect 4376 68516 4380 68572
rect 4380 68516 4436 68572
rect 4436 68516 4440 68572
rect 4376 68512 4440 68516
rect 4456 68572 4520 68576
rect 4456 68516 4460 68572
rect 4460 68516 4516 68572
rect 4516 68516 4520 68572
rect 4456 68512 4520 68516
rect 7480 68572 7544 68576
rect 7480 68516 7484 68572
rect 7484 68516 7540 68572
rect 7540 68516 7544 68572
rect 7480 68512 7544 68516
rect 7560 68572 7624 68576
rect 7560 68516 7564 68572
rect 7564 68516 7620 68572
rect 7620 68516 7624 68572
rect 7560 68512 7624 68516
rect 7640 68572 7704 68576
rect 7640 68516 7644 68572
rect 7644 68516 7700 68572
rect 7700 68516 7704 68572
rect 7640 68512 7704 68516
rect 7720 68572 7784 68576
rect 7720 68516 7724 68572
rect 7724 68516 7780 68572
rect 7780 68516 7784 68572
rect 7720 68512 7784 68516
rect 2584 68028 2648 68032
rect 2584 67972 2588 68028
rect 2588 67972 2644 68028
rect 2644 67972 2648 68028
rect 2584 67968 2648 67972
rect 2664 68028 2728 68032
rect 2664 67972 2668 68028
rect 2668 67972 2724 68028
rect 2724 67972 2728 68028
rect 2664 67968 2728 67972
rect 2744 68028 2808 68032
rect 2744 67972 2748 68028
rect 2748 67972 2804 68028
rect 2804 67972 2808 68028
rect 2744 67968 2808 67972
rect 2824 68028 2888 68032
rect 2824 67972 2828 68028
rect 2828 67972 2884 68028
rect 2884 67972 2888 68028
rect 2824 67968 2888 67972
rect 5848 68028 5912 68032
rect 5848 67972 5852 68028
rect 5852 67972 5908 68028
rect 5908 67972 5912 68028
rect 5848 67968 5912 67972
rect 5928 68028 5992 68032
rect 5928 67972 5932 68028
rect 5932 67972 5988 68028
rect 5988 67972 5992 68028
rect 5928 67968 5992 67972
rect 6008 68028 6072 68032
rect 6008 67972 6012 68028
rect 6012 67972 6068 68028
rect 6068 67972 6072 68028
rect 6008 67968 6072 67972
rect 6088 68028 6152 68032
rect 6088 67972 6092 68028
rect 6092 67972 6148 68028
rect 6148 67972 6152 68028
rect 6088 67968 6152 67972
rect 9112 68028 9176 68032
rect 9112 67972 9116 68028
rect 9116 67972 9172 68028
rect 9172 67972 9176 68028
rect 9112 67968 9176 67972
rect 9192 68028 9256 68032
rect 9192 67972 9196 68028
rect 9196 67972 9252 68028
rect 9252 67972 9256 68028
rect 9192 67968 9256 67972
rect 9272 68028 9336 68032
rect 9272 67972 9276 68028
rect 9276 67972 9332 68028
rect 9332 67972 9336 68028
rect 9272 67968 9336 67972
rect 9352 68028 9416 68032
rect 9352 67972 9356 68028
rect 9356 67972 9412 68028
rect 9412 67972 9416 68028
rect 9352 67968 9416 67972
rect 4216 67484 4280 67488
rect 4216 67428 4220 67484
rect 4220 67428 4276 67484
rect 4276 67428 4280 67484
rect 4216 67424 4280 67428
rect 4296 67484 4360 67488
rect 4296 67428 4300 67484
rect 4300 67428 4356 67484
rect 4356 67428 4360 67484
rect 4296 67424 4360 67428
rect 4376 67484 4440 67488
rect 4376 67428 4380 67484
rect 4380 67428 4436 67484
rect 4436 67428 4440 67484
rect 4376 67424 4440 67428
rect 4456 67484 4520 67488
rect 4456 67428 4460 67484
rect 4460 67428 4516 67484
rect 4516 67428 4520 67484
rect 4456 67424 4520 67428
rect 7480 67484 7544 67488
rect 7480 67428 7484 67484
rect 7484 67428 7540 67484
rect 7540 67428 7544 67484
rect 7480 67424 7544 67428
rect 7560 67484 7624 67488
rect 7560 67428 7564 67484
rect 7564 67428 7620 67484
rect 7620 67428 7624 67484
rect 7560 67424 7624 67428
rect 7640 67484 7704 67488
rect 7640 67428 7644 67484
rect 7644 67428 7700 67484
rect 7700 67428 7704 67484
rect 7640 67424 7704 67428
rect 7720 67484 7784 67488
rect 7720 67428 7724 67484
rect 7724 67428 7780 67484
rect 7780 67428 7784 67484
rect 7720 67424 7784 67428
rect 2584 66940 2648 66944
rect 2584 66884 2588 66940
rect 2588 66884 2644 66940
rect 2644 66884 2648 66940
rect 2584 66880 2648 66884
rect 2664 66940 2728 66944
rect 2664 66884 2668 66940
rect 2668 66884 2724 66940
rect 2724 66884 2728 66940
rect 2664 66880 2728 66884
rect 2744 66940 2808 66944
rect 2744 66884 2748 66940
rect 2748 66884 2804 66940
rect 2804 66884 2808 66940
rect 2744 66880 2808 66884
rect 2824 66940 2888 66944
rect 2824 66884 2828 66940
rect 2828 66884 2884 66940
rect 2884 66884 2888 66940
rect 2824 66880 2888 66884
rect 5848 66940 5912 66944
rect 5848 66884 5852 66940
rect 5852 66884 5908 66940
rect 5908 66884 5912 66940
rect 5848 66880 5912 66884
rect 5928 66940 5992 66944
rect 5928 66884 5932 66940
rect 5932 66884 5988 66940
rect 5988 66884 5992 66940
rect 5928 66880 5992 66884
rect 6008 66940 6072 66944
rect 6008 66884 6012 66940
rect 6012 66884 6068 66940
rect 6068 66884 6072 66940
rect 6008 66880 6072 66884
rect 6088 66940 6152 66944
rect 6088 66884 6092 66940
rect 6092 66884 6148 66940
rect 6148 66884 6152 66940
rect 6088 66880 6152 66884
rect 9112 66940 9176 66944
rect 9112 66884 9116 66940
rect 9116 66884 9172 66940
rect 9172 66884 9176 66940
rect 9112 66880 9176 66884
rect 9192 66940 9256 66944
rect 9192 66884 9196 66940
rect 9196 66884 9252 66940
rect 9252 66884 9256 66940
rect 9192 66880 9256 66884
rect 9272 66940 9336 66944
rect 9272 66884 9276 66940
rect 9276 66884 9332 66940
rect 9332 66884 9336 66940
rect 9272 66880 9336 66884
rect 9352 66940 9416 66944
rect 9352 66884 9356 66940
rect 9356 66884 9412 66940
rect 9412 66884 9416 66940
rect 9352 66880 9416 66884
rect 4216 66396 4280 66400
rect 4216 66340 4220 66396
rect 4220 66340 4276 66396
rect 4276 66340 4280 66396
rect 4216 66336 4280 66340
rect 4296 66396 4360 66400
rect 4296 66340 4300 66396
rect 4300 66340 4356 66396
rect 4356 66340 4360 66396
rect 4296 66336 4360 66340
rect 4376 66396 4440 66400
rect 4376 66340 4380 66396
rect 4380 66340 4436 66396
rect 4436 66340 4440 66396
rect 4376 66336 4440 66340
rect 4456 66396 4520 66400
rect 4456 66340 4460 66396
rect 4460 66340 4516 66396
rect 4516 66340 4520 66396
rect 4456 66336 4520 66340
rect 7480 66396 7544 66400
rect 7480 66340 7484 66396
rect 7484 66340 7540 66396
rect 7540 66340 7544 66396
rect 7480 66336 7544 66340
rect 7560 66396 7624 66400
rect 7560 66340 7564 66396
rect 7564 66340 7620 66396
rect 7620 66340 7624 66396
rect 7560 66336 7624 66340
rect 7640 66396 7704 66400
rect 7640 66340 7644 66396
rect 7644 66340 7700 66396
rect 7700 66340 7704 66396
rect 7640 66336 7704 66340
rect 7720 66396 7784 66400
rect 7720 66340 7724 66396
rect 7724 66340 7780 66396
rect 7780 66340 7784 66396
rect 7720 66336 7784 66340
rect 1532 66268 1596 66332
rect 3740 65996 3804 66060
rect 2584 65852 2648 65856
rect 2584 65796 2588 65852
rect 2588 65796 2644 65852
rect 2644 65796 2648 65852
rect 2584 65792 2648 65796
rect 2664 65852 2728 65856
rect 2664 65796 2668 65852
rect 2668 65796 2724 65852
rect 2724 65796 2728 65852
rect 2664 65792 2728 65796
rect 2744 65852 2808 65856
rect 2744 65796 2748 65852
rect 2748 65796 2804 65852
rect 2804 65796 2808 65852
rect 2744 65792 2808 65796
rect 2824 65852 2888 65856
rect 2824 65796 2828 65852
rect 2828 65796 2884 65852
rect 2884 65796 2888 65852
rect 2824 65792 2888 65796
rect 5848 65852 5912 65856
rect 5848 65796 5852 65852
rect 5852 65796 5908 65852
rect 5908 65796 5912 65852
rect 5848 65792 5912 65796
rect 5928 65852 5992 65856
rect 5928 65796 5932 65852
rect 5932 65796 5988 65852
rect 5988 65796 5992 65852
rect 5928 65792 5992 65796
rect 6008 65852 6072 65856
rect 6008 65796 6012 65852
rect 6012 65796 6068 65852
rect 6068 65796 6072 65852
rect 6008 65792 6072 65796
rect 6088 65852 6152 65856
rect 6088 65796 6092 65852
rect 6092 65796 6148 65852
rect 6148 65796 6152 65852
rect 6088 65792 6152 65796
rect 9112 65852 9176 65856
rect 9112 65796 9116 65852
rect 9116 65796 9172 65852
rect 9172 65796 9176 65852
rect 9112 65792 9176 65796
rect 9192 65852 9256 65856
rect 9192 65796 9196 65852
rect 9196 65796 9252 65852
rect 9252 65796 9256 65852
rect 9192 65792 9256 65796
rect 9272 65852 9336 65856
rect 9272 65796 9276 65852
rect 9276 65796 9332 65852
rect 9332 65796 9336 65852
rect 9272 65792 9336 65796
rect 9352 65852 9416 65856
rect 9352 65796 9356 65852
rect 9356 65796 9412 65852
rect 9412 65796 9416 65852
rect 9352 65792 9416 65796
rect 4216 65308 4280 65312
rect 4216 65252 4220 65308
rect 4220 65252 4276 65308
rect 4276 65252 4280 65308
rect 4216 65248 4280 65252
rect 4296 65308 4360 65312
rect 4296 65252 4300 65308
rect 4300 65252 4356 65308
rect 4356 65252 4360 65308
rect 4296 65248 4360 65252
rect 4376 65308 4440 65312
rect 4376 65252 4380 65308
rect 4380 65252 4436 65308
rect 4436 65252 4440 65308
rect 4376 65248 4440 65252
rect 4456 65308 4520 65312
rect 4456 65252 4460 65308
rect 4460 65252 4516 65308
rect 4516 65252 4520 65308
rect 4456 65248 4520 65252
rect 7480 65308 7544 65312
rect 7480 65252 7484 65308
rect 7484 65252 7540 65308
rect 7540 65252 7544 65308
rect 7480 65248 7544 65252
rect 7560 65308 7624 65312
rect 7560 65252 7564 65308
rect 7564 65252 7620 65308
rect 7620 65252 7624 65308
rect 7560 65248 7624 65252
rect 7640 65308 7704 65312
rect 7640 65252 7644 65308
rect 7644 65252 7700 65308
rect 7700 65252 7704 65308
rect 7640 65248 7704 65252
rect 7720 65308 7784 65312
rect 7720 65252 7724 65308
rect 7724 65252 7780 65308
rect 7780 65252 7784 65308
rect 7720 65248 7784 65252
rect 3556 65044 3620 65108
rect 1716 64968 1780 64972
rect 1716 64912 1730 64968
rect 1730 64912 1780 64968
rect 1716 64908 1780 64912
rect 2584 64764 2648 64768
rect 2584 64708 2588 64764
rect 2588 64708 2644 64764
rect 2644 64708 2648 64764
rect 2584 64704 2648 64708
rect 2664 64764 2728 64768
rect 2664 64708 2668 64764
rect 2668 64708 2724 64764
rect 2724 64708 2728 64764
rect 2664 64704 2728 64708
rect 2744 64764 2808 64768
rect 2744 64708 2748 64764
rect 2748 64708 2804 64764
rect 2804 64708 2808 64764
rect 2744 64704 2808 64708
rect 2824 64764 2888 64768
rect 2824 64708 2828 64764
rect 2828 64708 2884 64764
rect 2884 64708 2888 64764
rect 2824 64704 2888 64708
rect 5848 64764 5912 64768
rect 5848 64708 5852 64764
rect 5852 64708 5908 64764
rect 5908 64708 5912 64764
rect 5848 64704 5912 64708
rect 5928 64764 5992 64768
rect 5928 64708 5932 64764
rect 5932 64708 5988 64764
rect 5988 64708 5992 64764
rect 5928 64704 5992 64708
rect 6008 64764 6072 64768
rect 6008 64708 6012 64764
rect 6012 64708 6068 64764
rect 6068 64708 6072 64764
rect 6008 64704 6072 64708
rect 6088 64764 6152 64768
rect 6088 64708 6092 64764
rect 6092 64708 6148 64764
rect 6148 64708 6152 64764
rect 6088 64704 6152 64708
rect 9112 64764 9176 64768
rect 9112 64708 9116 64764
rect 9116 64708 9172 64764
rect 9172 64708 9176 64764
rect 9112 64704 9176 64708
rect 9192 64764 9256 64768
rect 9192 64708 9196 64764
rect 9196 64708 9252 64764
rect 9252 64708 9256 64764
rect 9192 64704 9256 64708
rect 9272 64764 9336 64768
rect 9272 64708 9276 64764
rect 9276 64708 9332 64764
rect 9332 64708 9336 64764
rect 9272 64704 9336 64708
rect 9352 64764 9416 64768
rect 9352 64708 9356 64764
rect 9356 64708 9412 64764
rect 9412 64708 9416 64764
rect 9352 64704 9416 64708
rect 4216 64220 4280 64224
rect 4216 64164 4220 64220
rect 4220 64164 4276 64220
rect 4276 64164 4280 64220
rect 4216 64160 4280 64164
rect 4296 64220 4360 64224
rect 4296 64164 4300 64220
rect 4300 64164 4356 64220
rect 4356 64164 4360 64220
rect 4296 64160 4360 64164
rect 4376 64220 4440 64224
rect 4376 64164 4380 64220
rect 4380 64164 4436 64220
rect 4436 64164 4440 64220
rect 4376 64160 4440 64164
rect 4456 64220 4520 64224
rect 4456 64164 4460 64220
rect 4460 64164 4516 64220
rect 4516 64164 4520 64220
rect 4456 64160 4520 64164
rect 7480 64220 7544 64224
rect 7480 64164 7484 64220
rect 7484 64164 7540 64220
rect 7540 64164 7544 64220
rect 7480 64160 7544 64164
rect 7560 64220 7624 64224
rect 7560 64164 7564 64220
rect 7564 64164 7620 64220
rect 7620 64164 7624 64220
rect 7560 64160 7624 64164
rect 7640 64220 7704 64224
rect 7640 64164 7644 64220
rect 7644 64164 7700 64220
rect 7700 64164 7704 64220
rect 7640 64160 7704 64164
rect 7720 64220 7784 64224
rect 7720 64164 7724 64220
rect 7724 64164 7780 64220
rect 7780 64164 7784 64220
rect 7720 64160 7784 64164
rect 3004 63820 3068 63884
rect 2584 63676 2648 63680
rect 2584 63620 2588 63676
rect 2588 63620 2644 63676
rect 2644 63620 2648 63676
rect 2584 63616 2648 63620
rect 2664 63676 2728 63680
rect 2664 63620 2668 63676
rect 2668 63620 2724 63676
rect 2724 63620 2728 63676
rect 2664 63616 2728 63620
rect 2744 63676 2808 63680
rect 2744 63620 2748 63676
rect 2748 63620 2804 63676
rect 2804 63620 2808 63676
rect 2744 63616 2808 63620
rect 2824 63676 2888 63680
rect 2824 63620 2828 63676
rect 2828 63620 2884 63676
rect 2884 63620 2888 63676
rect 2824 63616 2888 63620
rect 5848 63676 5912 63680
rect 5848 63620 5852 63676
rect 5852 63620 5908 63676
rect 5908 63620 5912 63676
rect 5848 63616 5912 63620
rect 5928 63676 5992 63680
rect 5928 63620 5932 63676
rect 5932 63620 5988 63676
rect 5988 63620 5992 63676
rect 5928 63616 5992 63620
rect 6008 63676 6072 63680
rect 6008 63620 6012 63676
rect 6012 63620 6068 63676
rect 6068 63620 6072 63676
rect 6008 63616 6072 63620
rect 6088 63676 6152 63680
rect 6088 63620 6092 63676
rect 6092 63620 6148 63676
rect 6148 63620 6152 63676
rect 6088 63616 6152 63620
rect 9112 63676 9176 63680
rect 9112 63620 9116 63676
rect 9116 63620 9172 63676
rect 9172 63620 9176 63676
rect 9112 63616 9176 63620
rect 9192 63676 9256 63680
rect 9192 63620 9196 63676
rect 9196 63620 9252 63676
rect 9252 63620 9256 63676
rect 9192 63616 9256 63620
rect 9272 63676 9336 63680
rect 9272 63620 9276 63676
rect 9276 63620 9332 63676
rect 9332 63620 9336 63676
rect 9272 63616 9336 63620
rect 9352 63676 9416 63680
rect 9352 63620 9356 63676
rect 9356 63620 9412 63676
rect 9412 63620 9416 63676
rect 9352 63616 9416 63620
rect 4216 63132 4280 63136
rect 4216 63076 4220 63132
rect 4220 63076 4276 63132
rect 4276 63076 4280 63132
rect 4216 63072 4280 63076
rect 4296 63132 4360 63136
rect 4296 63076 4300 63132
rect 4300 63076 4356 63132
rect 4356 63076 4360 63132
rect 4296 63072 4360 63076
rect 4376 63132 4440 63136
rect 4376 63076 4380 63132
rect 4380 63076 4436 63132
rect 4436 63076 4440 63132
rect 4376 63072 4440 63076
rect 4456 63132 4520 63136
rect 4456 63076 4460 63132
rect 4460 63076 4516 63132
rect 4516 63076 4520 63132
rect 4456 63072 4520 63076
rect 7480 63132 7544 63136
rect 7480 63076 7484 63132
rect 7484 63076 7540 63132
rect 7540 63076 7544 63132
rect 7480 63072 7544 63076
rect 7560 63132 7624 63136
rect 7560 63076 7564 63132
rect 7564 63076 7620 63132
rect 7620 63076 7624 63132
rect 7560 63072 7624 63076
rect 7640 63132 7704 63136
rect 7640 63076 7644 63132
rect 7644 63076 7700 63132
rect 7700 63076 7704 63132
rect 7640 63072 7704 63076
rect 7720 63132 7784 63136
rect 7720 63076 7724 63132
rect 7724 63076 7780 63132
rect 7780 63076 7784 63132
rect 7720 63072 7784 63076
rect 2268 62868 2332 62932
rect 1900 62596 1964 62660
rect 2584 62588 2648 62592
rect 2584 62532 2588 62588
rect 2588 62532 2644 62588
rect 2644 62532 2648 62588
rect 2584 62528 2648 62532
rect 2664 62588 2728 62592
rect 2664 62532 2668 62588
rect 2668 62532 2724 62588
rect 2724 62532 2728 62588
rect 2664 62528 2728 62532
rect 2744 62588 2808 62592
rect 2744 62532 2748 62588
rect 2748 62532 2804 62588
rect 2804 62532 2808 62588
rect 2744 62528 2808 62532
rect 2824 62588 2888 62592
rect 2824 62532 2828 62588
rect 2828 62532 2884 62588
rect 2884 62532 2888 62588
rect 2824 62528 2888 62532
rect 5848 62588 5912 62592
rect 5848 62532 5852 62588
rect 5852 62532 5908 62588
rect 5908 62532 5912 62588
rect 5848 62528 5912 62532
rect 5928 62588 5992 62592
rect 5928 62532 5932 62588
rect 5932 62532 5988 62588
rect 5988 62532 5992 62588
rect 5928 62528 5992 62532
rect 6008 62588 6072 62592
rect 6008 62532 6012 62588
rect 6012 62532 6068 62588
rect 6068 62532 6072 62588
rect 6008 62528 6072 62532
rect 6088 62588 6152 62592
rect 6088 62532 6092 62588
rect 6092 62532 6148 62588
rect 6148 62532 6152 62588
rect 6088 62528 6152 62532
rect 9112 62588 9176 62592
rect 9112 62532 9116 62588
rect 9116 62532 9172 62588
rect 9172 62532 9176 62588
rect 9112 62528 9176 62532
rect 9192 62588 9256 62592
rect 9192 62532 9196 62588
rect 9196 62532 9252 62588
rect 9252 62532 9256 62588
rect 9192 62528 9256 62532
rect 9272 62588 9336 62592
rect 9272 62532 9276 62588
rect 9276 62532 9332 62588
rect 9332 62532 9336 62588
rect 9272 62528 9336 62532
rect 9352 62588 9416 62592
rect 9352 62532 9356 62588
rect 9356 62532 9412 62588
rect 9412 62532 9416 62588
rect 9352 62528 9416 62532
rect 4216 62044 4280 62048
rect 4216 61988 4220 62044
rect 4220 61988 4276 62044
rect 4276 61988 4280 62044
rect 4216 61984 4280 61988
rect 4296 62044 4360 62048
rect 4296 61988 4300 62044
rect 4300 61988 4356 62044
rect 4356 61988 4360 62044
rect 4296 61984 4360 61988
rect 4376 62044 4440 62048
rect 4376 61988 4380 62044
rect 4380 61988 4436 62044
rect 4436 61988 4440 62044
rect 4376 61984 4440 61988
rect 4456 62044 4520 62048
rect 4456 61988 4460 62044
rect 4460 61988 4516 62044
rect 4516 61988 4520 62044
rect 4456 61984 4520 61988
rect 7480 62044 7544 62048
rect 7480 61988 7484 62044
rect 7484 61988 7540 62044
rect 7540 61988 7544 62044
rect 7480 61984 7544 61988
rect 7560 62044 7624 62048
rect 7560 61988 7564 62044
rect 7564 61988 7620 62044
rect 7620 61988 7624 62044
rect 7560 61984 7624 61988
rect 7640 62044 7704 62048
rect 7640 61988 7644 62044
rect 7644 61988 7700 62044
rect 7700 61988 7704 62044
rect 7640 61984 7704 61988
rect 7720 62044 7784 62048
rect 7720 61988 7724 62044
rect 7724 61988 7780 62044
rect 7780 61988 7784 62044
rect 7720 61984 7784 61988
rect 3188 61644 3252 61708
rect 2584 61500 2648 61504
rect 2584 61444 2588 61500
rect 2588 61444 2644 61500
rect 2644 61444 2648 61500
rect 2584 61440 2648 61444
rect 2664 61500 2728 61504
rect 2664 61444 2668 61500
rect 2668 61444 2724 61500
rect 2724 61444 2728 61500
rect 2664 61440 2728 61444
rect 2744 61500 2808 61504
rect 2744 61444 2748 61500
rect 2748 61444 2804 61500
rect 2804 61444 2808 61500
rect 2744 61440 2808 61444
rect 2824 61500 2888 61504
rect 2824 61444 2828 61500
rect 2828 61444 2884 61500
rect 2884 61444 2888 61500
rect 2824 61440 2888 61444
rect 5848 61500 5912 61504
rect 5848 61444 5852 61500
rect 5852 61444 5908 61500
rect 5908 61444 5912 61500
rect 5848 61440 5912 61444
rect 5928 61500 5992 61504
rect 5928 61444 5932 61500
rect 5932 61444 5988 61500
rect 5988 61444 5992 61500
rect 5928 61440 5992 61444
rect 6008 61500 6072 61504
rect 6008 61444 6012 61500
rect 6012 61444 6068 61500
rect 6068 61444 6072 61500
rect 6008 61440 6072 61444
rect 6088 61500 6152 61504
rect 6088 61444 6092 61500
rect 6092 61444 6148 61500
rect 6148 61444 6152 61500
rect 6088 61440 6152 61444
rect 9112 61500 9176 61504
rect 9112 61444 9116 61500
rect 9116 61444 9172 61500
rect 9172 61444 9176 61500
rect 9112 61440 9176 61444
rect 9192 61500 9256 61504
rect 9192 61444 9196 61500
rect 9196 61444 9252 61500
rect 9252 61444 9256 61500
rect 9192 61440 9256 61444
rect 9272 61500 9336 61504
rect 9272 61444 9276 61500
rect 9276 61444 9332 61500
rect 9332 61444 9336 61500
rect 9272 61440 9336 61444
rect 9352 61500 9416 61504
rect 9352 61444 9356 61500
rect 9356 61444 9412 61500
rect 9412 61444 9416 61500
rect 9352 61440 9416 61444
rect 2268 61100 2332 61164
rect 4216 60956 4280 60960
rect 4216 60900 4220 60956
rect 4220 60900 4276 60956
rect 4276 60900 4280 60956
rect 4216 60896 4280 60900
rect 4296 60956 4360 60960
rect 4296 60900 4300 60956
rect 4300 60900 4356 60956
rect 4356 60900 4360 60956
rect 4296 60896 4360 60900
rect 4376 60956 4440 60960
rect 4376 60900 4380 60956
rect 4380 60900 4436 60956
rect 4436 60900 4440 60956
rect 4376 60896 4440 60900
rect 4456 60956 4520 60960
rect 4456 60900 4460 60956
rect 4460 60900 4516 60956
rect 4516 60900 4520 60956
rect 4456 60896 4520 60900
rect 7480 60956 7544 60960
rect 7480 60900 7484 60956
rect 7484 60900 7540 60956
rect 7540 60900 7544 60956
rect 7480 60896 7544 60900
rect 7560 60956 7624 60960
rect 7560 60900 7564 60956
rect 7564 60900 7620 60956
rect 7620 60900 7624 60956
rect 7560 60896 7624 60900
rect 7640 60956 7704 60960
rect 7640 60900 7644 60956
rect 7644 60900 7700 60956
rect 7700 60900 7704 60956
rect 7640 60896 7704 60900
rect 7720 60956 7784 60960
rect 7720 60900 7724 60956
rect 7724 60900 7780 60956
rect 7780 60900 7784 60956
rect 7720 60896 7784 60900
rect 3188 60828 3252 60892
rect 3924 60888 3988 60892
rect 3924 60832 3974 60888
rect 3974 60832 3988 60888
rect 3924 60828 3988 60832
rect 3924 60616 3988 60620
rect 3924 60560 3974 60616
rect 3974 60560 3988 60616
rect 3924 60556 3988 60560
rect 2268 60420 2332 60484
rect 2584 60412 2648 60416
rect 2584 60356 2588 60412
rect 2588 60356 2644 60412
rect 2644 60356 2648 60412
rect 2584 60352 2648 60356
rect 2664 60412 2728 60416
rect 2664 60356 2668 60412
rect 2668 60356 2724 60412
rect 2724 60356 2728 60412
rect 2664 60352 2728 60356
rect 2744 60412 2808 60416
rect 2744 60356 2748 60412
rect 2748 60356 2804 60412
rect 2804 60356 2808 60412
rect 2744 60352 2808 60356
rect 2824 60412 2888 60416
rect 2824 60356 2828 60412
rect 2828 60356 2884 60412
rect 2884 60356 2888 60412
rect 2824 60352 2888 60356
rect 5848 60412 5912 60416
rect 5848 60356 5852 60412
rect 5852 60356 5908 60412
rect 5908 60356 5912 60412
rect 5848 60352 5912 60356
rect 5928 60412 5992 60416
rect 5928 60356 5932 60412
rect 5932 60356 5988 60412
rect 5988 60356 5992 60412
rect 5928 60352 5992 60356
rect 6008 60412 6072 60416
rect 6008 60356 6012 60412
rect 6012 60356 6068 60412
rect 6068 60356 6072 60412
rect 6008 60352 6072 60356
rect 6088 60412 6152 60416
rect 6088 60356 6092 60412
rect 6092 60356 6148 60412
rect 6148 60356 6152 60412
rect 6088 60352 6152 60356
rect 9112 60412 9176 60416
rect 9112 60356 9116 60412
rect 9116 60356 9172 60412
rect 9172 60356 9176 60412
rect 9112 60352 9176 60356
rect 9192 60412 9256 60416
rect 9192 60356 9196 60412
rect 9196 60356 9252 60412
rect 9252 60356 9256 60412
rect 9192 60352 9256 60356
rect 9272 60412 9336 60416
rect 9272 60356 9276 60412
rect 9276 60356 9332 60412
rect 9332 60356 9336 60412
rect 9272 60352 9336 60356
rect 9352 60412 9416 60416
rect 9352 60356 9356 60412
rect 9356 60356 9412 60412
rect 9412 60356 9416 60412
rect 9352 60352 9416 60356
rect 1348 60284 1412 60348
rect 2268 60284 2332 60348
rect 2084 60148 2148 60212
rect 2084 60012 2148 60076
rect 3372 59876 3436 59940
rect 4216 59868 4280 59872
rect 4216 59812 4220 59868
rect 4220 59812 4276 59868
rect 4276 59812 4280 59868
rect 4216 59808 4280 59812
rect 4296 59868 4360 59872
rect 4296 59812 4300 59868
rect 4300 59812 4356 59868
rect 4356 59812 4360 59868
rect 4296 59808 4360 59812
rect 4376 59868 4440 59872
rect 4376 59812 4380 59868
rect 4380 59812 4436 59868
rect 4436 59812 4440 59868
rect 4376 59808 4440 59812
rect 4456 59868 4520 59872
rect 4456 59812 4460 59868
rect 4460 59812 4516 59868
rect 4516 59812 4520 59868
rect 4456 59808 4520 59812
rect 7480 59868 7544 59872
rect 7480 59812 7484 59868
rect 7484 59812 7540 59868
rect 7540 59812 7544 59868
rect 7480 59808 7544 59812
rect 7560 59868 7624 59872
rect 7560 59812 7564 59868
rect 7564 59812 7620 59868
rect 7620 59812 7624 59868
rect 7560 59808 7624 59812
rect 7640 59868 7704 59872
rect 7640 59812 7644 59868
rect 7644 59812 7700 59868
rect 7700 59812 7704 59868
rect 7640 59808 7704 59812
rect 7720 59868 7784 59872
rect 7720 59812 7724 59868
rect 7724 59812 7780 59868
rect 7780 59812 7784 59868
rect 7720 59808 7784 59812
rect 2584 59324 2648 59328
rect 2584 59268 2588 59324
rect 2588 59268 2644 59324
rect 2644 59268 2648 59324
rect 2584 59264 2648 59268
rect 2664 59324 2728 59328
rect 2664 59268 2668 59324
rect 2668 59268 2724 59324
rect 2724 59268 2728 59324
rect 2664 59264 2728 59268
rect 2744 59324 2808 59328
rect 2744 59268 2748 59324
rect 2748 59268 2804 59324
rect 2804 59268 2808 59324
rect 2744 59264 2808 59268
rect 2824 59324 2888 59328
rect 2824 59268 2828 59324
rect 2828 59268 2884 59324
rect 2884 59268 2888 59324
rect 2824 59264 2888 59268
rect 5848 59324 5912 59328
rect 5848 59268 5852 59324
rect 5852 59268 5908 59324
rect 5908 59268 5912 59324
rect 5848 59264 5912 59268
rect 5928 59324 5992 59328
rect 5928 59268 5932 59324
rect 5932 59268 5988 59324
rect 5988 59268 5992 59324
rect 5928 59264 5992 59268
rect 6008 59324 6072 59328
rect 6008 59268 6012 59324
rect 6012 59268 6068 59324
rect 6068 59268 6072 59324
rect 6008 59264 6072 59268
rect 6088 59324 6152 59328
rect 6088 59268 6092 59324
rect 6092 59268 6148 59324
rect 6148 59268 6152 59324
rect 6088 59264 6152 59268
rect 9112 59324 9176 59328
rect 9112 59268 9116 59324
rect 9116 59268 9172 59324
rect 9172 59268 9176 59324
rect 9112 59264 9176 59268
rect 9192 59324 9256 59328
rect 9192 59268 9196 59324
rect 9196 59268 9252 59324
rect 9252 59268 9256 59324
rect 9192 59264 9256 59268
rect 9272 59324 9336 59328
rect 9272 59268 9276 59324
rect 9276 59268 9332 59324
rect 9332 59268 9336 59324
rect 9272 59264 9336 59268
rect 9352 59324 9416 59328
rect 9352 59268 9356 59324
rect 9356 59268 9412 59324
rect 9412 59268 9416 59324
rect 9352 59264 9416 59268
rect 3556 59196 3620 59260
rect 3556 59060 3620 59124
rect 4216 58780 4280 58784
rect 4216 58724 4220 58780
rect 4220 58724 4276 58780
rect 4276 58724 4280 58780
rect 4216 58720 4280 58724
rect 4296 58780 4360 58784
rect 4296 58724 4300 58780
rect 4300 58724 4356 58780
rect 4356 58724 4360 58780
rect 4296 58720 4360 58724
rect 4376 58780 4440 58784
rect 4376 58724 4380 58780
rect 4380 58724 4436 58780
rect 4436 58724 4440 58780
rect 4376 58720 4440 58724
rect 4456 58780 4520 58784
rect 4456 58724 4460 58780
rect 4460 58724 4516 58780
rect 4516 58724 4520 58780
rect 4456 58720 4520 58724
rect 7480 58780 7544 58784
rect 7480 58724 7484 58780
rect 7484 58724 7540 58780
rect 7540 58724 7544 58780
rect 7480 58720 7544 58724
rect 7560 58780 7624 58784
rect 7560 58724 7564 58780
rect 7564 58724 7620 58780
rect 7620 58724 7624 58780
rect 7560 58720 7624 58724
rect 7640 58780 7704 58784
rect 7640 58724 7644 58780
rect 7644 58724 7700 58780
rect 7700 58724 7704 58780
rect 7640 58720 7704 58724
rect 7720 58780 7784 58784
rect 7720 58724 7724 58780
rect 7724 58724 7780 58780
rect 7780 58724 7784 58780
rect 7720 58720 7784 58724
rect 3188 58380 3252 58444
rect 2584 58236 2648 58240
rect 2584 58180 2588 58236
rect 2588 58180 2644 58236
rect 2644 58180 2648 58236
rect 2584 58176 2648 58180
rect 2664 58236 2728 58240
rect 2664 58180 2668 58236
rect 2668 58180 2724 58236
rect 2724 58180 2728 58236
rect 2664 58176 2728 58180
rect 2744 58236 2808 58240
rect 2744 58180 2748 58236
rect 2748 58180 2804 58236
rect 2804 58180 2808 58236
rect 2744 58176 2808 58180
rect 2824 58236 2888 58240
rect 2824 58180 2828 58236
rect 2828 58180 2884 58236
rect 2884 58180 2888 58236
rect 2824 58176 2888 58180
rect 5848 58236 5912 58240
rect 5848 58180 5852 58236
rect 5852 58180 5908 58236
rect 5908 58180 5912 58236
rect 5848 58176 5912 58180
rect 5928 58236 5992 58240
rect 5928 58180 5932 58236
rect 5932 58180 5988 58236
rect 5988 58180 5992 58236
rect 5928 58176 5992 58180
rect 6008 58236 6072 58240
rect 6008 58180 6012 58236
rect 6012 58180 6068 58236
rect 6068 58180 6072 58236
rect 6008 58176 6072 58180
rect 6088 58236 6152 58240
rect 6088 58180 6092 58236
rect 6092 58180 6148 58236
rect 6148 58180 6152 58236
rect 6088 58176 6152 58180
rect 9112 58236 9176 58240
rect 9112 58180 9116 58236
rect 9116 58180 9172 58236
rect 9172 58180 9176 58236
rect 9112 58176 9176 58180
rect 9192 58236 9256 58240
rect 9192 58180 9196 58236
rect 9196 58180 9252 58236
rect 9252 58180 9256 58236
rect 9192 58176 9256 58180
rect 9272 58236 9336 58240
rect 9272 58180 9276 58236
rect 9276 58180 9332 58236
rect 9332 58180 9336 58236
rect 9272 58176 9336 58180
rect 9352 58236 9416 58240
rect 9352 58180 9356 58236
rect 9356 58180 9412 58236
rect 9412 58180 9416 58236
rect 9352 58176 9416 58180
rect 2084 57972 2148 58036
rect 3740 57972 3804 58036
rect 980 57836 1044 57900
rect 1164 57700 1228 57764
rect 3740 57700 3804 57764
rect 4216 57692 4280 57696
rect 4216 57636 4220 57692
rect 4220 57636 4276 57692
rect 4276 57636 4280 57692
rect 4216 57632 4280 57636
rect 4296 57692 4360 57696
rect 4296 57636 4300 57692
rect 4300 57636 4356 57692
rect 4356 57636 4360 57692
rect 4296 57632 4360 57636
rect 4376 57692 4440 57696
rect 4376 57636 4380 57692
rect 4380 57636 4436 57692
rect 4436 57636 4440 57692
rect 4376 57632 4440 57636
rect 4456 57692 4520 57696
rect 4456 57636 4460 57692
rect 4460 57636 4516 57692
rect 4516 57636 4520 57692
rect 4456 57632 4520 57636
rect 7480 57692 7544 57696
rect 7480 57636 7484 57692
rect 7484 57636 7540 57692
rect 7540 57636 7544 57692
rect 7480 57632 7544 57636
rect 7560 57692 7624 57696
rect 7560 57636 7564 57692
rect 7564 57636 7620 57692
rect 7620 57636 7624 57692
rect 7560 57632 7624 57636
rect 7640 57692 7704 57696
rect 7640 57636 7644 57692
rect 7644 57636 7700 57692
rect 7700 57636 7704 57692
rect 7640 57632 7704 57636
rect 7720 57692 7784 57696
rect 7720 57636 7724 57692
rect 7724 57636 7780 57692
rect 7780 57636 7784 57692
rect 7720 57632 7784 57636
rect 2084 57564 2148 57628
rect 3188 57624 3252 57628
rect 3188 57568 3202 57624
rect 3202 57568 3252 57624
rect 3188 57564 3252 57568
rect 1348 57428 1412 57492
rect 1164 57156 1228 57220
rect 1348 57020 1412 57084
rect 5580 57292 5644 57356
rect 2584 57148 2648 57152
rect 2584 57092 2588 57148
rect 2588 57092 2644 57148
rect 2644 57092 2648 57148
rect 2584 57088 2648 57092
rect 2664 57148 2728 57152
rect 2664 57092 2668 57148
rect 2668 57092 2724 57148
rect 2724 57092 2728 57148
rect 2664 57088 2728 57092
rect 2744 57148 2808 57152
rect 2744 57092 2748 57148
rect 2748 57092 2804 57148
rect 2804 57092 2808 57148
rect 2744 57088 2808 57092
rect 2824 57148 2888 57152
rect 2824 57092 2828 57148
rect 2828 57092 2884 57148
rect 2884 57092 2888 57148
rect 2824 57088 2888 57092
rect 5848 57148 5912 57152
rect 5848 57092 5852 57148
rect 5852 57092 5908 57148
rect 5908 57092 5912 57148
rect 5848 57088 5912 57092
rect 5928 57148 5992 57152
rect 5928 57092 5932 57148
rect 5932 57092 5988 57148
rect 5988 57092 5992 57148
rect 5928 57088 5992 57092
rect 6008 57148 6072 57152
rect 6008 57092 6012 57148
rect 6012 57092 6068 57148
rect 6068 57092 6072 57148
rect 6008 57088 6072 57092
rect 6088 57148 6152 57152
rect 6088 57092 6092 57148
rect 6092 57092 6148 57148
rect 6148 57092 6152 57148
rect 6088 57088 6152 57092
rect 9112 57148 9176 57152
rect 9112 57092 9116 57148
rect 9116 57092 9172 57148
rect 9172 57092 9176 57148
rect 9112 57088 9176 57092
rect 9192 57148 9256 57152
rect 9192 57092 9196 57148
rect 9196 57092 9252 57148
rect 9252 57092 9256 57148
rect 9192 57088 9256 57092
rect 9272 57148 9336 57152
rect 9272 57092 9276 57148
rect 9276 57092 9332 57148
rect 9332 57092 9336 57148
rect 9272 57088 9336 57092
rect 9352 57148 9416 57152
rect 9352 57092 9356 57148
rect 9356 57092 9412 57148
rect 9412 57092 9416 57148
rect 9352 57088 9416 57092
rect 796 56884 860 56948
rect 1164 56808 1228 56812
rect 1164 56752 1214 56808
rect 1214 56752 1228 56808
rect 1164 56748 1228 56752
rect 5396 56748 5460 56812
rect 2268 56612 2332 56676
rect 4216 56604 4280 56608
rect 4216 56548 4220 56604
rect 4220 56548 4276 56604
rect 4276 56548 4280 56604
rect 4216 56544 4280 56548
rect 4296 56604 4360 56608
rect 4296 56548 4300 56604
rect 4300 56548 4356 56604
rect 4356 56548 4360 56604
rect 4296 56544 4360 56548
rect 4376 56604 4440 56608
rect 4376 56548 4380 56604
rect 4380 56548 4436 56604
rect 4436 56548 4440 56604
rect 4376 56544 4440 56548
rect 4456 56604 4520 56608
rect 4456 56548 4460 56604
rect 4460 56548 4516 56604
rect 4516 56548 4520 56604
rect 4456 56544 4520 56548
rect 7480 56604 7544 56608
rect 7480 56548 7484 56604
rect 7484 56548 7540 56604
rect 7540 56548 7544 56604
rect 7480 56544 7544 56548
rect 7560 56604 7624 56608
rect 7560 56548 7564 56604
rect 7564 56548 7620 56604
rect 7620 56548 7624 56604
rect 7560 56544 7624 56548
rect 7640 56604 7704 56608
rect 7640 56548 7644 56604
rect 7644 56548 7700 56604
rect 7700 56548 7704 56604
rect 7640 56544 7704 56548
rect 7720 56604 7784 56608
rect 7720 56548 7724 56604
rect 7724 56548 7780 56604
rect 7780 56548 7784 56604
rect 7720 56544 7784 56548
rect 2084 56476 2148 56540
rect 3004 56400 3068 56404
rect 3004 56344 3018 56400
rect 3018 56344 3068 56400
rect 3004 56340 3068 56344
rect 2584 56060 2648 56064
rect 2584 56004 2588 56060
rect 2588 56004 2644 56060
rect 2644 56004 2648 56060
rect 2584 56000 2648 56004
rect 2664 56060 2728 56064
rect 2664 56004 2668 56060
rect 2668 56004 2724 56060
rect 2724 56004 2728 56060
rect 2664 56000 2728 56004
rect 2744 56060 2808 56064
rect 2744 56004 2748 56060
rect 2748 56004 2804 56060
rect 2804 56004 2808 56060
rect 2744 56000 2808 56004
rect 2824 56060 2888 56064
rect 2824 56004 2828 56060
rect 2828 56004 2884 56060
rect 2884 56004 2888 56060
rect 2824 56000 2888 56004
rect 5848 56060 5912 56064
rect 5848 56004 5852 56060
rect 5852 56004 5908 56060
rect 5908 56004 5912 56060
rect 5848 56000 5912 56004
rect 5928 56060 5992 56064
rect 5928 56004 5932 56060
rect 5932 56004 5988 56060
rect 5988 56004 5992 56060
rect 5928 56000 5992 56004
rect 6008 56060 6072 56064
rect 6008 56004 6012 56060
rect 6012 56004 6068 56060
rect 6068 56004 6072 56060
rect 6008 56000 6072 56004
rect 6088 56060 6152 56064
rect 6088 56004 6092 56060
rect 6092 56004 6148 56060
rect 6148 56004 6152 56060
rect 6088 56000 6152 56004
rect 9112 56060 9176 56064
rect 9112 56004 9116 56060
rect 9116 56004 9172 56060
rect 9172 56004 9176 56060
rect 9112 56000 9176 56004
rect 9192 56060 9256 56064
rect 9192 56004 9196 56060
rect 9196 56004 9252 56060
rect 9252 56004 9256 56060
rect 9192 56000 9256 56004
rect 9272 56060 9336 56064
rect 9272 56004 9276 56060
rect 9276 56004 9332 56060
rect 9332 56004 9336 56060
rect 9272 56000 9336 56004
rect 9352 56060 9416 56064
rect 9352 56004 9356 56060
rect 9356 56004 9412 56060
rect 9412 56004 9416 56060
rect 9352 56000 9416 56004
rect 3924 55796 3988 55860
rect 1900 55524 1964 55588
rect 4216 55516 4280 55520
rect 4216 55460 4220 55516
rect 4220 55460 4276 55516
rect 4276 55460 4280 55516
rect 4216 55456 4280 55460
rect 4296 55516 4360 55520
rect 4296 55460 4300 55516
rect 4300 55460 4356 55516
rect 4356 55460 4360 55516
rect 4296 55456 4360 55460
rect 4376 55516 4440 55520
rect 4376 55460 4380 55516
rect 4380 55460 4436 55516
rect 4436 55460 4440 55516
rect 4376 55456 4440 55460
rect 4456 55516 4520 55520
rect 4456 55460 4460 55516
rect 4460 55460 4516 55516
rect 4516 55460 4520 55516
rect 4456 55456 4520 55460
rect 7480 55516 7544 55520
rect 7480 55460 7484 55516
rect 7484 55460 7540 55516
rect 7540 55460 7544 55516
rect 7480 55456 7544 55460
rect 7560 55516 7624 55520
rect 7560 55460 7564 55516
rect 7564 55460 7620 55516
rect 7620 55460 7624 55516
rect 7560 55456 7624 55460
rect 7640 55516 7704 55520
rect 7640 55460 7644 55516
rect 7644 55460 7700 55516
rect 7700 55460 7704 55516
rect 7640 55456 7704 55460
rect 7720 55516 7784 55520
rect 7720 55460 7724 55516
rect 7724 55460 7780 55516
rect 7780 55460 7784 55516
rect 7720 55456 7784 55460
rect 2268 55312 2332 55316
rect 2268 55256 2318 55312
rect 2318 55256 2332 55312
rect 2268 55252 2332 55256
rect 6316 55252 6380 55316
rect 2584 54972 2648 54976
rect 2584 54916 2588 54972
rect 2588 54916 2644 54972
rect 2644 54916 2648 54972
rect 2584 54912 2648 54916
rect 2664 54972 2728 54976
rect 2664 54916 2668 54972
rect 2668 54916 2724 54972
rect 2724 54916 2728 54972
rect 2664 54912 2728 54916
rect 2744 54972 2808 54976
rect 2744 54916 2748 54972
rect 2748 54916 2804 54972
rect 2804 54916 2808 54972
rect 2744 54912 2808 54916
rect 2824 54972 2888 54976
rect 2824 54916 2828 54972
rect 2828 54916 2884 54972
rect 2884 54916 2888 54972
rect 2824 54912 2888 54916
rect 5848 54972 5912 54976
rect 5848 54916 5852 54972
rect 5852 54916 5908 54972
rect 5908 54916 5912 54972
rect 5848 54912 5912 54916
rect 5928 54972 5992 54976
rect 5928 54916 5932 54972
rect 5932 54916 5988 54972
rect 5988 54916 5992 54972
rect 5928 54912 5992 54916
rect 6008 54972 6072 54976
rect 6008 54916 6012 54972
rect 6012 54916 6068 54972
rect 6068 54916 6072 54972
rect 6008 54912 6072 54916
rect 6088 54972 6152 54976
rect 6088 54916 6092 54972
rect 6092 54916 6148 54972
rect 6148 54916 6152 54972
rect 6088 54912 6152 54916
rect 9112 54972 9176 54976
rect 9112 54916 9116 54972
rect 9116 54916 9172 54972
rect 9172 54916 9176 54972
rect 9112 54912 9176 54916
rect 9192 54972 9256 54976
rect 9192 54916 9196 54972
rect 9196 54916 9252 54972
rect 9252 54916 9256 54972
rect 9192 54912 9256 54916
rect 9272 54972 9336 54976
rect 9272 54916 9276 54972
rect 9276 54916 9332 54972
rect 9332 54916 9336 54972
rect 9272 54912 9336 54916
rect 9352 54972 9416 54976
rect 9352 54916 9356 54972
rect 9356 54916 9412 54972
rect 9412 54916 9416 54972
rect 9352 54912 9416 54916
rect 1348 54844 1412 54908
rect 1900 54844 1964 54908
rect 2084 54844 2148 54908
rect 2268 54436 2332 54500
rect 3188 54436 3252 54500
rect 4216 54428 4280 54432
rect 4216 54372 4220 54428
rect 4220 54372 4276 54428
rect 4276 54372 4280 54428
rect 4216 54368 4280 54372
rect 4296 54428 4360 54432
rect 4296 54372 4300 54428
rect 4300 54372 4356 54428
rect 4356 54372 4360 54428
rect 4296 54368 4360 54372
rect 4376 54428 4440 54432
rect 4376 54372 4380 54428
rect 4380 54372 4436 54428
rect 4436 54372 4440 54428
rect 4376 54368 4440 54372
rect 4456 54428 4520 54432
rect 4456 54372 4460 54428
rect 4460 54372 4516 54428
rect 4516 54372 4520 54428
rect 4456 54368 4520 54372
rect 7480 54428 7544 54432
rect 7480 54372 7484 54428
rect 7484 54372 7540 54428
rect 7540 54372 7544 54428
rect 7480 54368 7544 54372
rect 7560 54428 7624 54432
rect 7560 54372 7564 54428
rect 7564 54372 7620 54428
rect 7620 54372 7624 54428
rect 7560 54368 7624 54372
rect 7640 54428 7704 54432
rect 7640 54372 7644 54428
rect 7644 54372 7700 54428
rect 7700 54372 7704 54428
rect 7640 54368 7704 54372
rect 7720 54428 7784 54432
rect 7720 54372 7724 54428
rect 7724 54372 7780 54428
rect 7780 54372 7784 54428
rect 7720 54368 7784 54372
rect 3924 54300 3988 54364
rect 3188 54028 3252 54092
rect 2584 53884 2648 53888
rect 2584 53828 2588 53884
rect 2588 53828 2644 53884
rect 2644 53828 2648 53884
rect 2584 53824 2648 53828
rect 2664 53884 2728 53888
rect 2664 53828 2668 53884
rect 2668 53828 2724 53884
rect 2724 53828 2728 53884
rect 2664 53824 2728 53828
rect 2744 53884 2808 53888
rect 2744 53828 2748 53884
rect 2748 53828 2804 53884
rect 2804 53828 2808 53884
rect 2744 53824 2808 53828
rect 2824 53884 2888 53888
rect 2824 53828 2828 53884
rect 2828 53828 2884 53884
rect 2884 53828 2888 53884
rect 2824 53824 2888 53828
rect 5848 53884 5912 53888
rect 5848 53828 5852 53884
rect 5852 53828 5908 53884
rect 5908 53828 5912 53884
rect 5848 53824 5912 53828
rect 5928 53884 5992 53888
rect 5928 53828 5932 53884
rect 5932 53828 5988 53884
rect 5988 53828 5992 53884
rect 5928 53824 5992 53828
rect 6008 53884 6072 53888
rect 6008 53828 6012 53884
rect 6012 53828 6068 53884
rect 6068 53828 6072 53884
rect 6008 53824 6072 53828
rect 6088 53884 6152 53888
rect 6088 53828 6092 53884
rect 6092 53828 6148 53884
rect 6148 53828 6152 53884
rect 6088 53824 6152 53828
rect 9112 53884 9176 53888
rect 9112 53828 9116 53884
rect 9116 53828 9172 53884
rect 9172 53828 9176 53884
rect 9112 53824 9176 53828
rect 9192 53884 9256 53888
rect 9192 53828 9196 53884
rect 9196 53828 9252 53884
rect 9252 53828 9256 53884
rect 9192 53824 9256 53828
rect 9272 53884 9336 53888
rect 9272 53828 9276 53884
rect 9276 53828 9332 53884
rect 9332 53828 9336 53884
rect 9272 53824 9336 53828
rect 9352 53884 9416 53888
rect 9352 53828 9356 53884
rect 9356 53828 9412 53884
rect 9412 53828 9416 53884
rect 9352 53824 9416 53828
rect 244 53484 308 53548
rect 5212 53620 5276 53684
rect 4660 53484 4724 53548
rect 4216 53340 4280 53344
rect 4216 53284 4220 53340
rect 4220 53284 4276 53340
rect 4276 53284 4280 53340
rect 4216 53280 4280 53284
rect 4296 53340 4360 53344
rect 4296 53284 4300 53340
rect 4300 53284 4356 53340
rect 4356 53284 4360 53340
rect 4296 53280 4360 53284
rect 4376 53340 4440 53344
rect 4376 53284 4380 53340
rect 4380 53284 4436 53340
rect 4436 53284 4440 53340
rect 4376 53280 4440 53284
rect 4456 53340 4520 53344
rect 4456 53284 4460 53340
rect 4460 53284 4516 53340
rect 4516 53284 4520 53340
rect 4456 53280 4520 53284
rect 7480 53340 7544 53344
rect 7480 53284 7484 53340
rect 7484 53284 7540 53340
rect 7540 53284 7544 53340
rect 7480 53280 7544 53284
rect 7560 53340 7624 53344
rect 7560 53284 7564 53340
rect 7564 53284 7620 53340
rect 7620 53284 7624 53340
rect 7560 53280 7624 53284
rect 7640 53340 7704 53344
rect 7640 53284 7644 53340
rect 7644 53284 7700 53340
rect 7700 53284 7704 53340
rect 7640 53280 7704 53284
rect 7720 53340 7784 53344
rect 7720 53284 7724 53340
rect 7724 53284 7780 53340
rect 7780 53284 7784 53340
rect 7720 53280 7784 53284
rect 2084 53076 2148 53140
rect 5028 53136 5092 53140
rect 5028 53080 5078 53136
rect 5078 53080 5092 53136
rect 5028 53076 5092 53080
rect 2584 52796 2648 52800
rect 2584 52740 2588 52796
rect 2588 52740 2644 52796
rect 2644 52740 2648 52796
rect 2584 52736 2648 52740
rect 2664 52796 2728 52800
rect 2664 52740 2668 52796
rect 2668 52740 2724 52796
rect 2724 52740 2728 52796
rect 2664 52736 2728 52740
rect 2744 52796 2808 52800
rect 2744 52740 2748 52796
rect 2748 52740 2804 52796
rect 2804 52740 2808 52796
rect 2744 52736 2808 52740
rect 2824 52796 2888 52800
rect 2824 52740 2828 52796
rect 2828 52740 2884 52796
rect 2884 52740 2888 52796
rect 2824 52736 2888 52740
rect 5848 52796 5912 52800
rect 5848 52740 5852 52796
rect 5852 52740 5908 52796
rect 5908 52740 5912 52796
rect 5848 52736 5912 52740
rect 5928 52796 5992 52800
rect 5928 52740 5932 52796
rect 5932 52740 5988 52796
rect 5988 52740 5992 52796
rect 5928 52736 5992 52740
rect 6008 52796 6072 52800
rect 6008 52740 6012 52796
rect 6012 52740 6068 52796
rect 6068 52740 6072 52796
rect 6008 52736 6072 52740
rect 6088 52796 6152 52800
rect 6088 52740 6092 52796
rect 6092 52740 6148 52796
rect 6148 52740 6152 52796
rect 6088 52736 6152 52740
rect 9112 52796 9176 52800
rect 9112 52740 9116 52796
rect 9116 52740 9172 52796
rect 9172 52740 9176 52796
rect 9112 52736 9176 52740
rect 9192 52796 9256 52800
rect 9192 52740 9196 52796
rect 9196 52740 9252 52796
rect 9252 52740 9256 52796
rect 9192 52736 9256 52740
rect 9272 52796 9336 52800
rect 9272 52740 9276 52796
rect 9276 52740 9332 52796
rect 9332 52740 9336 52796
rect 9272 52736 9336 52740
rect 9352 52796 9416 52800
rect 9352 52740 9356 52796
rect 9356 52740 9412 52796
rect 9412 52740 9416 52796
rect 9352 52736 9416 52740
rect 980 52532 1044 52596
rect 4216 52252 4280 52256
rect 4216 52196 4220 52252
rect 4220 52196 4276 52252
rect 4276 52196 4280 52252
rect 4216 52192 4280 52196
rect 4296 52252 4360 52256
rect 4296 52196 4300 52252
rect 4300 52196 4356 52252
rect 4356 52196 4360 52252
rect 4296 52192 4360 52196
rect 4376 52252 4440 52256
rect 4376 52196 4380 52252
rect 4380 52196 4436 52252
rect 4436 52196 4440 52252
rect 4376 52192 4440 52196
rect 4456 52252 4520 52256
rect 4456 52196 4460 52252
rect 4460 52196 4516 52252
rect 4516 52196 4520 52252
rect 4456 52192 4520 52196
rect 7480 52252 7544 52256
rect 7480 52196 7484 52252
rect 7484 52196 7540 52252
rect 7540 52196 7544 52252
rect 7480 52192 7544 52196
rect 7560 52252 7624 52256
rect 7560 52196 7564 52252
rect 7564 52196 7620 52252
rect 7620 52196 7624 52252
rect 7560 52192 7624 52196
rect 7640 52252 7704 52256
rect 7640 52196 7644 52252
rect 7644 52196 7700 52252
rect 7700 52196 7704 52252
rect 7640 52192 7704 52196
rect 7720 52252 7784 52256
rect 7720 52196 7724 52252
rect 7724 52196 7780 52252
rect 7780 52196 7784 52252
rect 7720 52192 7784 52196
rect 2268 52124 2332 52188
rect 2084 51988 2148 52052
rect 2084 51852 2148 51916
rect 2584 51708 2648 51712
rect 2584 51652 2588 51708
rect 2588 51652 2644 51708
rect 2644 51652 2648 51708
rect 2584 51648 2648 51652
rect 2664 51708 2728 51712
rect 2664 51652 2668 51708
rect 2668 51652 2724 51708
rect 2724 51652 2728 51708
rect 2664 51648 2728 51652
rect 2744 51708 2808 51712
rect 2744 51652 2748 51708
rect 2748 51652 2804 51708
rect 2804 51652 2808 51708
rect 2744 51648 2808 51652
rect 2824 51708 2888 51712
rect 2824 51652 2828 51708
rect 2828 51652 2884 51708
rect 2884 51652 2888 51708
rect 2824 51648 2888 51652
rect 5848 51708 5912 51712
rect 5848 51652 5852 51708
rect 5852 51652 5908 51708
rect 5908 51652 5912 51708
rect 5848 51648 5912 51652
rect 5928 51708 5992 51712
rect 5928 51652 5932 51708
rect 5932 51652 5988 51708
rect 5988 51652 5992 51708
rect 5928 51648 5992 51652
rect 6008 51708 6072 51712
rect 6008 51652 6012 51708
rect 6012 51652 6068 51708
rect 6068 51652 6072 51708
rect 6008 51648 6072 51652
rect 6088 51708 6152 51712
rect 6088 51652 6092 51708
rect 6092 51652 6148 51708
rect 6148 51652 6152 51708
rect 6088 51648 6152 51652
rect 9112 51708 9176 51712
rect 9112 51652 9116 51708
rect 9116 51652 9172 51708
rect 9172 51652 9176 51708
rect 9112 51648 9176 51652
rect 9192 51708 9256 51712
rect 9192 51652 9196 51708
rect 9196 51652 9252 51708
rect 9252 51652 9256 51708
rect 9192 51648 9256 51652
rect 9272 51708 9336 51712
rect 9272 51652 9276 51708
rect 9276 51652 9332 51708
rect 9332 51652 9336 51708
rect 9272 51648 9336 51652
rect 9352 51708 9416 51712
rect 9352 51652 9356 51708
rect 9356 51652 9412 51708
rect 9412 51652 9416 51708
rect 9352 51648 9416 51652
rect 1164 51444 1228 51508
rect 3004 51504 3068 51508
rect 3004 51448 3054 51504
rect 3054 51448 3068 51504
rect 3004 51444 3068 51448
rect 1900 51308 1964 51372
rect 1900 51232 1964 51236
rect 1900 51176 1950 51232
rect 1950 51176 1964 51232
rect 1900 51172 1964 51176
rect 612 50934 676 50998
rect 2268 50900 2332 50964
rect 4844 51172 4908 51236
rect 4216 51164 4280 51168
rect 4216 51108 4220 51164
rect 4220 51108 4276 51164
rect 4276 51108 4280 51164
rect 4216 51104 4280 51108
rect 4296 51164 4360 51168
rect 4296 51108 4300 51164
rect 4300 51108 4356 51164
rect 4356 51108 4360 51164
rect 4296 51104 4360 51108
rect 4376 51164 4440 51168
rect 4376 51108 4380 51164
rect 4380 51108 4436 51164
rect 4436 51108 4440 51164
rect 4376 51104 4440 51108
rect 4456 51164 4520 51168
rect 4456 51108 4460 51164
rect 4460 51108 4516 51164
rect 4516 51108 4520 51164
rect 4456 51104 4520 51108
rect 7480 51164 7544 51168
rect 7480 51108 7484 51164
rect 7484 51108 7540 51164
rect 7540 51108 7544 51164
rect 7480 51104 7544 51108
rect 7560 51164 7624 51168
rect 7560 51108 7564 51164
rect 7564 51108 7620 51164
rect 7620 51108 7624 51164
rect 7560 51104 7624 51108
rect 7640 51164 7704 51168
rect 7640 51108 7644 51164
rect 7644 51108 7700 51164
rect 7700 51108 7704 51164
rect 7640 51104 7704 51108
rect 7720 51164 7784 51168
rect 7720 51108 7724 51164
rect 7724 51108 7780 51164
rect 7780 51108 7784 51164
rect 7720 51104 7784 51108
rect 5028 51096 5092 51100
rect 5028 51040 5078 51096
rect 5078 51040 5092 51096
rect 5028 51036 5092 51040
rect 4844 50900 4908 50964
rect 4660 50764 4724 50828
rect 2584 50620 2648 50624
rect 2584 50564 2588 50620
rect 2588 50564 2644 50620
rect 2644 50564 2648 50620
rect 2584 50560 2648 50564
rect 2664 50620 2728 50624
rect 2664 50564 2668 50620
rect 2668 50564 2724 50620
rect 2724 50564 2728 50620
rect 2664 50560 2728 50564
rect 2744 50620 2808 50624
rect 2744 50564 2748 50620
rect 2748 50564 2804 50620
rect 2804 50564 2808 50620
rect 2744 50560 2808 50564
rect 2824 50620 2888 50624
rect 2824 50564 2828 50620
rect 2828 50564 2884 50620
rect 2884 50564 2888 50620
rect 2824 50560 2888 50564
rect 5848 50620 5912 50624
rect 5848 50564 5852 50620
rect 5852 50564 5908 50620
rect 5908 50564 5912 50620
rect 5848 50560 5912 50564
rect 5928 50620 5992 50624
rect 5928 50564 5932 50620
rect 5932 50564 5988 50620
rect 5988 50564 5992 50620
rect 5928 50560 5992 50564
rect 6008 50620 6072 50624
rect 6008 50564 6012 50620
rect 6012 50564 6068 50620
rect 6068 50564 6072 50620
rect 6008 50560 6072 50564
rect 6088 50620 6152 50624
rect 6088 50564 6092 50620
rect 6092 50564 6148 50620
rect 6148 50564 6152 50620
rect 6088 50560 6152 50564
rect 9112 50620 9176 50624
rect 9112 50564 9116 50620
rect 9116 50564 9172 50620
rect 9172 50564 9176 50620
rect 9112 50560 9176 50564
rect 9192 50620 9256 50624
rect 9192 50564 9196 50620
rect 9196 50564 9252 50620
rect 9252 50564 9256 50620
rect 9192 50560 9256 50564
rect 9272 50620 9336 50624
rect 9272 50564 9276 50620
rect 9276 50564 9332 50620
rect 9332 50564 9336 50620
rect 9272 50560 9336 50564
rect 9352 50620 9416 50624
rect 9352 50564 9356 50620
rect 9356 50564 9412 50620
rect 9412 50564 9416 50620
rect 9352 50560 9416 50564
rect 1532 50356 1596 50420
rect 3740 50356 3804 50420
rect 5212 50220 5276 50284
rect 428 50084 492 50148
rect 1532 50084 1596 50148
rect 4216 50076 4280 50080
rect 4216 50020 4220 50076
rect 4220 50020 4276 50076
rect 4276 50020 4280 50076
rect 4216 50016 4280 50020
rect 4296 50076 4360 50080
rect 4296 50020 4300 50076
rect 4300 50020 4356 50076
rect 4356 50020 4360 50076
rect 4296 50016 4360 50020
rect 4376 50076 4440 50080
rect 4376 50020 4380 50076
rect 4380 50020 4436 50076
rect 4436 50020 4440 50076
rect 4376 50016 4440 50020
rect 4456 50076 4520 50080
rect 4456 50020 4460 50076
rect 4460 50020 4516 50076
rect 4516 50020 4520 50076
rect 4456 50016 4520 50020
rect 7480 50076 7544 50080
rect 7480 50020 7484 50076
rect 7484 50020 7540 50076
rect 7540 50020 7544 50076
rect 7480 50016 7544 50020
rect 7560 50076 7624 50080
rect 7560 50020 7564 50076
rect 7564 50020 7620 50076
rect 7620 50020 7624 50076
rect 7560 50016 7624 50020
rect 7640 50076 7704 50080
rect 7640 50020 7644 50076
rect 7644 50020 7700 50076
rect 7700 50020 7704 50076
rect 7640 50016 7704 50020
rect 7720 50076 7784 50080
rect 7720 50020 7724 50076
rect 7724 50020 7780 50076
rect 7780 50020 7784 50076
rect 7720 50016 7784 50020
rect 2268 50008 2332 50012
rect 2268 49952 2318 50008
rect 2318 49952 2332 50008
rect 2268 49948 2332 49952
rect 1164 49676 1228 49740
rect 1716 49600 1780 49604
rect 1716 49544 1730 49600
rect 1730 49544 1780 49600
rect 1716 49540 1780 49544
rect 2584 49532 2648 49536
rect 2584 49476 2588 49532
rect 2588 49476 2644 49532
rect 2644 49476 2648 49532
rect 2584 49472 2648 49476
rect 2664 49532 2728 49536
rect 2664 49476 2668 49532
rect 2668 49476 2724 49532
rect 2724 49476 2728 49532
rect 2664 49472 2728 49476
rect 2744 49532 2808 49536
rect 2744 49476 2748 49532
rect 2748 49476 2804 49532
rect 2804 49476 2808 49532
rect 2744 49472 2808 49476
rect 2824 49532 2888 49536
rect 2824 49476 2828 49532
rect 2828 49476 2884 49532
rect 2884 49476 2888 49532
rect 2824 49472 2888 49476
rect 5848 49532 5912 49536
rect 5848 49476 5852 49532
rect 5852 49476 5908 49532
rect 5908 49476 5912 49532
rect 5848 49472 5912 49476
rect 5928 49532 5992 49536
rect 5928 49476 5932 49532
rect 5932 49476 5988 49532
rect 5988 49476 5992 49532
rect 5928 49472 5992 49476
rect 6008 49532 6072 49536
rect 6008 49476 6012 49532
rect 6012 49476 6068 49532
rect 6068 49476 6072 49532
rect 6008 49472 6072 49476
rect 6088 49532 6152 49536
rect 6088 49476 6092 49532
rect 6092 49476 6148 49532
rect 6148 49476 6152 49532
rect 6088 49472 6152 49476
rect 9112 49532 9176 49536
rect 9112 49476 9116 49532
rect 9116 49476 9172 49532
rect 9172 49476 9176 49532
rect 9112 49472 9176 49476
rect 9192 49532 9256 49536
rect 9192 49476 9196 49532
rect 9196 49476 9252 49532
rect 9252 49476 9256 49532
rect 9192 49472 9256 49476
rect 9272 49532 9336 49536
rect 9272 49476 9276 49532
rect 9276 49476 9332 49532
rect 9332 49476 9336 49532
rect 9272 49472 9336 49476
rect 9352 49532 9416 49536
rect 9352 49476 9356 49532
rect 9356 49476 9412 49532
rect 9412 49476 9416 49532
rect 9352 49472 9416 49476
rect 4660 49404 4724 49468
rect 3924 49268 3988 49332
rect 1716 49132 1780 49196
rect 3556 49132 3620 49196
rect 3924 49192 3988 49196
rect 3924 49136 3974 49192
rect 3974 49136 3988 49192
rect 3924 49132 3988 49136
rect 5212 49132 5276 49196
rect 4216 48988 4280 48992
rect 4216 48932 4220 48988
rect 4220 48932 4276 48988
rect 4276 48932 4280 48988
rect 4216 48928 4280 48932
rect 4296 48988 4360 48992
rect 4296 48932 4300 48988
rect 4300 48932 4356 48988
rect 4356 48932 4360 48988
rect 4296 48928 4360 48932
rect 4376 48988 4440 48992
rect 4376 48932 4380 48988
rect 4380 48932 4436 48988
rect 4436 48932 4440 48988
rect 4376 48928 4440 48932
rect 4456 48988 4520 48992
rect 4456 48932 4460 48988
rect 4460 48932 4516 48988
rect 4516 48932 4520 48988
rect 4456 48928 4520 48932
rect 7480 48988 7544 48992
rect 7480 48932 7484 48988
rect 7484 48932 7540 48988
rect 7540 48932 7544 48988
rect 7480 48928 7544 48932
rect 7560 48988 7624 48992
rect 7560 48932 7564 48988
rect 7564 48932 7620 48988
rect 7620 48932 7624 48988
rect 7560 48928 7624 48932
rect 7640 48988 7704 48992
rect 7640 48932 7644 48988
rect 7644 48932 7700 48988
rect 7700 48932 7704 48988
rect 7640 48928 7704 48932
rect 7720 48988 7784 48992
rect 7720 48932 7724 48988
rect 7724 48932 7780 48988
rect 7780 48932 7784 48988
rect 7720 48928 7784 48932
rect 1532 48452 1596 48516
rect 1900 48452 1964 48516
rect 2584 48444 2648 48448
rect 2584 48388 2588 48444
rect 2588 48388 2644 48444
rect 2644 48388 2648 48444
rect 2584 48384 2648 48388
rect 2664 48444 2728 48448
rect 2664 48388 2668 48444
rect 2668 48388 2724 48444
rect 2724 48388 2728 48444
rect 2664 48384 2728 48388
rect 2744 48444 2808 48448
rect 2744 48388 2748 48444
rect 2748 48388 2804 48444
rect 2804 48388 2808 48444
rect 2744 48384 2808 48388
rect 2824 48444 2888 48448
rect 2824 48388 2828 48444
rect 2828 48388 2884 48444
rect 2884 48388 2888 48444
rect 2824 48384 2888 48388
rect 3556 48588 3620 48652
rect 5848 48444 5912 48448
rect 5848 48388 5852 48444
rect 5852 48388 5908 48444
rect 5908 48388 5912 48444
rect 5848 48384 5912 48388
rect 5928 48444 5992 48448
rect 5928 48388 5932 48444
rect 5932 48388 5988 48444
rect 5988 48388 5992 48444
rect 5928 48384 5992 48388
rect 6008 48444 6072 48448
rect 6008 48388 6012 48444
rect 6012 48388 6068 48444
rect 6068 48388 6072 48444
rect 6008 48384 6072 48388
rect 6088 48444 6152 48448
rect 6088 48388 6092 48444
rect 6092 48388 6148 48444
rect 6148 48388 6152 48444
rect 6088 48384 6152 48388
rect 9112 48444 9176 48448
rect 9112 48388 9116 48444
rect 9116 48388 9172 48444
rect 9172 48388 9176 48444
rect 9112 48384 9176 48388
rect 9192 48444 9256 48448
rect 9192 48388 9196 48444
rect 9196 48388 9252 48444
rect 9252 48388 9256 48444
rect 9192 48384 9256 48388
rect 9272 48444 9336 48448
rect 9272 48388 9276 48444
rect 9276 48388 9332 48444
rect 9332 48388 9336 48444
rect 9272 48384 9336 48388
rect 9352 48444 9416 48448
rect 9352 48388 9356 48444
rect 9356 48388 9412 48444
rect 9412 48388 9416 48444
rect 9352 48384 9416 48388
rect 4660 48316 4724 48380
rect 1348 48044 1412 48108
rect 1900 48044 1964 48108
rect 5396 48044 5460 48108
rect 1532 47908 1596 47972
rect 4216 47900 4280 47904
rect 4216 47844 4220 47900
rect 4220 47844 4276 47900
rect 4276 47844 4280 47900
rect 4216 47840 4280 47844
rect 4296 47900 4360 47904
rect 4296 47844 4300 47900
rect 4300 47844 4356 47900
rect 4356 47844 4360 47900
rect 4296 47840 4360 47844
rect 4376 47900 4440 47904
rect 4376 47844 4380 47900
rect 4380 47844 4436 47900
rect 4436 47844 4440 47900
rect 4376 47840 4440 47844
rect 4456 47900 4520 47904
rect 4456 47844 4460 47900
rect 4460 47844 4516 47900
rect 4516 47844 4520 47900
rect 4456 47840 4520 47844
rect 7480 47900 7544 47904
rect 7480 47844 7484 47900
rect 7484 47844 7540 47900
rect 7540 47844 7544 47900
rect 7480 47840 7544 47844
rect 7560 47900 7624 47904
rect 7560 47844 7564 47900
rect 7564 47844 7620 47900
rect 7620 47844 7624 47900
rect 7560 47840 7624 47844
rect 7640 47900 7704 47904
rect 7640 47844 7644 47900
rect 7644 47844 7700 47900
rect 7700 47844 7704 47900
rect 7640 47840 7704 47844
rect 7720 47900 7784 47904
rect 7720 47844 7724 47900
rect 7724 47844 7780 47900
rect 7780 47844 7784 47900
rect 7720 47840 7784 47844
rect 5396 47500 5460 47564
rect 2584 47356 2648 47360
rect 2584 47300 2588 47356
rect 2588 47300 2644 47356
rect 2644 47300 2648 47356
rect 2584 47296 2648 47300
rect 2664 47356 2728 47360
rect 2664 47300 2668 47356
rect 2668 47300 2724 47356
rect 2724 47300 2728 47356
rect 2664 47296 2728 47300
rect 2744 47356 2808 47360
rect 2744 47300 2748 47356
rect 2748 47300 2804 47356
rect 2804 47300 2808 47356
rect 2744 47296 2808 47300
rect 2824 47356 2888 47360
rect 2824 47300 2828 47356
rect 2828 47300 2884 47356
rect 2884 47300 2888 47356
rect 2824 47296 2888 47300
rect 5848 47356 5912 47360
rect 5848 47300 5852 47356
rect 5852 47300 5908 47356
rect 5908 47300 5912 47356
rect 5848 47296 5912 47300
rect 5928 47356 5992 47360
rect 5928 47300 5932 47356
rect 5932 47300 5988 47356
rect 5988 47300 5992 47356
rect 5928 47296 5992 47300
rect 6008 47356 6072 47360
rect 6008 47300 6012 47356
rect 6012 47300 6068 47356
rect 6068 47300 6072 47356
rect 6008 47296 6072 47300
rect 6088 47356 6152 47360
rect 6088 47300 6092 47356
rect 6092 47300 6148 47356
rect 6148 47300 6152 47356
rect 6088 47296 6152 47300
rect 9112 47356 9176 47360
rect 9112 47300 9116 47356
rect 9116 47300 9172 47356
rect 9172 47300 9176 47356
rect 9112 47296 9176 47300
rect 9192 47356 9256 47360
rect 9192 47300 9196 47356
rect 9196 47300 9252 47356
rect 9252 47300 9256 47356
rect 9192 47296 9256 47300
rect 9272 47356 9336 47360
rect 9272 47300 9276 47356
rect 9276 47300 9332 47356
rect 9332 47300 9336 47356
rect 9272 47296 9336 47300
rect 9352 47356 9416 47360
rect 9352 47300 9356 47356
rect 9356 47300 9412 47356
rect 9412 47300 9416 47356
rect 9352 47296 9416 47300
rect 3188 47092 3252 47156
rect 4660 46956 4724 47020
rect 3004 46820 3068 46884
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 7480 46812 7544 46816
rect 7480 46756 7484 46812
rect 7484 46756 7540 46812
rect 7540 46756 7544 46812
rect 7480 46752 7544 46756
rect 7560 46812 7624 46816
rect 7560 46756 7564 46812
rect 7564 46756 7620 46812
rect 7620 46756 7624 46812
rect 7560 46752 7624 46756
rect 7640 46812 7704 46816
rect 7640 46756 7644 46812
rect 7644 46756 7700 46812
rect 7700 46756 7704 46812
rect 7640 46752 7704 46756
rect 7720 46812 7784 46816
rect 7720 46756 7724 46812
rect 7724 46756 7780 46812
rect 7780 46756 7784 46812
rect 7720 46752 7784 46756
rect 428 46684 492 46748
rect 1532 46684 1596 46748
rect 3188 46684 3252 46748
rect 3556 46684 3620 46748
rect 3556 46548 3620 46612
rect 2584 46268 2648 46272
rect 2584 46212 2588 46268
rect 2588 46212 2644 46268
rect 2644 46212 2648 46268
rect 2584 46208 2648 46212
rect 2664 46268 2728 46272
rect 2664 46212 2668 46268
rect 2668 46212 2724 46268
rect 2724 46212 2728 46268
rect 2664 46208 2728 46212
rect 2744 46268 2808 46272
rect 2744 46212 2748 46268
rect 2748 46212 2804 46268
rect 2804 46212 2808 46268
rect 2744 46208 2808 46212
rect 2824 46268 2888 46272
rect 2824 46212 2828 46268
rect 2828 46212 2884 46268
rect 2884 46212 2888 46268
rect 2824 46208 2888 46212
rect 5028 46412 5092 46476
rect 5848 46268 5912 46272
rect 5848 46212 5852 46268
rect 5852 46212 5908 46268
rect 5908 46212 5912 46268
rect 5848 46208 5912 46212
rect 5928 46268 5992 46272
rect 5928 46212 5932 46268
rect 5932 46212 5988 46268
rect 5988 46212 5992 46268
rect 5928 46208 5992 46212
rect 6008 46268 6072 46272
rect 6008 46212 6012 46268
rect 6012 46212 6068 46268
rect 6068 46212 6072 46268
rect 6008 46208 6072 46212
rect 6088 46268 6152 46272
rect 6088 46212 6092 46268
rect 6092 46212 6148 46268
rect 6148 46212 6152 46268
rect 6088 46208 6152 46212
rect 9112 46268 9176 46272
rect 9112 46212 9116 46268
rect 9116 46212 9172 46268
rect 9172 46212 9176 46268
rect 9112 46208 9176 46212
rect 9192 46268 9256 46272
rect 9192 46212 9196 46268
rect 9196 46212 9252 46268
rect 9252 46212 9256 46268
rect 9192 46208 9256 46212
rect 9272 46268 9336 46272
rect 9272 46212 9276 46268
rect 9276 46212 9332 46268
rect 9332 46212 9336 46268
rect 9272 46208 9336 46212
rect 9352 46268 9416 46272
rect 9352 46212 9356 46268
rect 9356 46212 9412 46268
rect 9412 46212 9416 46268
rect 9352 46208 9416 46212
rect 612 45766 676 45830
rect 4844 45732 4908 45796
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 7480 45724 7544 45728
rect 7480 45668 7484 45724
rect 7484 45668 7540 45724
rect 7540 45668 7544 45724
rect 7480 45664 7544 45668
rect 7560 45724 7624 45728
rect 7560 45668 7564 45724
rect 7564 45668 7620 45724
rect 7620 45668 7624 45724
rect 7560 45664 7624 45668
rect 7640 45724 7704 45728
rect 7640 45668 7644 45724
rect 7644 45668 7700 45724
rect 7700 45668 7704 45724
rect 7640 45664 7704 45668
rect 7720 45724 7784 45728
rect 7720 45668 7724 45724
rect 7724 45668 7780 45724
rect 7780 45668 7784 45724
rect 7720 45664 7784 45668
rect 1348 45460 1412 45524
rect 1716 45460 1780 45524
rect 3004 45460 3068 45524
rect 2584 45180 2648 45184
rect 2584 45124 2588 45180
rect 2588 45124 2644 45180
rect 2644 45124 2648 45180
rect 2584 45120 2648 45124
rect 2664 45180 2728 45184
rect 2664 45124 2668 45180
rect 2668 45124 2724 45180
rect 2724 45124 2728 45180
rect 2664 45120 2728 45124
rect 2744 45180 2808 45184
rect 2744 45124 2748 45180
rect 2748 45124 2804 45180
rect 2804 45124 2808 45180
rect 2744 45120 2808 45124
rect 2824 45180 2888 45184
rect 2824 45124 2828 45180
rect 2828 45124 2884 45180
rect 2884 45124 2888 45180
rect 2824 45120 2888 45124
rect 5848 45180 5912 45184
rect 5848 45124 5852 45180
rect 5852 45124 5908 45180
rect 5908 45124 5912 45180
rect 5848 45120 5912 45124
rect 5928 45180 5992 45184
rect 5928 45124 5932 45180
rect 5932 45124 5988 45180
rect 5988 45124 5992 45180
rect 5928 45120 5992 45124
rect 6008 45180 6072 45184
rect 6008 45124 6012 45180
rect 6012 45124 6068 45180
rect 6068 45124 6072 45180
rect 6008 45120 6072 45124
rect 6088 45180 6152 45184
rect 6088 45124 6092 45180
rect 6092 45124 6148 45180
rect 6148 45124 6152 45180
rect 6088 45120 6152 45124
rect 9112 45180 9176 45184
rect 9112 45124 9116 45180
rect 9116 45124 9172 45180
rect 9172 45124 9176 45180
rect 9112 45120 9176 45124
rect 9192 45180 9256 45184
rect 9192 45124 9196 45180
rect 9196 45124 9252 45180
rect 9252 45124 9256 45180
rect 9192 45120 9256 45124
rect 9272 45180 9336 45184
rect 9272 45124 9276 45180
rect 9276 45124 9332 45180
rect 9332 45124 9336 45180
rect 9272 45120 9336 45124
rect 9352 45180 9416 45184
rect 9352 45124 9356 45180
rect 9356 45124 9412 45180
rect 9412 45124 9416 45180
rect 9352 45120 9416 45124
rect 3372 44780 3436 44844
rect 1532 44508 1596 44572
rect 3740 44916 3804 44980
rect 3740 44780 3804 44844
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 7480 44636 7544 44640
rect 7480 44580 7484 44636
rect 7484 44580 7540 44636
rect 7540 44580 7544 44636
rect 7480 44576 7544 44580
rect 7560 44636 7624 44640
rect 7560 44580 7564 44636
rect 7564 44580 7620 44636
rect 7620 44580 7624 44636
rect 7560 44576 7624 44580
rect 7640 44636 7704 44640
rect 7640 44580 7644 44636
rect 7644 44580 7700 44636
rect 7700 44580 7704 44636
rect 7640 44576 7704 44580
rect 7720 44636 7784 44640
rect 7720 44580 7724 44636
rect 7724 44580 7780 44636
rect 7780 44580 7784 44636
rect 7720 44576 7784 44580
rect 3188 44296 3252 44300
rect 3188 44240 3202 44296
rect 3202 44240 3252 44296
rect 3188 44236 3252 44240
rect 2584 44092 2648 44096
rect 2584 44036 2588 44092
rect 2588 44036 2644 44092
rect 2644 44036 2648 44092
rect 2584 44032 2648 44036
rect 2664 44092 2728 44096
rect 2664 44036 2668 44092
rect 2668 44036 2724 44092
rect 2724 44036 2728 44092
rect 2664 44032 2728 44036
rect 2744 44092 2808 44096
rect 2744 44036 2748 44092
rect 2748 44036 2804 44092
rect 2804 44036 2808 44092
rect 2744 44032 2808 44036
rect 2824 44092 2888 44096
rect 2824 44036 2828 44092
rect 2828 44036 2884 44092
rect 2884 44036 2888 44092
rect 2824 44032 2888 44036
rect 5848 44092 5912 44096
rect 5848 44036 5852 44092
rect 5852 44036 5908 44092
rect 5908 44036 5912 44092
rect 5848 44032 5912 44036
rect 5928 44092 5992 44096
rect 5928 44036 5932 44092
rect 5932 44036 5988 44092
rect 5988 44036 5992 44092
rect 5928 44032 5992 44036
rect 6008 44092 6072 44096
rect 6008 44036 6012 44092
rect 6012 44036 6068 44092
rect 6068 44036 6072 44092
rect 6008 44032 6072 44036
rect 6088 44092 6152 44096
rect 6088 44036 6092 44092
rect 6092 44036 6148 44092
rect 6148 44036 6152 44092
rect 6088 44032 6152 44036
rect 9112 44092 9176 44096
rect 9112 44036 9116 44092
rect 9116 44036 9172 44092
rect 9172 44036 9176 44092
rect 9112 44032 9176 44036
rect 9192 44092 9256 44096
rect 9192 44036 9196 44092
rect 9196 44036 9252 44092
rect 9252 44036 9256 44092
rect 9192 44032 9256 44036
rect 9272 44092 9336 44096
rect 9272 44036 9276 44092
rect 9276 44036 9332 44092
rect 9332 44036 9336 44092
rect 9272 44032 9336 44036
rect 9352 44092 9416 44096
rect 9352 44036 9356 44092
rect 9356 44036 9412 44092
rect 9412 44036 9416 44092
rect 9352 44032 9416 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 7480 43548 7544 43552
rect 7480 43492 7484 43548
rect 7484 43492 7540 43548
rect 7540 43492 7544 43548
rect 7480 43488 7544 43492
rect 7560 43548 7624 43552
rect 7560 43492 7564 43548
rect 7564 43492 7620 43548
rect 7620 43492 7624 43548
rect 7560 43488 7624 43492
rect 7640 43548 7704 43552
rect 7640 43492 7644 43548
rect 7644 43492 7700 43548
rect 7700 43492 7704 43548
rect 7640 43488 7704 43492
rect 7720 43548 7784 43552
rect 7720 43492 7724 43548
rect 7724 43492 7780 43548
rect 7780 43492 7784 43548
rect 7720 43488 7784 43492
rect 1716 43420 1780 43484
rect 796 43284 860 43348
rect 3372 43012 3436 43076
rect 2584 43004 2648 43008
rect 2584 42948 2588 43004
rect 2588 42948 2644 43004
rect 2644 42948 2648 43004
rect 2584 42944 2648 42948
rect 2664 43004 2728 43008
rect 2664 42948 2668 43004
rect 2668 42948 2724 43004
rect 2724 42948 2728 43004
rect 2664 42944 2728 42948
rect 2744 43004 2808 43008
rect 2744 42948 2748 43004
rect 2748 42948 2804 43004
rect 2804 42948 2808 43004
rect 2744 42944 2808 42948
rect 2824 43004 2888 43008
rect 2824 42948 2828 43004
rect 2828 42948 2884 43004
rect 2884 42948 2888 43004
rect 2824 42944 2888 42948
rect 5848 43004 5912 43008
rect 5848 42948 5852 43004
rect 5852 42948 5908 43004
rect 5908 42948 5912 43004
rect 5848 42944 5912 42948
rect 5928 43004 5992 43008
rect 5928 42948 5932 43004
rect 5932 42948 5988 43004
rect 5988 42948 5992 43004
rect 5928 42944 5992 42948
rect 6008 43004 6072 43008
rect 6008 42948 6012 43004
rect 6012 42948 6068 43004
rect 6068 42948 6072 43004
rect 6008 42944 6072 42948
rect 6088 43004 6152 43008
rect 6088 42948 6092 43004
rect 6092 42948 6148 43004
rect 6148 42948 6152 43004
rect 6088 42944 6152 42948
rect 9112 43004 9176 43008
rect 9112 42948 9116 43004
rect 9116 42948 9172 43004
rect 9172 42948 9176 43004
rect 9112 42944 9176 42948
rect 9192 43004 9256 43008
rect 9192 42948 9196 43004
rect 9196 42948 9252 43004
rect 9252 42948 9256 43004
rect 9192 42944 9256 42948
rect 9272 43004 9336 43008
rect 9272 42948 9276 43004
rect 9276 42948 9332 43004
rect 9332 42948 9336 43004
rect 9272 42944 9336 42948
rect 9352 43004 9416 43008
rect 9352 42948 9356 43004
rect 9356 42948 9412 43004
rect 9412 42948 9416 43004
rect 9352 42944 9416 42948
rect 3372 42740 3436 42804
rect 4660 42740 4724 42804
rect 1900 42468 1964 42532
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 7480 42460 7544 42464
rect 7480 42404 7484 42460
rect 7484 42404 7540 42460
rect 7540 42404 7544 42460
rect 7480 42400 7544 42404
rect 7560 42460 7624 42464
rect 7560 42404 7564 42460
rect 7564 42404 7620 42460
rect 7620 42404 7624 42460
rect 7560 42400 7624 42404
rect 7640 42460 7704 42464
rect 7640 42404 7644 42460
rect 7644 42404 7700 42460
rect 7700 42404 7704 42460
rect 7640 42400 7704 42404
rect 7720 42460 7784 42464
rect 7720 42404 7724 42460
rect 7724 42404 7780 42460
rect 7780 42404 7784 42460
rect 7720 42400 7784 42404
rect 2268 42332 2332 42396
rect 3556 42196 3620 42260
rect 1900 42060 1964 42124
rect 5212 42060 5276 42124
rect 5212 41924 5276 41988
rect 2584 41916 2648 41920
rect 2584 41860 2588 41916
rect 2588 41860 2644 41916
rect 2644 41860 2648 41916
rect 2584 41856 2648 41860
rect 2664 41916 2728 41920
rect 2664 41860 2668 41916
rect 2668 41860 2724 41916
rect 2724 41860 2728 41916
rect 2664 41856 2728 41860
rect 2744 41916 2808 41920
rect 2744 41860 2748 41916
rect 2748 41860 2804 41916
rect 2804 41860 2808 41916
rect 2744 41856 2808 41860
rect 2824 41916 2888 41920
rect 2824 41860 2828 41916
rect 2828 41860 2884 41916
rect 2884 41860 2888 41916
rect 2824 41856 2888 41860
rect 5848 41916 5912 41920
rect 5848 41860 5852 41916
rect 5852 41860 5908 41916
rect 5908 41860 5912 41916
rect 5848 41856 5912 41860
rect 5928 41916 5992 41920
rect 5928 41860 5932 41916
rect 5932 41860 5988 41916
rect 5988 41860 5992 41916
rect 5928 41856 5992 41860
rect 6008 41916 6072 41920
rect 6008 41860 6012 41916
rect 6012 41860 6068 41916
rect 6068 41860 6072 41916
rect 6008 41856 6072 41860
rect 6088 41916 6152 41920
rect 6088 41860 6092 41916
rect 6092 41860 6148 41916
rect 6148 41860 6152 41916
rect 6088 41856 6152 41860
rect 9112 41916 9176 41920
rect 9112 41860 9116 41916
rect 9116 41860 9172 41916
rect 9172 41860 9176 41916
rect 9112 41856 9176 41860
rect 9192 41916 9256 41920
rect 9192 41860 9196 41916
rect 9196 41860 9252 41916
rect 9252 41860 9256 41916
rect 9192 41856 9256 41860
rect 9272 41916 9336 41920
rect 9272 41860 9276 41916
rect 9276 41860 9332 41916
rect 9332 41860 9336 41916
rect 9272 41856 9336 41860
rect 9352 41916 9416 41920
rect 9352 41860 9356 41916
rect 9356 41860 9412 41916
rect 9412 41860 9416 41916
rect 9352 41856 9416 41860
rect 3004 41516 3068 41580
rect 1900 41108 1964 41172
rect 3004 41032 3068 41036
rect 4660 41516 4724 41580
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 7480 41372 7544 41376
rect 7480 41316 7484 41372
rect 7484 41316 7540 41372
rect 7540 41316 7544 41372
rect 7480 41312 7544 41316
rect 7560 41372 7624 41376
rect 7560 41316 7564 41372
rect 7564 41316 7620 41372
rect 7620 41316 7624 41372
rect 7560 41312 7624 41316
rect 7640 41372 7704 41376
rect 7640 41316 7644 41372
rect 7644 41316 7700 41372
rect 7700 41316 7704 41372
rect 7640 41312 7704 41316
rect 7720 41372 7784 41376
rect 7720 41316 7724 41372
rect 7724 41316 7780 41372
rect 7780 41316 7784 41372
rect 7720 41312 7784 41316
rect 3004 40976 3054 41032
rect 3054 40976 3068 41032
rect 3004 40972 3068 40976
rect 1532 40836 1596 40900
rect 2584 40828 2648 40832
rect 2584 40772 2588 40828
rect 2588 40772 2644 40828
rect 2644 40772 2648 40828
rect 2584 40768 2648 40772
rect 2664 40828 2728 40832
rect 2664 40772 2668 40828
rect 2668 40772 2724 40828
rect 2724 40772 2728 40828
rect 2664 40768 2728 40772
rect 2744 40828 2808 40832
rect 2744 40772 2748 40828
rect 2748 40772 2804 40828
rect 2804 40772 2808 40828
rect 2744 40768 2808 40772
rect 2824 40828 2888 40832
rect 2824 40772 2828 40828
rect 2828 40772 2884 40828
rect 2884 40772 2888 40828
rect 2824 40768 2888 40772
rect 5848 40828 5912 40832
rect 5848 40772 5852 40828
rect 5852 40772 5908 40828
rect 5908 40772 5912 40828
rect 5848 40768 5912 40772
rect 5928 40828 5992 40832
rect 5928 40772 5932 40828
rect 5932 40772 5988 40828
rect 5988 40772 5992 40828
rect 5928 40768 5992 40772
rect 6008 40828 6072 40832
rect 6008 40772 6012 40828
rect 6012 40772 6068 40828
rect 6068 40772 6072 40828
rect 6008 40768 6072 40772
rect 6088 40828 6152 40832
rect 6088 40772 6092 40828
rect 6092 40772 6148 40828
rect 6148 40772 6152 40828
rect 6088 40768 6152 40772
rect 9112 40828 9176 40832
rect 9112 40772 9116 40828
rect 9116 40772 9172 40828
rect 9172 40772 9176 40828
rect 9112 40768 9176 40772
rect 9192 40828 9256 40832
rect 9192 40772 9196 40828
rect 9196 40772 9252 40828
rect 9252 40772 9256 40828
rect 9192 40768 9256 40772
rect 9272 40828 9336 40832
rect 9272 40772 9276 40828
rect 9276 40772 9332 40828
rect 9332 40772 9336 40828
rect 9272 40768 9336 40772
rect 9352 40828 9416 40832
rect 9352 40772 9356 40828
rect 9356 40772 9412 40828
rect 9412 40772 9416 40828
rect 9352 40768 9416 40772
rect 1716 40760 1780 40764
rect 1716 40704 1766 40760
rect 1766 40704 1780 40760
rect 1716 40700 1780 40704
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 7480 40284 7544 40288
rect 7480 40228 7484 40284
rect 7484 40228 7540 40284
rect 7540 40228 7544 40284
rect 7480 40224 7544 40228
rect 7560 40284 7624 40288
rect 7560 40228 7564 40284
rect 7564 40228 7620 40284
rect 7620 40228 7624 40284
rect 7560 40224 7624 40228
rect 7640 40284 7704 40288
rect 7640 40228 7644 40284
rect 7644 40228 7700 40284
rect 7700 40228 7704 40284
rect 7640 40224 7704 40228
rect 7720 40284 7784 40288
rect 7720 40228 7724 40284
rect 7724 40228 7780 40284
rect 7780 40228 7784 40284
rect 7720 40224 7784 40228
rect 2268 40020 2332 40084
rect 3188 40020 3252 40084
rect 244 39884 308 39948
rect 428 39884 492 39948
rect 3556 39884 3620 39948
rect 2584 39740 2648 39744
rect 2584 39684 2588 39740
rect 2588 39684 2644 39740
rect 2644 39684 2648 39740
rect 2584 39680 2648 39684
rect 2664 39740 2728 39744
rect 2664 39684 2668 39740
rect 2668 39684 2724 39740
rect 2724 39684 2728 39740
rect 2664 39680 2728 39684
rect 2744 39740 2808 39744
rect 2744 39684 2748 39740
rect 2748 39684 2804 39740
rect 2804 39684 2808 39740
rect 2744 39680 2808 39684
rect 2824 39740 2888 39744
rect 2824 39684 2828 39740
rect 2828 39684 2884 39740
rect 2884 39684 2888 39740
rect 2824 39680 2888 39684
rect 5848 39740 5912 39744
rect 5848 39684 5852 39740
rect 5852 39684 5908 39740
rect 5908 39684 5912 39740
rect 5848 39680 5912 39684
rect 5928 39740 5992 39744
rect 5928 39684 5932 39740
rect 5932 39684 5988 39740
rect 5988 39684 5992 39740
rect 5928 39680 5992 39684
rect 6008 39740 6072 39744
rect 6008 39684 6012 39740
rect 6012 39684 6068 39740
rect 6068 39684 6072 39740
rect 6008 39680 6072 39684
rect 6088 39740 6152 39744
rect 6088 39684 6092 39740
rect 6092 39684 6148 39740
rect 6148 39684 6152 39740
rect 6088 39680 6152 39684
rect 9112 39740 9176 39744
rect 9112 39684 9116 39740
rect 9116 39684 9172 39740
rect 9172 39684 9176 39740
rect 9112 39680 9176 39684
rect 9192 39740 9256 39744
rect 9192 39684 9196 39740
rect 9196 39684 9252 39740
rect 9252 39684 9256 39740
rect 9192 39680 9256 39684
rect 9272 39740 9336 39744
rect 9272 39684 9276 39740
rect 9276 39684 9332 39740
rect 9332 39684 9336 39740
rect 9272 39680 9336 39684
rect 9352 39740 9416 39744
rect 9352 39684 9356 39740
rect 9356 39684 9412 39740
rect 9412 39684 9416 39740
rect 9352 39680 9416 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 7480 39196 7544 39200
rect 7480 39140 7484 39196
rect 7484 39140 7540 39196
rect 7540 39140 7544 39196
rect 7480 39136 7544 39140
rect 7560 39196 7624 39200
rect 7560 39140 7564 39196
rect 7564 39140 7620 39196
rect 7620 39140 7624 39196
rect 7560 39136 7624 39140
rect 7640 39196 7704 39200
rect 7640 39140 7644 39196
rect 7644 39140 7700 39196
rect 7700 39140 7704 39196
rect 7640 39136 7704 39140
rect 7720 39196 7784 39200
rect 7720 39140 7724 39196
rect 7724 39140 7780 39196
rect 7780 39140 7784 39196
rect 7720 39136 7784 39140
rect 2268 39068 2332 39132
rect 3004 39068 3068 39132
rect 3188 38932 3252 38996
rect 3740 38932 3804 38996
rect 3004 38796 3068 38860
rect 5212 38796 5276 38860
rect 2584 38652 2648 38656
rect 2584 38596 2588 38652
rect 2588 38596 2644 38652
rect 2644 38596 2648 38652
rect 2584 38592 2648 38596
rect 2664 38652 2728 38656
rect 2664 38596 2668 38652
rect 2668 38596 2724 38652
rect 2724 38596 2728 38652
rect 2664 38592 2728 38596
rect 2744 38652 2808 38656
rect 2744 38596 2748 38652
rect 2748 38596 2804 38652
rect 2804 38596 2808 38652
rect 2744 38592 2808 38596
rect 2824 38652 2888 38656
rect 2824 38596 2828 38652
rect 2828 38596 2884 38652
rect 2884 38596 2888 38652
rect 2824 38592 2888 38596
rect 5848 38652 5912 38656
rect 5848 38596 5852 38652
rect 5852 38596 5908 38652
rect 5908 38596 5912 38652
rect 5848 38592 5912 38596
rect 5928 38652 5992 38656
rect 5928 38596 5932 38652
rect 5932 38596 5988 38652
rect 5988 38596 5992 38652
rect 5928 38592 5992 38596
rect 6008 38652 6072 38656
rect 6008 38596 6012 38652
rect 6012 38596 6068 38652
rect 6068 38596 6072 38652
rect 6008 38592 6072 38596
rect 6088 38652 6152 38656
rect 6088 38596 6092 38652
rect 6092 38596 6148 38652
rect 6148 38596 6152 38652
rect 6088 38592 6152 38596
rect 9112 38652 9176 38656
rect 9112 38596 9116 38652
rect 9116 38596 9172 38652
rect 9172 38596 9176 38652
rect 9112 38592 9176 38596
rect 9192 38652 9256 38656
rect 9192 38596 9196 38652
rect 9196 38596 9252 38652
rect 9252 38596 9256 38652
rect 9192 38592 9256 38596
rect 9272 38652 9336 38656
rect 9272 38596 9276 38652
rect 9276 38596 9332 38652
rect 9332 38596 9336 38652
rect 9272 38592 9336 38596
rect 9352 38652 9416 38656
rect 9352 38596 9356 38652
rect 9356 38596 9412 38652
rect 9412 38596 9416 38652
rect 9352 38592 9416 38596
rect 5212 38252 5276 38316
rect 1900 38116 1964 38180
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 7480 38108 7544 38112
rect 7480 38052 7484 38108
rect 7484 38052 7540 38108
rect 7540 38052 7544 38108
rect 7480 38048 7544 38052
rect 7560 38108 7624 38112
rect 7560 38052 7564 38108
rect 7564 38052 7620 38108
rect 7620 38052 7624 38108
rect 7560 38048 7624 38052
rect 7640 38108 7704 38112
rect 7640 38052 7644 38108
rect 7644 38052 7700 38108
rect 7700 38052 7704 38108
rect 7640 38048 7704 38052
rect 7720 38108 7784 38112
rect 7720 38052 7724 38108
rect 7724 38052 7780 38108
rect 7780 38052 7784 38108
rect 7720 38048 7784 38052
rect 3188 37844 3252 37908
rect 1532 37708 1596 37772
rect 2584 37564 2648 37568
rect 2584 37508 2588 37564
rect 2588 37508 2644 37564
rect 2644 37508 2648 37564
rect 2584 37504 2648 37508
rect 2664 37564 2728 37568
rect 2664 37508 2668 37564
rect 2668 37508 2724 37564
rect 2724 37508 2728 37564
rect 2664 37504 2728 37508
rect 2744 37564 2808 37568
rect 2744 37508 2748 37564
rect 2748 37508 2804 37564
rect 2804 37508 2808 37564
rect 2744 37504 2808 37508
rect 2824 37564 2888 37568
rect 2824 37508 2828 37564
rect 2828 37508 2884 37564
rect 2884 37508 2888 37564
rect 2824 37504 2888 37508
rect 5848 37564 5912 37568
rect 5848 37508 5852 37564
rect 5852 37508 5908 37564
rect 5908 37508 5912 37564
rect 5848 37504 5912 37508
rect 5928 37564 5992 37568
rect 5928 37508 5932 37564
rect 5932 37508 5988 37564
rect 5988 37508 5992 37564
rect 5928 37504 5992 37508
rect 6008 37564 6072 37568
rect 6008 37508 6012 37564
rect 6012 37508 6068 37564
rect 6068 37508 6072 37564
rect 6008 37504 6072 37508
rect 6088 37564 6152 37568
rect 6088 37508 6092 37564
rect 6092 37508 6148 37564
rect 6148 37508 6152 37564
rect 6088 37504 6152 37508
rect 9112 37564 9176 37568
rect 9112 37508 9116 37564
rect 9116 37508 9172 37564
rect 9172 37508 9176 37564
rect 9112 37504 9176 37508
rect 9192 37564 9256 37568
rect 9192 37508 9196 37564
rect 9196 37508 9252 37564
rect 9252 37508 9256 37564
rect 9192 37504 9256 37508
rect 9272 37564 9336 37568
rect 9272 37508 9276 37564
rect 9276 37508 9332 37564
rect 9332 37508 9336 37564
rect 9272 37504 9336 37508
rect 9352 37564 9416 37568
rect 9352 37508 9356 37564
rect 9356 37508 9412 37564
rect 9412 37508 9416 37564
rect 9352 37504 9416 37508
rect 4660 37300 4724 37364
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 7480 37020 7544 37024
rect 7480 36964 7484 37020
rect 7484 36964 7540 37020
rect 7540 36964 7544 37020
rect 7480 36960 7544 36964
rect 7560 37020 7624 37024
rect 7560 36964 7564 37020
rect 7564 36964 7620 37020
rect 7620 36964 7624 37020
rect 7560 36960 7624 36964
rect 7640 37020 7704 37024
rect 7640 36964 7644 37020
rect 7644 36964 7700 37020
rect 7700 36964 7704 37020
rect 7640 36960 7704 36964
rect 7720 37020 7784 37024
rect 7720 36964 7724 37020
rect 7724 36964 7780 37020
rect 7780 36964 7784 37020
rect 7720 36960 7784 36964
rect 4660 36756 4724 36820
rect 5396 36756 5460 36820
rect 2584 36476 2648 36480
rect 2584 36420 2588 36476
rect 2588 36420 2644 36476
rect 2644 36420 2648 36476
rect 2584 36416 2648 36420
rect 2664 36476 2728 36480
rect 2664 36420 2668 36476
rect 2668 36420 2724 36476
rect 2724 36420 2728 36476
rect 2664 36416 2728 36420
rect 2744 36476 2808 36480
rect 2744 36420 2748 36476
rect 2748 36420 2804 36476
rect 2804 36420 2808 36476
rect 2744 36416 2808 36420
rect 2824 36476 2888 36480
rect 2824 36420 2828 36476
rect 2828 36420 2884 36476
rect 2884 36420 2888 36476
rect 2824 36416 2888 36420
rect 5848 36476 5912 36480
rect 5848 36420 5852 36476
rect 5852 36420 5908 36476
rect 5908 36420 5912 36476
rect 5848 36416 5912 36420
rect 5928 36476 5992 36480
rect 5928 36420 5932 36476
rect 5932 36420 5988 36476
rect 5988 36420 5992 36476
rect 5928 36416 5992 36420
rect 6008 36476 6072 36480
rect 6008 36420 6012 36476
rect 6012 36420 6068 36476
rect 6068 36420 6072 36476
rect 6008 36416 6072 36420
rect 6088 36476 6152 36480
rect 6088 36420 6092 36476
rect 6092 36420 6148 36476
rect 6148 36420 6152 36476
rect 6088 36416 6152 36420
rect 9112 36476 9176 36480
rect 9112 36420 9116 36476
rect 9116 36420 9172 36476
rect 9172 36420 9176 36476
rect 9112 36416 9176 36420
rect 9192 36476 9256 36480
rect 9192 36420 9196 36476
rect 9196 36420 9252 36476
rect 9252 36420 9256 36476
rect 9192 36416 9256 36420
rect 9272 36476 9336 36480
rect 9272 36420 9276 36476
rect 9276 36420 9332 36476
rect 9332 36420 9336 36476
rect 9272 36416 9336 36420
rect 9352 36476 9416 36480
rect 9352 36420 9356 36476
rect 9356 36420 9412 36476
rect 9412 36420 9416 36476
rect 9352 36416 9416 36420
rect 5212 36076 5276 36140
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 7480 35932 7544 35936
rect 7480 35876 7484 35932
rect 7484 35876 7540 35932
rect 7540 35876 7544 35932
rect 7480 35872 7544 35876
rect 7560 35932 7624 35936
rect 7560 35876 7564 35932
rect 7564 35876 7620 35932
rect 7620 35876 7624 35932
rect 7560 35872 7624 35876
rect 7640 35932 7704 35936
rect 7640 35876 7644 35932
rect 7644 35876 7700 35932
rect 7700 35876 7704 35932
rect 7640 35872 7704 35876
rect 7720 35932 7784 35936
rect 7720 35876 7724 35932
rect 7724 35876 7780 35932
rect 7780 35876 7784 35932
rect 7720 35872 7784 35876
rect 2584 35388 2648 35392
rect 2584 35332 2588 35388
rect 2588 35332 2644 35388
rect 2644 35332 2648 35388
rect 2584 35328 2648 35332
rect 2664 35388 2728 35392
rect 2664 35332 2668 35388
rect 2668 35332 2724 35388
rect 2724 35332 2728 35388
rect 2664 35328 2728 35332
rect 2744 35388 2808 35392
rect 2744 35332 2748 35388
rect 2748 35332 2804 35388
rect 2804 35332 2808 35388
rect 2744 35328 2808 35332
rect 2824 35388 2888 35392
rect 2824 35332 2828 35388
rect 2828 35332 2884 35388
rect 2884 35332 2888 35388
rect 2824 35328 2888 35332
rect 5848 35388 5912 35392
rect 5848 35332 5852 35388
rect 5852 35332 5908 35388
rect 5908 35332 5912 35388
rect 5848 35328 5912 35332
rect 5928 35388 5992 35392
rect 5928 35332 5932 35388
rect 5932 35332 5988 35388
rect 5988 35332 5992 35388
rect 5928 35328 5992 35332
rect 6008 35388 6072 35392
rect 6008 35332 6012 35388
rect 6012 35332 6068 35388
rect 6068 35332 6072 35388
rect 6008 35328 6072 35332
rect 6088 35388 6152 35392
rect 6088 35332 6092 35388
rect 6092 35332 6148 35388
rect 6148 35332 6152 35388
rect 6088 35328 6152 35332
rect 9112 35388 9176 35392
rect 9112 35332 9116 35388
rect 9116 35332 9172 35388
rect 9172 35332 9176 35388
rect 9112 35328 9176 35332
rect 9192 35388 9256 35392
rect 9192 35332 9196 35388
rect 9196 35332 9252 35388
rect 9252 35332 9256 35388
rect 9192 35328 9256 35332
rect 9272 35388 9336 35392
rect 9272 35332 9276 35388
rect 9276 35332 9332 35388
rect 9332 35332 9336 35388
rect 9272 35328 9336 35332
rect 9352 35388 9416 35392
rect 9352 35332 9356 35388
rect 9356 35332 9412 35388
rect 9412 35332 9416 35388
rect 9352 35328 9416 35332
rect 1716 34912 1780 34916
rect 1716 34856 1730 34912
rect 1730 34856 1780 34912
rect 1716 34852 1780 34856
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 7480 34844 7544 34848
rect 7480 34788 7484 34844
rect 7484 34788 7540 34844
rect 7540 34788 7544 34844
rect 7480 34784 7544 34788
rect 7560 34844 7624 34848
rect 7560 34788 7564 34844
rect 7564 34788 7620 34844
rect 7620 34788 7624 34844
rect 7560 34784 7624 34788
rect 7640 34844 7704 34848
rect 7640 34788 7644 34844
rect 7644 34788 7700 34844
rect 7700 34788 7704 34844
rect 7640 34784 7704 34788
rect 7720 34844 7784 34848
rect 7720 34788 7724 34844
rect 7724 34788 7780 34844
rect 7780 34788 7784 34844
rect 7720 34784 7784 34788
rect 2584 34300 2648 34304
rect 2584 34244 2588 34300
rect 2588 34244 2644 34300
rect 2644 34244 2648 34300
rect 2584 34240 2648 34244
rect 2664 34300 2728 34304
rect 2664 34244 2668 34300
rect 2668 34244 2724 34300
rect 2724 34244 2728 34300
rect 2664 34240 2728 34244
rect 2744 34300 2808 34304
rect 2744 34244 2748 34300
rect 2748 34244 2804 34300
rect 2804 34244 2808 34300
rect 2744 34240 2808 34244
rect 2824 34300 2888 34304
rect 2824 34244 2828 34300
rect 2828 34244 2884 34300
rect 2884 34244 2888 34300
rect 2824 34240 2888 34244
rect 5848 34300 5912 34304
rect 5848 34244 5852 34300
rect 5852 34244 5908 34300
rect 5908 34244 5912 34300
rect 5848 34240 5912 34244
rect 5928 34300 5992 34304
rect 5928 34244 5932 34300
rect 5932 34244 5988 34300
rect 5988 34244 5992 34300
rect 5928 34240 5992 34244
rect 6008 34300 6072 34304
rect 6008 34244 6012 34300
rect 6012 34244 6068 34300
rect 6068 34244 6072 34300
rect 6008 34240 6072 34244
rect 6088 34300 6152 34304
rect 6088 34244 6092 34300
rect 6092 34244 6148 34300
rect 6148 34244 6152 34300
rect 6088 34240 6152 34244
rect 9112 34300 9176 34304
rect 9112 34244 9116 34300
rect 9116 34244 9172 34300
rect 9172 34244 9176 34300
rect 9112 34240 9176 34244
rect 9192 34300 9256 34304
rect 9192 34244 9196 34300
rect 9196 34244 9252 34300
rect 9252 34244 9256 34300
rect 9192 34240 9256 34244
rect 9272 34300 9336 34304
rect 9272 34244 9276 34300
rect 9276 34244 9332 34300
rect 9332 34244 9336 34300
rect 9272 34240 9336 34244
rect 9352 34300 9416 34304
rect 9352 34244 9356 34300
rect 9356 34244 9412 34300
rect 9412 34244 9416 34300
rect 9352 34240 9416 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 7480 33756 7544 33760
rect 7480 33700 7484 33756
rect 7484 33700 7540 33756
rect 7540 33700 7544 33756
rect 7480 33696 7544 33700
rect 7560 33756 7624 33760
rect 7560 33700 7564 33756
rect 7564 33700 7620 33756
rect 7620 33700 7624 33756
rect 7560 33696 7624 33700
rect 7640 33756 7704 33760
rect 7640 33700 7644 33756
rect 7644 33700 7700 33756
rect 7700 33700 7704 33756
rect 7640 33696 7704 33700
rect 7720 33756 7784 33760
rect 7720 33700 7724 33756
rect 7724 33700 7780 33756
rect 7780 33700 7784 33756
rect 7720 33696 7784 33700
rect 2584 33212 2648 33216
rect 2584 33156 2588 33212
rect 2588 33156 2644 33212
rect 2644 33156 2648 33212
rect 2584 33152 2648 33156
rect 2664 33212 2728 33216
rect 2664 33156 2668 33212
rect 2668 33156 2724 33212
rect 2724 33156 2728 33212
rect 2664 33152 2728 33156
rect 2744 33212 2808 33216
rect 2744 33156 2748 33212
rect 2748 33156 2804 33212
rect 2804 33156 2808 33212
rect 2744 33152 2808 33156
rect 2824 33212 2888 33216
rect 2824 33156 2828 33212
rect 2828 33156 2884 33212
rect 2884 33156 2888 33212
rect 2824 33152 2888 33156
rect 5848 33212 5912 33216
rect 5848 33156 5852 33212
rect 5852 33156 5908 33212
rect 5908 33156 5912 33212
rect 5848 33152 5912 33156
rect 5928 33212 5992 33216
rect 5928 33156 5932 33212
rect 5932 33156 5988 33212
rect 5988 33156 5992 33212
rect 5928 33152 5992 33156
rect 6008 33212 6072 33216
rect 6008 33156 6012 33212
rect 6012 33156 6068 33212
rect 6068 33156 6072 33212
rect 6008 33152 6072 33156
rect 6088 33212 6152 33216
rect 6088 33156 6092 33212
rect 6092 33156 6148 33212
rect 6148 33156 6152 33212
rect 6088 33152 6152 33156
rect 9112 33212 9176 33216
rect 9112 33156 9116 33212
rect 9116 33156 9172 33212
rect 9172 33156 9176 33212
rect 9112 33152 9176 33156
rect 9192 33212 9256 33216
rect 9192 33156 9196 33212
rect 9196 33156 9252 33212
rect 9252 33156 9256 33212
rect 9192 33152 9256 33156
rect 9272 33212 9336 33216
rect 9272 33156 9276 33212
rect 9276 33156 9332 33212
rect 9332 33156 9336 33212
rect 9272 33152 9336 33156
rect 9352 33212 9416 33216
rect 9352 33156 9356 33212
rect 9356 33156 9412 33212
rect 9412 33156 9416 33212
rect 9352 33152 9416 33156
rect 3556 32948 3620 33012
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 7480 32668 7544 32672
rect 7480 32612 7484 32668
rect 7484 32612 7540 32668
rect 7540 32612 7544 32668
rect 7480 32608 7544 32612
rect 7560 32668 7624 32672
rect 7560 32612 7564 32668
rect 7564 32612 7620 32668
rect 7620 32612 7624 32668
rect 7560 32608 7624 32612
rect 7640 32668 7704 32672
rect 7640 32612 7644 32668
rect 7644 32612 7700 32668
rect 7700 32612 7704 32668
rect 7640 32608 7704 32612
rect 7720 32668 7784 32672
rect 7720 32612 7724 32668
rect 7724 32612 7780 32668
rect 7780 32612 7784 32668
rect 7720 32608 7784 32612
rect 5212 32404 5276 32468
rect 1900 32192 1964 32196
rect 1900 32136 1950 32192
rect 1950 32136 1964 32192
rect 1900 32132 1964 32136
rect 3188 32132 3252 32196
rect 2584 32124 2648 32128
rect 2584 32068 2588 32124
rect 2588 32068 2644 32124
rect 2644 32068 2648 32124
rect 2584 32064 2648 32068
rect 2664 32124 2728 32128
rect 2664 32068 2668 32124
rect 2668 32068 2724 32124
rect 2724 32068 2728 32124
rect 2664 32064 2728 32068
rect 2744 32124 2808 32128
rect 2744 32068 2748 32124
rect 2748 32068 2804 32124
rect 2804 32068 2808 32124
rect 2744 32064 2808 32068
rect 2824 32124 2888 32128
rect 2824 32068 2828 32124
rect 2828 32068 2884 32124
rect 2884 32068 2888 32124
rect 2824 32064 2888 32068
rect 3188 31996 3252 32060
rect 3740 32132 3804 32196
rect 3740 31996 3804 32060
rect 5848 32124 5912 32128
rect 5848 32068 5852 32124
rect 5852 32068 5908 32124
rect 5908 32068 5912 32124
rect 5848 32064 5912 32068
rect 5928 32124 5992 32128
rect 5928 32068 5932 32124
rect 5932 32068 5988 32124
rect 5988 32068 5992 32124
rect 5928 32064 5992 32068
rect 6008 32124 6072 32128
rect 6008 32068 6012 32124
rect 6012 32068 6068 32124
rect 6068 32068 6072 32124
rect 6008 32064 6072 32068
rect 6088 32124 6152 32128
rect 6088 32068 6092 32124
rect 6092 32068 6148 32124
rect 6148 32068 6152 32124
rect 6088 32064 6152 32068
rect 9112 32124 9176 32128
rect 9112 32068 9116 32124
rect 9116 32068 9172 32124
rect 9172 32068 9176 32124
rect 9112 32064 9176 32068
rect 9192 32124 9256 32128
rect 9192 32068 9196 32124
rect 9196 32068 9252 32124
rect 9252 32068 9256 32124
rect 9192 32064 9256 32068
rect 9272 32124 9336 32128
rect 9272 32068 9276 32124
rect 9276 32068 9332 32124
rect 9332 32068 9336 32124
rect 9272 32064 9336 32068
rect 9352 32124 9416 32128
rect 9352 32068 9356 32124
rect 9356 32068 9412 32124
rect 9412 32068 9416 32124
rect 9352 32064 9416 32068
rect 5212 31996 5276 32060
rect 5396 31724 5460 31788
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 3004 31452 3068 31516
rect 3740 31452 3804 31516
rect 1900 31316 1964 31380
rect 3004 31316 3068 31380
rect 7480 31580 7544 31584
rect 7480 31524 7484 31580
rect 7484 31524 7540 31580
rect 7540 31524 7544 31580
rect 7480 31520 7544 31524
rect 7560 31580 7624 31584
rect 7560 31524 7564 31580
rect 7564 31524 7620 31580
rect 7620 31524 7624 31580
rect 7560 31520 7624 31524
rect 7640 31580 7704 31584
rect 7640 31524 7644 31580
rect 7644 31524 7700 31580
rect 7700 31524 7704 31580
rect 7640 31520 7704 31524
rect 7720 31580 7784 31584
rect 7720 31524 7724 31580
rect 7724 31524 7780 31580
rect 7780 31524 7784 31580
rect 7720 31520 7784 31524
rect 980 31044 1044 31108
rect 2584 31036 2648 31040
rect 2584 30980 2588 31036
rect 2588 30980 2644 31036
rect 2644 30980 2648 31036
rect 2584 30976 2648 30980
rect 2664 31036 2728 31040
rect 2664 30980 2668 31036
rect 2668 30980 2724 31036
rect 2724 30980 2728 31036
rect 2664 30976 2728 30980
rect 2744 31036 2808 31040
rect 2744 30980 2748 31036
rect 2748 30980 2804 31036
rect 2804 30980 2808 31036
rect 2744 30976 2808 30980
rect 2824 31036 2888 31040
rect 2824 30980 2828 31036
rect 2828 30980 2884 31036
rect 2884 30980 2888 31036
rect 2824 30976 2888 30980
rect 5848 31036 5912 31040
rect 5848 30980 5852 31036
rect 5852 30980 5908 31036
rect 5908 30980 5912 31036
rect 5848 30976 5912 30980
rect 5928 31036 5992 31040
rect 5928 30980 5932 31036
rect 5932 30980 5988 31036
rect 5988 30980 5992 31036
rect 5928 30976 5992 30980
rect 6008 31036 6072 31040
rect 6008 30980 6012 31036
rect 6012 30980 6068 31036
rect 6068 30980 6072 31036
rect 6008 30976 6072 30980
rect 6088 31036 6152 31040
rect 6088 30980 6092 31036
rect 6092 30980 6148 31036
rect 6148 30980 6152 31036
rect 6088 30976 6152 30980
rect 9112 31036 9176 31040
rect 9112 30980 9116 31036
rect 9116 30980 9172 31036
rect 9172 30980 9176 31036
rect 9112 30976 9176 30980
rect 9192 31036 9256 31040
rect 9192 30980 9196 31036
rect 9196 30980 9252 31036
rect 9252 30980 9256 31036
rect 9192 30976 9256 30980
rect 9272 31036 9336 31040
rect 9272 30980 9276 31036
rect 9276 30980 9332 31036
rect 9332 30980 9336 31036
rect 9272 30976 9336 30980
rect 9352 31036 9416 31040
rect 9352 30980 9356 31036
rect 9356 30980 9412 31036
rect 9412 30980 9416 31036
rect 9352 30976 9416 30980
rect 3740 30908 3804 30972
rect 1532 30636 1596 30700
rect 1348 30500 1412 30564
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 7480 30492 7544 30496
rect 7480 30436 7484 30492
rect 7484 30436 7540 30492
rect 7540 30436 7544 30492
rect 7480 30432 7544 30436
rect 7560 30492 7624 30496
rect 7560 30436 7564 30492
rect 7564 30436 7620 30492
rect 7620 30436 7624 30492
rect 7560 30432 7624 30436
rect 7640 30492 7704 30496
rect 7640 30436 7644 30492
rect 7644 30436 7700 30492
rect 7700 30436 7704 30492
rect 7640 30432 7704 30436
rect 7720 30492 7784 30496
rect 7720 30436 7724 30492
rect 7724 30436 7780 30492
rect 7780 30436 7784 30492
rect 7720 30432 7784 30436
rect 3372 30364 3436 30428
rect 1164 30228 1228 30292
rect 1532 29956 1596 30020
rect 2584 29948 2648 29952
rect 2584 29892 2588 29948
rect 2588 29892 2644 29948
rect 2644 29892 2648 29948
rect 2584 29888 2648 29892
rect 2664 29948 2728 29952
rect 2664 29892 2668 29948
rect 2668 29892 2724 29948
rect 2724 29892 2728 29948
rect 2664 29888 2728 29892
rect 2744 29948 2808 29952
rect 2744 29892 2748 29948
rect 2748 29892 2804 29948
rect 2804 29892 2808 29948
rect 2744 29888 2808 29892
rect 2824 29948 2888 29952
rect 2824 29892 2828 29948
rect 2828 29892 2884 29948
rect 2884 29892 2888 29948
rect 2824 29888 2888 29892
rect 5848 29948 5912 29952
rect 5848 29892 5852 29948
rect 5852 29892 5908 29948
rect 5908 29892 5912 29948
rect 5848 29888 5912 29892
rect 5928 29948 5992 29952
rect 5928 29892 5932 29948
rect 5932 29892 5988 29948
rect 5988 29892 5992 29948
rect 5928 29888 5992 29892
rect 6008 29948 6072 29952
rect 6008 29892 6012 29948
rect 6012 29892 6068 29948
rect 6068 29892 6072 29948
rect 6008 29888 6072 29892
rect 6088 29948 6152 29952
rect 6088 29892 6092 29948
rect 6092 29892 6148 29948
rect 6148 29892 6152 29948
rect 6088 29888 6152 29892
rect 9112 29948 9176 29952
rect 9112 29892 9116 29948
rect 9116 29892 9172 29948
rect 9172 29892 9176 29948
rect 9112 29888 9176 29892
rect 9192 29948 9256 29952
rect 9192 29892 9196 29948
rect 9196 29892 9252 29948
rect 9252 29892 9256 29948
rect 9192 29888 9256 29892
rect 9272 29948 9336 29952
rect 9272 29892 9276 29948
rect 9276 29892 9332 29948
rect 9332 29892 9336 29948
rect 9272 29888 9336 29892
rect 9352 29948 9416 29952
rect 9352 29892 9356 29948
rect 9356 29892 9412 29948
rect 9412 29892 9416 29948
rect 9352 29888 9416 29892
rect 2084 29880 2148 29884
rect 2084 29824 2098 29880
rect 2098 29824 2148 29880
rect 2084 29820 2148 29824
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 7480 29404 7544 29408
rect 7480 29348 7484 29404
rect 7484 29348 7540 29404
rect 7540 29348 7544 29404
rect 7480 29344 7544 29348
rect 7560 29404 7624 29408
rect 7560 29348 7564 29404
rect 7564 29348 7620 29404
rect 7620 29348 7624 29404
rect 7560 29344 7624 29348
rect 7640 29404 7704 29408
rect 7640 29348 7644 29404
rect 7644 29348 7700 29404
rect 7700 29348 7704 29404
rect 7640 29344 7704 29348
rect 7720 29404 7784 29408
rect 7720 29348 7724 29404
rect 7724 29348 7780 29404
rect 7780 29348 7784 29404
rect 7720 29344 7784 29348
rect 2268 29276 2332 29340
rect 1900 28928 1964 28932
rect 1900 28872 1950 28928
rect 1950 28872 1964 28928
rect 1900 28868 1964 28872
rect 2084 28928 2148 28932
rect 2084 28872 2134 28928
rect 2134 28872 2148 28928
rect 2084 28868 2148 28872
rect 2268 28460 2332 28524
rect 2584 28860 2648 28864
rect 2584 28804 2588 28860
rect 2588 28804 2644 28860
rect 2644 28804 2648 28860
rect 2584 28800 2648 28804
rect 2664 28860 2728 28864
rect 2664 28804 2668 28860
rect 2668 28804 2724 28860
rect 2724 28804 2728 28860
rect 2664 28800 2728 28804
rect 2744 28860 2808 28864
rect 2744 28804 2748 28860
rect 2748 28804 2804 28860
rect 2804 28804 2808 28860
rect 2744 28800 2808 28804
rect 2824 28860 2888 28864
rect 2824 28804 2828 28860
rect 2828 28804 2884 28860
rect 2884 28804 2888 28860
rect 2824 28800 2888 28804
rect 5848 28860 5912 28864
rect 5848 28804 5852 28860
rect 5852 28804 5908 28860
rect 5908 28804 5912 28860
rect 5848 28800 5912 28804
rect 5928 28860 5992 28864
rect 5928 28804 5932 28860
rect 5932 28804 5988 28860
rect 5988 28804 5992 28860
rect 5928 28800 5992 28804
rect 6008 28860 6072 28864
rect 6008 28804 6012 28860
rect 6012 28804 6068 28860
rect 6068 28804 6072 28860
rect 6008 28800 6072 28804
rect 6088 28860 6152 28864
rect 6088 28804 6092 28860
rect 6092 28804 6148 28860
rect 6148 28804 6152 28860
rect 6088 28800 6152 28804
rect 9112 28860 9176 28864
rect 9112 28804 9116 28860
rect 9116 28804 9172 28860
rect 9172 28804 9176 28860
rect 9112 28800 9176 28804
rect 9192 28860 9256 28864
rect 9192 28804 9196 28860
rect 9196 28804 9252 28860
rect 9252 28804 9256 28860
rect 9192 28800 9256 28804
rect 9272 28860 9336 28864
rect 9272 28804 9276 28860
rect 9276 28804 9332 28860
rect 9332 28804 9336 28860
rect 9272 28800 9336 28804
rect 9352 28860 9416 28864
rect 9352 28804 9356 28860
rect 9356 28804 9412 28860
rect 9412 28804 9416 28860
rect 9352 28800 9416 28804
rect 3004 28596 3068 28660
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 7480 28316 7544 28320
rect 7480 28260 7484 28316
rect 7484 28260 7540 28316
rect 7540 28260 7544 28316
rect 7480 28256 7544 28260
rect 7560 28316 7624 28320
rect 7560 28260 7564 28316
rect 7564 28260 7620 28316
rect 7620 28260 7624 28316
rect 7560 28256 7624 28260
rect 7640 28316 7704 28320
rect 7640 28260 7644 28316
rect 7644 28260 7700 28316
rect 7700 28260 7704 28316
rect 7640 28256 7704 28260
rect 7720 28316 7784 28320
rect 7720 28260 7724 28316
rect 7724 28260 7780 28316
rect 7780 28260 7784 28316
rect 7720 28256 7784 28260
rect 1900 28188 1964 28252
rect 1532 28112 1596 28116
rect 1532 28056 1546 28112
rect 1546 28056 1596 28112
rect 1532 28052 1596 28056
rect 5580 28052 5644 28116
rect 2084 27916 2148 27980
rect 3556 27916 3620 27980
rect 2584 27772 2648 27776
rect 2584 27716 2588 27772
rect 2588 27716 2644 27772
rect 2644 27716 2648 27772
rect 2584 27712 2648 27716
rect 2664 27772 2728 27776
rect 2664 27716 2668 27772
rect 2668 27716 2724 27772
rect 2724 27716 2728 27772
rect 2664 27712 2728 27716
rect 2744 27772 2808 27776
rect 2744 27716 2748 27772
rect 2748 27716 2804 27772
rect 2804 27716 2808 27772
rect 2744 27712 2808 27716
rect 2824 27772 2888 27776
rect 2824 27716 2828 27772
rect 2828 27716 2884 27772
rect 2884 27716 2888 27772
rect 2824 27712 2888 27716
rect 5848 27772 5912 27776
rect 5848 27716 5852 27772
rect 5852 27716 5908 27772
rect 5908 27716 5912 27772
rect 5848 27712 5912 27716
rect 5928 27772 5992 27776
rect 5928 27716 5932 27772
rect 5932 27716 5988 27772
rect 5988 27716 5992 27772
rect 5928 27712 5992 27716
rect 6008 27772 6072 27776
rect 6008 27716 6012 27772
rect 6012 27716 6068 27772
rect 6068 27716 6072 27772
rect 6008 27712 6072 27716
rect 6088 27772 6152 27776
rect 6088 27716 6092 27772
rect 6092 27716 6148 27772
rect 6148 27716 6152 27772
rect 6088 27712 6152 27716
rect 9112 27772 9176 27776
rect 9112 27716 9116 27772
rect 9116 27716 9172 27772
rect 9172 27716 9176 27772
rect 9112 27712 9176 27716
rect 9192 27772 9256 27776
rect 9192 27716 9196 27772
rect 9196 27716 9252 27772
rect 9252 27716 9256 27772
rect 9192 27712 9256 27716
rect 9272 27772 9336 27776
rect 9272 27716 9276 27772
rect 9276 27716 9332 27772
rect 9332 27716 9336 27772
rect 9272 27712 9336 27716
rect 9352 27772 9416 27776
rect 9352 27716 9356 27772
rect 9356 27716 9412 27772
rect 9412 27716 9416 27772
rect 9352 27712 9416 27716
rect 3740 27372 3804 27436
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 7480 27228 7544 27232
rect 7480 27172 7484 27228
rect 7484 27172 7540 27228
rect 7540 27172 7544 27228
rect 7480 27168 7544 27172
rect 7560 27228 7624 27232
rect 7560 27172 7564 27228
rect 7564 27172 7620 27228
rect 7620 27172 7624 27228
rect 7560 27168 7624 27172
rect 7640 27228 7704 27232
rect 7640 27172 7644 27228
rect 7644 27172 7700 27228
rect 7700 27172 7704 27228
rect 7640 27168 7704 27172
rect 7720 27228 7784 27232
rect 7720 27172 7724 27228
rect 7724 27172 7780 27228
rect 7780 27172 7784 27228
rect 7720 27168 7784 27172
rect 5212 26964 5276 27028
rect 6316 26828 6380 26892
rect 2584 26684 2648 26688
rect 2584 26628 2588 26684
rect 2588 26628 2644 26684
rect 2644 26628 2648 26684
rect 2584 26624 2648 26628
rect 2664 26684 2728 26688
rect 2664 26628 2668 26684
rect 2668 26628 2724 26684
rect 2724 26628 2728 26684
rect 2664 26624 2728 26628
rect 2744 26684 2808 26688
rect 2744 26628 2748 26684
rect 2748 26628 2804 26684
rect 2804 26628 2808 26684
rect 2744 26624 2808 26628
rect 2824 26684 2888 26688
rect 2824 26628 2828 26684
rect 2828 26628 2884 26684
rect 2884 26628 2888 26684
rect 2824 26624 2888 26628
rect 5848 26684 5912 26688
rect 5848 26628 5852 26684
rect 5852 26628 5908 26684
rect 5908 26628 5912 26684
rect 5848 26624 5912 26628
rect 5928 26684 5992 26688
rect 5928 26628 5932 26684
rect 5932 26628 5988 26684
rect 5988 26628 5992 26684
rect 5928 26624 5992 26628
rect 6008 26684 6072 26688
rect 6008 26628 6012 26684
rect 6012 26628 6068 26684
rect 6068 26628 6072 26684
rect 6008 26624 6072 26628
rect 6088 26684 6152 26688
rect 6088 26628 6092 26684
rect 6092 26628 6148 26684
rect 6148 26628 6152 26684
rect 6088 26624 6152 26628
rect 9112 26684 9176 26688
rect 9112 26628 9116 26684
rect 9116 26628 9172 26684
rect 9172 26628 9176 26684
rect 9112 26624 9176 26628
rect 9192 26684 9256 26688
rect 9192 26628 9196 26684
rect 9196 26628 9252 26684
rect 9252 26628 9256 26684
rect 9192 26624 9256 26628
rect 9272 26684 9336 26688
rect 9272 26628 9276 26684
rect 9276 26628 9332 26684
rect 9332 26628 9336 26684
rect 9272 26624 9336 26628
rect 9352 26684 9416 26688
rect 9352 26628 9356 26684
rect 9356 26628 9412 26684
rect 9412 26628 9416 26684
rect 9352 26624 9416 26628
rect 3188 26344 3252 26348
rect 3188 26288 3202 26344
rect 3202 26288 3252 26344
rect 3188 26284 3252 26288
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 7480 26140 7544 26144
rect 7480 26084 7484 26140
rect 7484 26084 7540 26140
rect 7540 26084 7544 26140
rect 7480 26080 7544 26084
rect 7560 26140 7624 26144
rect 7560 26084 7564 26140
rect 7564 26084 7620 26140
rect 7620 26084 7624 26140
rect 7560 26080 7624 26084
rect 7640 26140 7704 26144
rect 7640 26084 7644 26140
rect 7644 26084 7700 26140
rect 7700 26084 7704 26140
rect 7640 26080 7704 26084
rect 7720 26140 7784 26144
rect 7720 26084 7724 26140
rect 7724 26084 7780 26140
rect 7780 26084 7784 26140
rect 7720 26080 7784 26084
rect 3556 25800 3620 25804
rect 3556 25744 3606 25800
rect 3606 25744 3620 25800
rect 3556 25740 3620 25744
rect 2584 25596 2648 25600
rect 2584 25540 2588 25596
rect 2588 25540 2644 25596
rect 2644 25540 2648 25596
rect 2584 25536 2648 25540
rect 2664 25596 2728 25600
rect 2664 25540 2668 25596
rect 2668 25540 2724 25596
rect 2724 25540 2728 25596
rect 2664 25536 2728 25540
rect 2744 25596 2808 25600
rect 2744 25540 2748 25596
rect 2748 25540 2804 25596
rect 2804 25540 2808 25596
rect 2744 25536 2808 25540
rect 2824 25596 2888 25600
rect 2824 25540 2828 25596
rect 2828 25540 2884 25596
rect 2884 25540 2888 25596
rect 2824 25536 2888 25540
rect 5848 25596 5912 25600
rect 5848 25540 5852 25596
rect 5852 25540 5908 25596
rect 5908 25540 5912 25596
rect 5848 25536 5912 25540
rect 5928 25596 5992 25600
rect 5928 25540 5932 25596
rect 5932 25540 5988 25596
rect 5988 25540 5992 25596
rect 5928 25536 5992 25540
rect 6008 25596 6072 25600
rect 6008 25540 6012 25596
rect 6012 25540 6068 25596
rect 6068 25540 6072 25596
rect 6008 25536 6072 25540
rect 6088 25596 6152 25600
rect 6088 25540 6092 25596
rect 6092 25540 6148 25596
rect 6148 25540 6152 25596
rect 6088 25536 6152 25540
rect 9112 25596 9176 25600
rect 9112 25540 9116 25596
rect 9116 25540 9172 25596
rect 9172 25540 9176 25596
rect 9112 25536 9176 25540
rect 9192 25596 9256 25600
rect 9192 25540 9196 25596
rect 9196 25540 9252 25596
rect 9252 25540 9256 25596
rect 9192 25536 9256 25540
rect 9272 25596 9336 25600
rect 9272 25540 9276 25596
rect 9276 25540 9332 25596
rect 9332 25540 9336 25596
rect 9272 25536 9336 25540
rect 9352 25596 9416 25600
rect 9352 25540 9356 25596
rect 9356 25540 9412 25596
rect 9412 25540 9416 25596
rect 9352 25536 9416 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 7480 25052 7544 25056
rect 7480 24996 7484 25052
rect 7484 24996 7540 25052
rect 7540 24996 7544 25052
rect 7480 24992 7544 24996
rect 7560 25052 7624 25056
rect 7560 24996 7564 25052
rect 7564 24996 7620 25052
rect 7620 24996 7624 25052
rect 7560 24992 7624 24996
rect 7640 25052 7704 25056
rect 7640 24996 7644 25052
rect 7644 24996 7700 25052
rect 7700 24996 7704 25052
rect 7640 24992 7704 24996
rect 7720 25052 7784 25056
rect 7720 24996 7724 25052
rect 7724 24996 7780 25052
rect 7780 24996 7784 25052
rect 7720 24992 7784 24996
rect 2584 24508 2648 24512
rect 2584 24452 2588 24508
rect 2588 24452 2644 24508
rect 2644 24452 2648 24508
rect 2584 24448 2648 24452
rect 2664 24508 2728 24512
rect 2664 24452 2668 24508
rect 2668 24452 2724 24508
rect 2724 24452 2728 24508
rect 2664 24448 2728 24452
rect 2744 24508 2808 24512
rect 2744 24452 2748 24508
rect 2748 24452 2804 24508
rect 2804 24452 2808 24508
rect 2744 24448 2808 24452
rect 2824 24508 2888 24512
rect 2824 24452 2828 24508
rect 2828 24452 2884 24508
rect 2884 24452 2888 24508
rect 2824 24448 2888 24452
rect 5848 24508 5912 24512
rect 5848 24452 5852 24508
rect 5852 24452 5908 24508
rect 5908 24452 5912 24508
rect 5848 24448 5912 24452
rect 5928 24508 5992 24512
rect 5928 24452 5932 24508
rect 5932 24452 5988 24508
rect 5988 24452 5992 24508
rect 5928 24448 5992 24452
rect 6008 24508 6072 24512
rect 6008 24452 6012 24508
rect 6012 24452 6068 24508
rect 6068 24452 6072 24508
rect 6008 24448 6072 24452
rect 6088 24508 6152 24512
rect 6088 24452 6092 24508
rect 6092 24452 6148 24508
rect 6148 24452 6152 24508
rect 6088 24448 6152 24452
rect 9112 24508 9176 24512
rect 9112 24452 9116 24508
rect 9116 24452 9172 24508
rect 9172 24452 9176 24508
rect 9112 24448 9176 24452
rect 9192 24508 9256 24512
rect 9192 24452 9196 24508
rect 9196 24452 9252 24508
rect 9252 24452 9256 24508
rect 9192 24448 9256 24452
rect 9272 24508 9336 24512
rect 9272 24452 9276 24508
rect 9276 24452 9332 24508
rect 9332 24452 9336 24508
rect 9272 24448 9336 24452
rect 9352 24508 9416 24512
rect 9352 24452 9356 24508
rect 9356 24452 9412 24508
rect 9412 24452 9416 24508
rect 9352 24448 9416 24452
rect 2268 24108 2332 24172
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 7480 23964 7544 23968
rect 7480 23908 7484 23964
rect 7484 23908 7540 23964
rect 7540 23908 7544 23964
rect 7480 23904 7544 23908
rect 7560 23964 7624 23968
rect 7560 23908 7564 23964
rect 7564 23908 7620 23964
rect 7620 23908 7624 23964
rect 7560 23904 7624 23908
rect 7640 23964 7704 23968
rect 7640 23908 7644 23964
rect 7644 23908 7700 23964
rect 7700 23908 7704 23964
rect 7640 23904 7704 23908
rect 7720 23964 7784 23968
rect 7720 23908 7724 23964
rect 7724 23908 7780 23964
rect 7780 23908 7784 23964
rect 7720 23904 7784 23908
rect 2584 23420 2648 23424
rect 2584 23364 2588 23420
rect 2588 23364 2644 23420
rect 2644 23364 2648 23420
rect 2584 23360 2648 23364
rect 2664 23420 2728 23424
rect 2664 23364 2668 23420
rect 2668 23364 2724 23420
rect 2724 23364 2728 23420
rect 2664 23360 2728 23364
rect 2744 23420 2808 23424
rect 2744 23364 2748 23420
rect 2748 23364 2804 23420
rect 2804 23364 2808 23420
rect 2744 23360 2808 23364
rect 2824 23420 2888 23424
rect 2824 23364 2828 23420
rect 2828 23364 2884 23420
rect 2884 23364 2888 23420
rect 2824 23360 2888 23364
rect 5848 23420 5912 23424
rect 5848 23364 5852 23420
rect 5852 23364 5908 23420
rect 5908 23364 5912 23420
rect 5848 23360 5912 23364
rect 5928 23420 5992 23424
rect 5928 23364 5932 23420
rect 5932 23364 5988 23420
rect 5988 23364 5992 23420
rect 5928 23360 5992 23364
rect 6008 23420 6072 23424
rect 6008 23364 6012 23420
rect 6012 23364 6068 23420
rect 6068 23364 6072 23420
rect 6008 23360 6072 23364
rect 6088 23420 6152 23424
rect 6088 23364 6092 23420
rect 6092 23364 6148 23420
rect 6148 23364 6152 23420
rect 6088 23360 6152 23364
rect 9112 23420 9176 23424
rect 9112 23364 9116 23420
rect 9116 23364 9172 23420
rect 9172 23364 9176 23420
rect 9112 23360 9176 23364
rect 9192 23420 9256 23424
rect 9192 23364 9196 23420
rect 9196 23364 9252 23420
rect 9252 23364 9256 23420
rect 9192 23360 9256 23364
rect 9272 23420 9336 23424
rect 9272 23364 9276 23420
rect 9276 23364 9332 23420
rect 9332 23364 9336 23420
rect 9272 23360 9336 23364
rect 9352 23420 9416 23424
rect 9352 23364 9356 23420
rect 9356 23364 9412 23420
rect 9412 23364 9416 23420
rect 9352 23360 9416 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 7480 22876 7544 22880
rect 7480 22820 7484 22876
rect 7484 22820 7540 22876
rect 7540 22820 7544 22876
rect 7480 22816 7544 22820
rect 7560 22876 7624 22880
rect 7560 22820 7564 22876
rect 7564 22820 7620 22876
rect 7620 22820 7624 22876
rect 7560 22816 7624 22820
rect 7640 22876 7704 22880
rect 7640 22820 7644 22876
rect 7644 22820 7700 22876
rect 7700 22820 7704 22876
rect 7640 22816 7704 22820
rect 7720 22876 7784 22880
rect 7720 22820 7724 22876
rect 7724 22820 7780 22876
rect 7780 22820 7784 22876
rect 7720 22816 7784 22820
rect 2584 22332 2648 22336
rect 2584 22276 2588 22332
rect 2588 22276 2644 22332
rect 2644 22276 2648 22332
rect 2584 22272 2648 22276
rect 2664 22332 2728 22336
rect 2664 22276 2668 22332
rect 2668 22276 2724 22332
rect 2724 22276 2728 22332
rect 2664 22272 2728 22276
rect 2744 22332 2808 22336
rect 2744 22276 2748 22332
rect 2748 22276 2804 22332
rect 2804 22276 2808 22332
rect 2744 22272 2808 22276
rect 2824 22332 2888 22336
rect 2824 22276 2828 22332
rect 2828 22276 2884 22332
rect 2884 22276 2888 22332
rect 2824 22272 2888 22276
rect 5848 22332 5912 22336
rect 5848 22276 5852 22332
rect 5852 22276 5908 22332
rect 5908 22276 5912 22332
rect 5848 22272 5912 22276
rect 5928 22332 5992 22336
rect 5928 22276 5932 22332
rect 5932 22276 5988 22332
rect 5988 22276 5992 22332
rect 5928 22272 5992 22276
rect 6008 22332 6072 22336
rect 6008 22276 6012 22332
rect 6012 22276 6068 22332
rect 6068 22276 6072 22332
rect 6008 22272 6072 22276
rect 6088 22332 6152 22336
rect 6088 22276 6092 22332
rect 6092 22276 6148 22332
rect 6148 22276 6152 22332
rect 6088 22272 6152 22276
rect 9112 22332 9176 22336
rect 9112 22276 9116 22332
rect 9116 22276 9172 22332
rect 9172 22276 9176 22332
rect 9112 22272 9176 22276
rect 9192 22332 9256 22336
rect 9192 22276 9196 22332
rect 9196 22276 9252 22332
rect 9252 22276 9256 22332
rect 9192 22272 9256 22276
rect 9272 22332 9336 22336
rect 9272 22276 9276 22332
rect 9276 22276 9332 22332
rect 9332 22276 9336 22332
rect 9272 22272 9336 22276
rect 9352 22332 9416 22336
rect 9352 22276 9356 22332
rect 9356 22276 9412 22332
rect 9412 22276 9416 22332
rect 9352 22272 9416 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 7480 21788 7544 21792
rect 7480 21732 7484 21788
rect 7484 21732 7540 21788
rect 7540 21732 7544 21788
rect 7480 21728 7544 21732
rect 7560 21788 7624 21792
rect 7560 21732 7564 21788
rect 7564 21732 7620 21788
rect 7620 21732 7624 21788
rect 7560 21728 7624 21732
rect 7640 21788 7704 21792
rect 7640 21732 7644 21788
rect 7644 21732 7700 21788
rect 7700 21732 7704 21788
rect 7640 21728 7704 21732
rect 7720 21788 7784 21792
rect 7720 21732 7724 21788
rect 7724 21732 7780 21788
rect 7780 21732 7784 21788
rect 7720 21728 7784 21732
rect 2584 21244 2648 21248
rect 2584 21188 2588 21244
rect 2588 21188 2644 21244
rect 2644 21188 2648 21244
rect 2584 21184 2648 21188
rect 2664 21244 2728 21248
rect 2664 21188 2668 21244
rect 2668 21188 2724 21244
rect 2724 21188 2728 21244
rect 2664 21184 2728 21188
rect 2744 21244 2808 21248
rect 2744 21188 2748 21244
rect 2748 21188 2804 21244
rect 2804 21188 2808 21244
rect 2744 21184 2808 21188
rect 2824 21244 2888 21248
rect 2824 21188 2828 21244
rect 2828 21188 2884 21244
rect 2884 21188 2888 21244
rect 2824 21184 2888 21188
rect 5848 21244 5912 21248
rect 5848 21188 5852 21244
rect 5852 21188 5908 21244
rect 5908 21188 5912 21244
rect 5848 21184 5912 21188
rect 5928 21244 5992 21248
rect 5928 21188 5932 21244
rect 5932 21188 5988 21244
rect 5988 21188 5992 21244
rect 5928 21184 5992 21188
rect 6008 21244 6072 21248
rect 6008 21188 6012 21244
rect 6012 21188 6068 21244
rect 6068 21188 6072 21244
rect 6008 21184 6072 21188
rect 6088 21244 6152 21248
rect 6088 21188 6092 21244
rect 6092 21188 6148 21244
rect 6148 21188 6152 21244
rect 6088 21184 6152 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 9272 21244 9336 21248
rect 9272 21188 9276 21244
rect 9276 21188 9332 21244
rect 9332 21188 9336 21244
rect 9272 21184 9336 21188
rect 9352 21244 9416 21248
rect 9352 21188 9356 21244
rect 9356 21188 9412 21244
rect 9412 21188 9416 21244
rect 9352 21184 9416 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 7480 20700 7544 20704
rect 7480 20644 7484 20700
rect 7484 20644 7540 20700
rect 7540 20644 7544 20700
rect 7480 20640 7544 20644
rect 7560 20700 7624 20704
rect 7560 20644 7564 20700
rect 7564 20644 7620 20700
rect 7620 20644 7624 20700
rect 7560 20640 7624 20644
rect 7640 20700 7704 20704
rect 7640 20644 7644 20700
rect 7644 20644 7700 20700
rect 7700 20644 7704 20700
rect 7640 20640 7704 20644
rect 7720 20700 7784 20704
rect 7720 20644 7724 20700
rect 7724 20644 7780 20700
rect 7780 20644 7784 20700
rect 7720 20640 7784 20644
rect 2584 20156 2648 20160
rect 2584 20100 2588 20156
rect 2588 20100 2644 20156
rect 2644 20100 2648 20156
rect 2584 20096 2648 20100
rect 2664 20156 2728 20160
rect 2664 20100 2668 20156
rect 2668 20100 2724 20156
rect 2724 20100 2728 20156
rect 2664 20096 2728 20100
rect 2744 20156 2808 20160
rect 2744 20100 2748 20156
rect 2748 20100 2804 20156
rect 2804 20100 2808 20156
rect 2744 20096 2808 20100
rect 2824 20156 2888 20160
rect 2824 20100 2828 20156
rect 2828 20100 2884 20156
rect 2884 20100 2888 20156
rect 2824 20096 2888 20100
rect 5848 20156 5912 20160
rect 5848 20100 5852 20156
rect 5852 20100 5908 20156
rect 5908 20100 5912 20156
rect 5848 20096 5912 20100
rect 5928 20156 5992 20160
rect 5928 20100 5932 20156
rect 5932 20100 5988 20156
rect 5988 20100 5992 20156
rect 5928 20096 5992 20100
rect 6008 20156 6072 20160
rect 6008 20100 6012 20156
rect 6012 20100 6068 20156
rect 6068 20100 6072 20156
rect 6008 20096 6072 20100
rect 6088 20156 6152 20160
rect 6088 20100 6092 20156
rect 6092 20100 6148 20156
rect 6148 20100 6152 20156
rect 6088 20096 6152 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 9272 20156 9336 20160
rect 9272 20100 9276 20156
rect 9276 20100 9332 20156
rect 9332 20100 9336 20156
rect 9272 20096 9336 20100
rect 9352 20156 9416 20160
rect 9352 20100 9356 20156
rect 9356 20100 9412 20156
rect 9412 20100 9416 20156
rect 9352 20096 9416 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 7480 19612 7544 19616
rect 7480 19556 7484 19612
rect 7484 19556 7540 19612
rect 7540 19556 7544 19612
rect 7480 19552 7544 19556
rect 7560 19612 7624 19616
rect 7560 19556 7564 19612
rect 7564 19556 7620 19612
rect 7620 19556 7624 19612
rect 7560 19552 7624 19556
rect 7640 19612 7704 19616
rect 7640 19556 7644 19612
rect 7644 19556 7700 19612
rect 7700 19556 7704 19612
rect 7640 19552 7704 19556
rect 7720 19612 7784 19616
rect 7720 19556 7724 19612
rect 7724 19556 7780 19612
rect 7780 19556 7784 19612
rect 7720 19552 7784 19556
rect 2584 19068 2648 19072
rect 2584 19012 2588 19068
rect 2588 19012 2644 19068
rect 2644 19012 2648 19068
rect 2584 19008 2648 19012
rect 2664 19068 2728 19072
rect 2664 19012 2668 19068
rect 2668 19012 2724 19068
rect 2724 19012 2728 19068
rect 2664 19008 2728 19012
rect 2744 19068 2808 19072
rect 2744 19012 2748 19068
rect 2748 19012 2804 19068
rect 2804 19012 2808 19068
rect 2744 19008 2808 19012
rect 2824 19068 2888 19072
rect 2824 19012 2828 19068
rect 2828 19012 2884 19068
rect 2884 19012 2888 19068
rect 2824 19008 2888 19012
rect 5848 19068 5912 19072
rect 5848 19012 5852 19068
rect 5852 19012 5908 19068
rect 5908 19012 5912 19068
rect 5848 19008 5912 19012
rect 5928 19068 5992 19072
rect 5928 19012 5932 19068
rect 5932 19012 5988 19068
rect 5988 19012 5992 19068
rect 5928 19008 5992 19012
rect 6008 19068 6072 19072
rect 6008 19012 6012 19068
rect 6012 19012 6068 19068
rect 6068 19012 6072 19068
rect 6008 19008 6072 19012
rect 6088 19068 6152 19072
rect 6088 19012 6092 19068
rect 6092 19012 6148 19068
rect 6148 19012 6152 19068
rect 6088 19008 6152 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 9272 19068 9336 19072
rect 9272 19012 9276 19068
rect 9276 19012 9332 19068
rect 9332 19012 9336 19068
rect 9272 19008 9336 19012
rect 9352 19068 9416 19072
rect 9352 19012 9356 19068
rect 9356 19012 9412 19068
rect 9412 19012 9416 19068
rect 9352 19008 9416 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 7480 18524 7544 18528
rect 7480 18468 7484 18524
rect 7484 18468 7540 18524
rect 7540 18468 7544 18524
rect 7480 18464 7544 18468
rect 7560 18524 7624 18528
rect 7560 18468 7564 18524
rect 7564 18468 7620 18524
rect 7620 18468 7624 18524
rect 7560 18464 7624 18468
rect 7640 18524 7704 18528
rect 7640 18468 7644 18524
rect 7644 18468 7700 18524
rect 7700 18468 7704 18524
rect 7640 18464 7704 18468
rect 7720 18524 7784 18528
rect 7720 18468 7724 18524
rect 7724 18468 7780 18524
rect 7780 18468 7784 18524
rect 7720 18464 7784 18468
rect 2584 17980 2648 17984
rect 2584 17924 2588 17980
rect 2588 17924 2644 17980
rect 2644 17924 2648 17980
rect 2584 17920 2648 17924
rect 2664 17980 2728 17984
rect 2664 17924 2668 17980
rect 2668 17924 2724 17980
rect 2724 17924 2728 17980
rect 2664 17920 2728 17924
rect 2744 17980 2808 17984
rect 2744 17924 2748 17980
rect 2748 17924 2804 17980
rect 2804 17924 2808 17980
rect 2744 17920 2808 17924
rect 2824 17980 2888 17984
rect 2824 17924 2828 17980
rect 2828 17924 2884 17980
rect 2884 17924 2888 17980
rect 2824 17920 2888 17924
rect 5848 17980 5912 17984
rect 5848 17924 5852 17980
rect 5852 17924 5908 17980
rect 5908 17924 5912 17980
rect 5848 17920 5912 17924
rect 5928 17980 5992 17984
rect 5928 17924 5932 17980
rect 5932 17924 5988 17980
rect 5988 17924 5992 17980
rect 5928 17920 5992 17924
rect 6008 17980 6072 17984
rect 6008 17924 6012 17980
rect 6012 17924 6068 17980
rect 6068 17924 6072 17980
rect 6008 17920 6072 17924
rect 6088 17980 6152 17984
rect 6088 17924 6092 17980
rect 6092 17924 6148 17980
rect 6148 17924 6152 17980
rect 6088 17920 6152 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 9272 17980 9336 17984
rect 9272 17924 9276 17980
rect 9276 17924 9332 17980
rect 9332 17924 9336 17980
rect 9272 17920 9336 17924
rect 9352 17980 9416 17984
rect 9352 17924 9356 17980
rect 9356 17924 9412 17980
rect 9412 17924 9416 17980
rect 9352 17920 9416 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 7480 17436 7544 17440
rect 7480 17380 7484 17436
rect 7484 17380 7540 17436
rect 7540 17380 7544 17436
rect 7480 17376 7544 17380
rect 7560 17436 7624 17440
rect 7560 17380 7564 17436
rect 7564 17380 7620 17436
rect 7620 17380 7624 17436
rect 7560 17376 7624 17380
rect 7640 17436 7704 17440
rect 7640 17380 7644 17436
rect 7644 17380 7700 17436
rect 7700 17380 7704 17436
rect 7640 17376 7704 17380
rect 7720 17436 7784 17440
rect 7720 17380 7724 17436
rect 7724 17380 7780 17436
rect 7780 17380 7784 17436
rect 7720 17376 7784 17380
rect 3004 17036 3068 17100
rect 2584 16892 2648 16896
rect 2584 16836 2588 16892
rect 2588 16836 2644 16892
rect 2644 16836 2648 16892
rect 2584 16832 2648 16836
rect 2664 16892 2728 16896
rect 2664 16836 2668 16892
rect 2668 16836 2724 16892
rect 2724 16836 2728 16892
rect 2664 16832 2728 16836
rect 2744 16892 2808 16896
rect 2744 16836 2748 16892
rect 2748 16836 2804 16892
rect 2804 16836 2808 16892
rect 2744 16832 2808 16836
rect 2824 16892 2888 16896
rect 2824 16836 2828 16892
rect 2828 16836 2884 16892
rect 2884 16836 2888 16892
rect 2824 16832 2888 16836
rect 5848 16892 5912 16896
rect 5848 16836 5852 16892
rect 5852 16836 5908 16892
rect 5908 16836 5912 16892
rect 5848 16832 5912 16836
rect 5928 16892 5992 16896
rect 5928 16836 5932 16892
rect 5932 16836 5988 16892
rect 5988 16836 5992 16892
rect 5928 16832 5992 16836
rect 6008 16892 6072 16896
rect 6008 16836 6012 16892
rect 6012 16836 6068 16892
rect 6068 16836 6072 16892
rect 6008 16832 6072 16836
rect 6088 16892 6152 16896
rect 6088 16836 6092 16892
rect 6092 16836 6148 16892
rect 6148 16836 6152 16892
rect 6088 16832 6152 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 9272 16892 9336 16896
rect 9272 16836 9276 16892
rect 9276 16836 9332 16892
rect 9332 16836 9336 16892
rect 9272 16832 9336 16836
rect 9352 16892 9416 16896
rect 9352 16836 9356 16892
rect 9356 16836 9412 16892
rect 9412 16836 9416 16892
rect 9352 16832 9416 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 7480 16348 7544 16352
rect 7480 16292 7484 16348
rect 7484 16292 7540 16348
rect 7540 16292 7544 16348
rect 7480 16288 7544 16292
rect 7560 16348 7624 16352
rect 7560 16292 7564 16348
rect 7564 16292 7620 16348
rect 7620 16292 7624 16348
rect 7560 16288 7624 16292
rect 7640 16348 7704 16352
rect 7640 16292 7644 16348
rect 7644 16292 7700 16348
rect 7700 16292 7704 16348
rect 7640 16288 7704 16292
rect 7720 16348 7784 16352
rect 7720 16292 7724 16348
rect 7724 16292 7780 16348
rect 7780 16292 7784 16348
rect 7720 16288 7784 16292
rect 2584 15804 2648 15808
rect 2584 15748 2588 15804
rect 2588 15748 2644 15804
rect 2644 15748 2648 15804
rect 2584 15744 2648 15748
rect 2664 15804 2728 15808
rect 2664 15748 2668 15804
rect 2668 15748 2724 15804
rect 2724 15748 2728 15804
rect 2664 15744 2728 15748
rect 2744 15804 2808 15808
rect 2744 15748 2748 15804
rect 2748 15748 2804 15804
rect 2804 15748 2808 15804
rect 2744 15744 2808 15748
rect 2824 15804 2888 15808
rect 2824 15748 2828 15804
rect 2828 15748 2884 15804
rect 2884 15748 2888 15804
rect 2824 15744 2888 15748
rect 5848 15804 5912 15808
rect 5848 15748 5852 15804
rect 5852 15748 5908 15804
rect 5908 15748 5912 15804
rect 5848 15744 5912 15748
rect 5928 15804 5992 15808
rect 5928 15748 5932 15804
rect 5932 15748 5988 15804
rect 5988 15748 5992 15804
rect 5928 15744 5992 15748
rect 6008 15804 6072 15808
rect 6008 15748 6012 15804
rect 6012 15748 6068 15804
rect 6068 15748 6072 15804
rect 6008 15744 6072 15748
rect 6088 15804 6152 15808
rect 6088 15748 6092 15804
rect 6092 15748 6148 15804
rect 6148 15748 6152 15804
rect 6088 15744 6152 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 9272 15804 9336 15808
rect 9272 15748 9276 15804
rect 9276 15748 9332 15804
rect 9332 15748 9336 15804
rect 9272 15744 9336 15748
rect 9352 15804 9416 15808
rect 9352 15748 9356 15804
rect 9356 15748 9412 15804
rect 9412 15748 9416 15804
rect 9352 15744 9416 15748
rect 3372 15736 3436 15740
rect 3372 15680 3422 15736
rect 3422 15680 3436 15736
rect 3372 15676 3436 15680
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 7480 15260 7544 15264
rect 7480 15204 7484 15260
rect 7484 15204 7540 15260
rect 7540 15204 7544 15260
rect 7480 15200 7544 15204
rect 7560 15260 7624 15264
rect 7560 15204 7564 15260
rect 7564 15204 7620 15260
rect 7620 15204 7624 15260
rect 7560 15200 7624 15204
rect 7640 15260 7704 15264
rect 7640 15204 7644 15260
rect 7644 15204 7700 15260
rect 7700 15204 7704 15260
rect 7640 15200 7704 15204
rect 7720 15260 7784 15264
rect 7720 15204 7724 15260
rect 7724 15204 7780 15260
rect 7780 15204 7784 15260
rect 7720 15200 7784 15204
rect 2584 14716 2648 14720
rect 2584 14660 2588 14716
rect 2588 14660 2644 14716
rect 2644 14660 2648 14716
rect 2584 14656 2648 14660
rect 2664 14716 2728 14720
rect 2664 14660 2668 14716
rect 2668 14660 2724 14716
rect 2724 14660 2728 14716
rect 2664 14656 2728 14660
rect 2744 14716 2808 14720
rect 2744 14660 2748 14716
rect 2748 14660 2804 14716
rect 2804 14660 2808 14716
rect 2744 14656 2808 14660
rect 2824 14716 2888 14720
rect 2824 14660 2828 14716
rect 2828 14660 2884 14716
rect 2884 14660 2888 14716
rect 2824 14656 2888 14660
rect 5848 14716 5912 14720
rect 5848 14660 5852 14716
rect 5852 14660 5908 14716
rect 5908 14660 5912 14716
rect 5848 14656 5912 14660
rect 5928 14716 5992 14720
rect 5928 14660 5932 14716
rect 5932 14660 5988 14716
rect 5988 14660 5992 14716
rect 5928 14656 5992 14660
rect 6008 14716 6072 14720
rect 6008 14660 6012 14716
rect 6012 14660 6068 14716
rect 6068 14660 6072 14716
rect 6008 14656 6072 14660
rect 6088 14716 6152 14720
rect 6088 14660 6092 14716
rect 6092 14660 6148 14716
rect 6148 14660 6152 14716
rect 6088 14656 6152 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 9272 14716 9336 14720
rect 9272 14660 9276 14716
rect 9276 14660 9332 14716
rect 9332 14660 9336 14716
rect 9272 14656 9336 14660
rect 9352 14716 9416 14720
rect 9352 14660 9356 14716
rect 9356 14660 9412 14716
rect 9412 14660 9416 14716
rect 9352 14656 9416 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 7480 14172 7544 14176
rect 7480 14116 7484 14172
rect 7484 14116 7540 14172
rect 7540 14116 7544 14172
rect 7480 14112 7544 14116
rect 7560 14172 7624 14176
rect 7560 14116 7564 14172
rect 7564 14116 7620 14172
rect 7620 14116 7624 14172
rect 7560 14112 7624 14116
rect 7640 14172 7704 14176
rect 7640 14116 7644 14172
rect 7644 14116 7700 14172
rect 7700 14116 7704 14172
rect 7640 14112 7704 14116
rect 7720 14172 7784 14176
rect 7720 14116 7724 14172
rect 7724 14116 7780 14172
rect 7780 14116 7784 14172
rect 7720 14112 7784 14116
rect 3556 14104 3620 14108
rect 3556 14048 3606 14104
rect 3606 14048 3620 14104
rect 3556 14044 3620 14048
rect 2584 13628 2648 13632
rect 2584 13572 2588 13628
rect 2588 13572 2644 13628
rect 2644 13572 2648 13628
rect 2584 13568 2648 13572
rect 2664 13628 2728 13632
rect 2664 13572 2668 13628
rect 2668 13572 2724 13628
rect 2724 13572 2728 13628
rect 2664 13568 2728 13572
rect 2744 13628 2808 13632
rect 2744 13572 2748 13628
rect 2748 13572 2804 13628
rect 2804 13572 2808 13628
rect 2744 13568 2808 13572
rect 2824 13628 2888 13632
rect 2824 13572 2828 13628
rect 2828 13572 2884 13628
rect 2884 13572 2888 13628
rect 2824 13568 2888 13572
rect 5848 13628 5912 13632
rect 5848 13572 5852 13628
rect 5852 13572 5908 13628
rect 5908 13572 5912 13628
rect 5848 13568 5912 13572
rect 5928 13628 5992 13632
rect 5928 13572 5932 13628
rect 5932 13572 5988 13628
rect 5988 13572 5992 13628
rect 5928 13568 5992 13572
rect 6008 13628 6072 13632
rect 6008 13572 6012 13628
rect 6012 13572 6068 13628
rect 6068 13572 6072 13628
rect 6008 13568 6072 13572
rect 6088 13628 6152 13632
rect 6088 13572 6092 13628
rect 6092 13572 6148 13628
rect 6148 13572 6152 13628
rect 6088 13568 6152 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 9272 13628 9336 13632
rect 9272 13572 9276 13628
rect 9276 13572 9332 13628
rect 9332 13572 9336 13628
rect 9272 13568 9336 13572
rect 9352 13628 9416 13632
rect 9352 13572 9356 13628
rect 9356 13572 9412 13628
rect 9412 13572 9416 13628
rect 9352 13568 9416 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 7480 13084 7544 13088
rect 7480 13028 7484 13084
rect 7484 13028 7540 13084
rect 7540 13028 7544 13084
rect 7480 13024 7544 13028
rect 7560 13084 7624 13088
rect 7560 13028 7564 13084
rect 7564 13028 7620 13084
rect 7620 13028 7624 13084
rect 7560 13024 7624 13028
rect 7640 13084 7704 13088
rect 7640 13028 7644 13084
rect 7644 13028 7700 13084
rect 7700 13028 7704 13084
rect 7640 13024 7704 13028
rect 7720 13084 7784 13088
rect 7720 13028 7724 13084
rect 7724 13028 7780 13084
rect 7780 13028 7784 13084
rect 7720 13024 7784 13028
rect 2584 12540 2648 12544
rect 2584 12484 2588 12540
rect 2588 12484 2644 12540
rect 2644 12484 2648 12540
rect 2584 12480 2648 12484
rect 2664 12540 2728 12544
rect 2664 12484 2668 12540
rect 2668 12484 2724 12540
rect 2724 12484 2728 12540
rect 2664 12480 2728 12484
rect 2744 12540 2808 12544
rect 2744 12484 2748 12540
rect 2748 12484 2804 12540
rect 2804 12484 2808 12540
rect 2744 12480 2808 12484
rect 2824 12540 2888 12544
rect 2824 12484 2828 12540
rect 2828 12484 2884 12540
rect 2884 12484 2888 12540
rect 2824 12480 2888 12484
rect 5848 12540 5912 12544
rect 5848 12484 5852 12540
rect 5852 12484 5908 12540
rect 5908 12484 5912 12540
rect 5848 12480 5912 12484
rect 5928 12540 5992 12544
rect 5928 12484 5932 12540
rect 5932 12484 5988 12540
rect 5988 12484 5992 12540
rect 5928 12480 5992 12484
rect 6008 12540 6072 12544
rect 6008 12484 6012 12540
rect 6012 12484 6068 12540
rect 6068 12484 6072 12540
rect 6008 12480 6072 12484
rect 6088 12540 6152 12544
rect 6088 12484 6092 12540
rect 6092 12484 6148 12540
rect 6148 12484 6152 12540
rect 6088 12480 6152 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 9272 12540 9336 12544
rect 9272 12484 9276 12540
rect 9276 12484 9332 12540
rect 9332 12484 9336 12540
rect 9272 12480 9336 12484
rect 9352 12540 9416 12544
rect 9352 12484 9356 12540
rect 9356 12484 9412 12540
rect 9412 12484 9416 12540
rect 9352 12480 9416 12484
rect 3556 12412 3620 12476
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 7480 11996 7544 12000
rect 7480 11940 7484 11996
rect 7484 11940 7540 11996
rect 7540 11940 7544 11996
rect 7480 11936 7544 11940
rect 7560 11996 7624 12000
rect 7560 11940 7564 11996
rect 7564 11940 7620 11996
rect 7620 11940 7624 11996
rect 7560 11936 7624 11940
rect 7640 11996 7704 12000
rect 7640 11940 7644 11996
rect 7644 11940 7700 11996
rect 7700 11940 7704 11996
rect 7640 11936 7704 11940
rect 7720 11996 7784 12000
rect 7720 11940 7724 11996
rect 7724 11940 7780 11996
rect 7780 11940 7784 11996
rect 7720 11936 7784 11940
rect 3004 11792 3068 11796
rect 3004 11736 3054 11792
rect 3054 11736 3068 11792
rect 3004 11732 3068 11736
rect 3372 11460 3436 11524
rect 2584 11452 2648 11456
rect 2584 11396 2588 11452
rect 2588 11396 2644 11452
rect 2644 11396 2648 11452
rect 2584 11392 2648 11396
rect 2664 11452 2728 11456
rect 2664 11396 2668 11452
rect 2668 11396 2724 11452
rect 2724 11396 2728 11452
rect 2664 11392 2728 11396
rect 2744 11452 2808 11456
rect 2744 11396 2748 11452
rect 2748 11396 2804 11452
rect 2804 11396 2808 11452
rect 2744 11392 2808 11396
rect 2824 11452 2888 11456
rect 2824 11396 2828 11452
rect 2828 11396 2884 11452
rect 2884 11396 2888 11452
rect 2824 11392 2888 11396
rect 5848 11452 5912 11456
rect 5848 11396 5852 11452
rect 5852 11396 5908 11452
rect 5908 11396 5912 11452
rect 5848 11392 5912 11396
rect 5928 11452 5992 11456
rect 5928 11396 5932 11452
rect 5932 11396 5988 11452
rect 5988 11396 5992 11452
rect 5928 11392 5992 11396
rect 6008 11452 6072 11456
rect 6008 11396 6012 11452
rect 6012 11396 6068 11452
rect 6068 11396 6072 11452
rect 6008 11392 6072 11396
rect 6088 11452 6152 11456
rect 6088 11396 6092 11452
rect 6092 11396 6148 11452
rect 6148 11396 6152 11452
rect 6088 11392 6152 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 9272 11452 9336 11456
rect 9272 11396 9276 11452
rect 9276 11396 9332 11452
rect 9332 11396 9336 11452
rect 9272 11392 9336 11396
rect 9352 11452 9416 11456
rect 9352 11396 9356 11452
rect 9356 11396 9412 11452
rect 9412 11396 9416 11452
rect 9352 11392 9416 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 7480 10908 7544 10912
rect 7480 10852 7484 10908
rect 7484 10852 7540 10908
rect 7540 10852 7544 10908
rect 7480 10848 7544 10852
rect 7560 10908 7624 10912
rect 7560 10852 7564 10908
rect 7564 10852 7620 10908
rect 7620 10852 7624 10908
rect 7560 10848 7624 10852
rect 7640 10908 7704 10912
rect 7640 10852 7644 10908
rect 7644 10852 7700 10908
rect 7700 10852 7704 10908
rect 7640 10848 7704 10852
rect 7720 10908 7784 10912
rect 7720 10852 7724 10908
rect 7724 10852 7780 10908
rect 7780 10852 7784 10908
rect 7720 10848 7784 10852
rect 2584 10364 2648 10368
rect 2584 10308 2588 10364
rect 2588 10308 2644 10364
rect 2644 10308 2648 10364
rect 2584 10304 2648 10308
rect 2664 10364 2728 10368
rect 2664 10308 2668 10364
rect 2668 10308 2724 10364
rect 2724 10308 2728 10364
rect 2664 10304 2728 10308
rect 2744 10364 2808 10368
rect 2744 10308 2748 10364
rect 2748 10308 2804 10364
rect 2804 10308 2808 10364
rect 2744 10304 2808 10308
rect 2824 10364 2888 10368
rect 2824 10308 2828 10364
rect 2828 10308 2884 10364
rect 2884 10308 2888 10364
rect 2824 10304 2888 10308
rect 5848 10364 5912 10368
rect 5848 10308 5852 10364
rect 5852 10308 5908 10364
rect 5908 10308 5912 10364
rect 5848 10304 5912 10308
rect 5928 10364 5992 10368
rect 5928 10308 5932 10364
rect 5932 10308 5988 10364
rect 5988 10308 5992 10364
rect 5928 10304 5992 10308
rect 6008 10364 6072 10368
rect 6008 10308 6012 10364
rect 6012 10308 6068 10364
rect 6068 10308 6072 10364
rect 6008 10304 6072 10308
rect 6088 10364 6152 10368
rect 6088 10308 6092 10364
rect 6092 10308 6148 10364
rect 6148 10308 6152 10364
rect 6088 10304 6152 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 9272 10364 9336 10368
rect 9272 10308 9276 10364
rect 9276 10308 9332 10364
rect 9332 10308 9336 10364
rect 9272 10304 9336 10308
rect 9352 10364 9416 10368
rect 9352 10308 9356 10364
rect 9356 10308 9412 10364
rect 9412 10308 9416 10364
rect 9352 10304 9416 10308
rect 3924 10296 3988 10300
rect 3924 10240 3974 10296
rect 3974 10240 3988 10296
rect 3924 10236 3988 10240
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 7480 9820 7544 9824
rect 7480 9764 7484 9820
rect 7484 9764 7540 9820
rect 7540 9764 7544 9820
rect 7480 9760 7544 9764
rect 7560 9820 7624 9824
rect 7560 9764 7564 9820
rect 7564 9764 7620 9820
rect 7620 9764 7624 9820
rect 7560 9760 7624 9764
rect 7640 9820 7704 9824
rect 7640 9764 7644 9820
rect 7644 9764 7700 9820
rect 7700 9764 7704 9820
rect 7640 9760 7704 9764
rect 7720 9820 7784 9824
rect 7720 9764 7724 9820
rect 7724 9764 7780 9820
rect 7780 9764 7784 9820
rect 7720 9760 7784 9764
rect 2584 9276 2648 9280
rect 2584 9220 2588 9276
rect 2588 9220 2644 9276
rect 2644 9220 2648 9276
rect 2584 9216 2648 9220
rect 2664 9276 2728 9280
rect 2664 9220 2668 9276
rect 2668 9220 2724 9276
rect 2724 9220 2728 9276
rect 2664 9216 2728 9220
rect 2744 9276 2808 9280
rect 2744 9220 2748 9276
rect 2748 9220 2804 9276
rect 2804 9220 2808 9276
rect 2744 9216 2808 9220
rect 2824 9276 2888 9280
rect 2824 9220 2828 9276
rect 2828 9220 2884 9276
rect 2884 9220 2888 9276
rect 2824 9216 2888 9220
rect 5848 9276 5912 9280
rect 5848 9220 5852 9276
rect 5852 9220 5908 9276
rect 5908 9220 5912 9276
rect 5848 9216 5912 9220
rect 5928 9276 5992 9280
rect 5928 9220 5932 9276
rect 5932 9220 5988 9276
rect 5988 9220 5992 9276
rect 5928 9216 5992 9220
rect 6008 9276 6072 9280
rect 6008 9220 6012 9276
rect 6012 9220 6068 9276
rect 6068 9220 6072 9276
rect 6008 9216 6072 9220
rect 6088 9276 6152 9280
rect 6088 9220 6092 9276
rect 6092 9220 6148 9276
rect 6148 9220 6152 9276
rect 6088 9216 6152 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 9272 9276 9336 9280
rect 9272 9220 9276 9276
rect 9276 9220 9332 9276
rect 9332 9220 9336 9276
rect 9272 9216 9336 9220
rect 9352 9276 9416 9280
rect 9352 9220 9356 9276
rect 9356 9220 9412 9276
rect 9412 9220 9416 9276
rect 9352 9216 9416 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 7480 8732 7544 8736
rect 7480 8676 7484 8732
rect 7484 8676 7540 8732
rect 7540 8676 7544 8732
rect 7480 8672 7544 8676
rect 7560 8732 7624 8736
rect 7560 8676 7564 8732
rect 7564 8676 7620 8732
rect 7620 8676 7624 8732
rect 7560 8672 7624 8676
rect 7640 8732 7704 8736
rect 7640 8676 7644 8732
rect 7644 8676 7700 8732
rect 7700 8676 7704 8732
rect 7640 8672 7704 8676
rect 7720 8732 7784 8736
rect 7720 8676 7724 8732
rect 7724 8676 7780 8732
rect 7780 8676 7784 8732
rect 7720 8672 7784 8676
rect 2584 8188 2648 8192
rect 2584 8132 2588 8188
rect 2588 8132 2644 8188
rect 2644 8132 2648 8188
rect 2584 8128 2648 8132
rect 2664 8188 2728 8192
rect 2664 8132 2668 8188
rect 2668 8132 2724 8188
rect 2724 8132 2728 8188
rect 2664 8128 2728 8132
rect 2744 8188 2808 8192
rect 2744 8132 2748 8188
rect 2748 8132 2804 8188
rect 2804 8132 2808 8188
rect 2744 8128 2808 8132
rect 2824 8188 2888 8192
rect 2824 8132 2828 8188
rect 2828 8132 2884 8188
rect 2884 8132 2888 8188
rect 2824 8128 2888 8132
rect 5848 8188 5912 8192
rect 5848 8132 5852 8188
rect 5852 8132 5908 8188
rect 5908 8132 5912 8188
rect 5848 8128 5912 8132
rect 5928 8188 5992 8192
rect 5928 8132 5932 8188
rect 5932 8132 5988 8188
rect 5988 8132 5992 8188
rect 5928 8128 5992 8132
rect 6008 8188 6072 8192
rect 6008 8132 6012 8188
rect 6012 8132 6068 8188
rect 6068 8132 6072 8188
rect 6008 8128 6072 8132
rect 6088 8188 6152 8192
rect 6088 8132 6092 8188
rect 6092 8132 6148 8188
rect 6148 8132 6152 8188
rect 6088 8128 6152 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 9272 8188 9336 8192
rect 9272 8132 9276 8188
rect 9276 8132 9332 8188
rect 9332 8132 9336 8188
rect 9272 8128 9336 8132
rect 9352 8188 9416 8192
rect 9352 8132 9356 8188
rect 9356 8132 9412 8188
rect 9412 8132 9416 8188
rect 9352 8128 9416 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 7480 7644 7544 7648
rect 7480 7588 7484 7644
rect 7484 7588 7540 7644
rect 7540 7588 7544 7644
rect 7480 7584 7544 7588
rect 7560 7644 7624 7648
rect 7560 7588 7564 7644
rect 7564 7588 7620 7644
rect 7620 7588 7624 7644
rect 7560 7584 7624 7588
rect 7640 7644 7704 7648
rect 7640 7588 7644 7644
rect 7644 7588 7700 7644
rect 7700 7588 7704 7644
rect 7640 7584 7704 7588
rect 7720 7644 7784 7648
rect 7720 7588 7724 7644
rect 7724 7588 7780 7644
rect 7780 7588 7784 7644
rect 7720 7584 7784 7588
rect 2584 7100 2648 7104
rect 2584 7044 2588 7100
rect 2588 7044 2644 7100
rect 2644 7044 2648 7100
rect 2584 7040 2648 7044
rect 2664 7100 2728 7104
rect 2664 7044 2668 7100
rect 2668 7044 2724 7100
rect 2724 7044 2728 7100
rect 2664 7040 2728 7044
rect 2744 7100 2808 7104
rect 2744 7044 2748 7100
rect 2748 7044 2804 7100
rect 2804 7044 2808 7100
rect 2744 7040 2808 7044
rect 2824 7100 2888 7104
rect 2824 7044 2828 7100
rect 2828 7044 2884 7100
rect 2884 7044 2888 7100
rect 2824 7040 2888 7044
rect 5848 7100 5912 7104
rect 5848 7044 5852 7100
rect 5852 7044 5908 7100
rect 5908 7044 5912 7100
rect 5848 7040 5912 7044
rect 5928 7100 5992 7104
rect 5928 7044 5932 7100
rect 5932 7044 5988 7100
rect 5988 7044 5992 7100
rect 5928 7040 5992 7044
rect 6008 7100 6072 7104
rect 6008 7044 6012 7100
rect 6012 7044 6068 7100
rect 6068 7044 6072 7100
rect 6008 7040 6072 7044
rect 6088 7100 6152 7104
rect 6088 7044 6092 7100
rect 6092 7044 6148 7100
rect 6148 7044 6152 7100
rect 6088 7040 6152 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 9272 7100 9336 7104
rect 9272 7044 9276 7100
rect 9276 7044 9332 7100
rect 9332 7044 9336 7100
rect 9272 7040 9336 7044
rect 9352 7100 9416 7104
rect 9352 7044 9356 7100
rect 9356 7044 9412 7100
rect 9412 7044 9416 7100
rect 9352 7040 9416 7044
rect 5028 6700 5092 6764
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 7480 6556 7544 6560
rect 7480 6500 7484 6556
rect 7484 6500 7540 6556
rect 7540 6500 7544 6556
rect 7480 6496 7544 6500
rect 7560 6556 7624 6560
rect 7560 6500 7564 6556
rect 7564 6500 7620 6556
rect 7620 6500 7624 6556
rect 7560 6496 7624 6500
rect 7640 6556 7704 6560
rect 7640 6500 7644 6556
rect 7644 6500 7700 6556
rect 7700 6500 7704 6556
rect 7640 6496 7704 6500
rect 7720 6556 7784 6560
rect 7720 6500 7724 6556
rect 7724 6500 7780 6556
rect 7780 6500 7784 6556
rect 7720 6496 7784 6500
rect 2584 6012 2648 6016
rect 2584 5956 2588 6012
rect 2588 5956 2644 6012
rect 2644 5956 2648 6012
rect 2584 5952 2648 5956
rect 2664 6012 2728 6016
rect 2664 5956 2668 6012
rect 2668 5956 2724 6012
rect 2724 5956 2728 6012
rect 2664 5952 2728 5956
rect 2744 6012 2808 6016
rect 2744 5956 2748 6012
rect 2748 5956 2804 6012
rect 2804 5956 2808 6012
rect 2744 5952 2808 5956
rect 2824 6012 2888 6016
rect 2824 5956 2828 6012
rect 2828 5956 2884 6012
rect 2884 5956 2888 6012
rect 2824 5952 2888 5956
rect 5848 6012 5912 6016
rect 5848 5956 5852 6012
rect 5852 5956 5908 6012
rect 5908 5956 5912 6012
rect 5848 5952 5912 5956
rect 5928 6012 5992 6016
rect 5928 5956 5932 6012
rect 5932 5956 5988 6012
rect 5988 5956 5992 6012
rect 5928 5952 5992 5956
rect 6008 6012 6072 6016
rect 6008 5956 6012 6012
rect 6012 5956 6068 6012
rect 6068 5956 6072 6012
rect 6008 5952 6072 5956
rect 6088 6012 6152 6016
rect 6088 5956 6092 6012
rect 6092 5956 6148 6012
rect 6148 5956 6152 6012
rect 6088 5952 6152 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 9272 6012 9336 6016
rect 9272 5956 9276 6012
rect 9276 5956 9332 6012
rect 9332 5956 9336 6012
rect 9272 5952 9336 5956
rect 9352 6012 9416 6016
rect 9352 5956 9356 6012
rect 9356 5956 9412 6012
rect 9412 5956 9416 6012
rect 9352 5952 9416 5956
rect 4660 5884 4724 5948
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 7480 5468 7544 5472
rect 7480 5412 7484 5468
rect 7484 5412 7540 5468
rect 7540 5412 7544 5468
rect 7480 5408 7544 5412
rect 7560 5468 7624 5472
rect 7560 5412 7564 5468
rect 7564 5412 7620 5468
rect 7620 5412 7624 5468
rect 7560 5408 7624 5412
rect 7640 5468 7704 5472
rect 7640 5412 7644 5468
rect 7644 5412 7700 5468
rect 7700 5412 7704 5468
rect 7640 5408 7704 5412
rect 7720 5468 7784 5472
rect 7720 5412 7724 5468
rect 7724 5412 7780 5468
rect 7780 5412 7784 5468
rect 7720 5408 7784 5412
rect 4844 5204 4908 5268
rect 2584 4924 2648 4928
rect 2584 4868 2588 4924
rect 2588 4868 2644 4924
rect 2644 4868 2648 4924
rect 2584 4864 2648 4868
rect 2664 4924 2728 4928
rect 2664 4868 2668 4924
rect 2668 4868 2724 4924
rect 2724 4868 2728 4924
rect 2664 4864 2728 4868
rect 2744 4924 2808 4928
rect 2744 4868 2748 4924
rect 2748 4868 2804 4924
rect 2804 4868 2808 4924
rect 2744 4864 2808 4868
rect 2824 4924 2888 4928
rect 2824 4868 2828 4924
rect 2828 4868 2884 4924
rect 2884 4868 2888 4924
rect 2824 4864 2888 4868
rect 5848 4924 5912 4928
rect 5848 4868 5852 4924
rect 5852 4868 5908 4924
rect 5908 4868 5912 4924
rect 5848 4864 5912 4868
rect 5928 4924 5992 4928
rect 5928 4868 5932 4924
rect 5932 4868 5988 4924
rect 5988 4868 5992 4924
rect 5928 4864 5992 4868
rect 6008 4924 6072 4928
rect 6008 4868 6012 4924
rect 6012 4868 6068 4924
rect 6068 4868 6072 4924
rect 6008 4864 6072 4868
rect 6088 4924 6152 4928
rect 6088 4868 6092 4924
rect 6092 4868 6148 4924
rect 6148 4868 6152 4924
rect 6088 4864 6152 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 9272 4924 9336 4928
rect 9272 4868 9276 4924
rect 9276 4868 9332 4924
rect 9332 4868 9336 4924
rect 9272 4864 9336 4868
rect 9352 4924 9416 4928
rect 9352 4868 9356 4924
rect 9356 4868 9412 4924
rect 9412 4868 9416 4924
rect 9352 4864 9416 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 7480 4380 7544 4384
rect 7480 4324 7484 4380
rect 7484 4324 7540 4380
rect 7540 4324 7544 4380
rect 7480 4320 7544 4324
rect 7560 4380 7624 4384
rect 7560 4324 7564 4380
rect 7564 4324 7620 4380
rect 7620 4324 7624 4380
rect 7560 4320 7624 4324
rect 7640 4380 7704 4384
rect 7640 4324 7644 4380
rect 7644 4324 7700 4380
rect 7700 4324 7704 4380
rect 7640 4320 7704 4324
rect 7720 4380 7784 4384
rect 7720 4324 7724 4380
rect 7724 4324 7780 4380
rect 7780 4324 7784 4380
rect 7720 4320 7784 4324
rect 2584 3836 2648 3840
rect 2584 3780 2588 3836
rect 2588 3780 2644 3836
rect 2644 3780 2648 3836
rect 2584 3776 2648 3780
rect 2664 3836 2728 3840
rect 2664 3780 2668 3836
rect 2668 3780 2724 3836
rect 2724 3780 2728 3836
rect 2664 3776 2728 3780
rect 2744 3836 2808 3840
rect 2744 3780 2748 3836
rect 2748 3780 2804 3836
rect 2804 3780 2808 3836
rect 2744 3776 2808 3780
rect 2824 3836 2888 3840
rect 2824 3780 2828 3836
rect 2828 3780 2884 3836
rect 2884 3780 2888 3836
rect 2824 3776 2888 3780
rect 5848 3836 5912 3840
rect 5848 3780 5852 3836
rect 5852 3780 5908 3836
rect 5908 3780 5912 3836
rect 5848 3776 5912 3780
rect 5928 3836 5992 3840
rect 5928 3780 5932 3836
rect 5932 3780 5988 3836
rect 5988 3780 5992 3836
rect 5928 3776 5992 3780
rect 6008 3836 6072 3840
rect 6008 3780 6012 3836
rect 6012 3780 6068 3836
rect 6068 3780 6072 3836
rect 6008 3776 6072 3780
rect 6088 3836 6152 3840
rect 6088 3780 6092 3836
rect 6092 3780 6148 3836
rect 6148 3780 6152 3836
rect 6088 3776 6152 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 9272 3836 9336 3840
rect 9272 3780 9276 3836
rect 9276 3780 9332 3836
rect 9332 3780 9336 3836
rect 9272 3776 9336 3780
rect 9352 3836 9416 3840
rect 9352 3780 9356 3836
rect 9356 3780 9412 3836
rect 9412 3780 9416 3836
rect 9352 3776 9416 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 7480 3292 7544 3296
rect 7480 3236 7484 3292
rect 7484 3236 7540 3292
rect 7540 3236 7544 3292
rect 7480 3232 7544 3236
rect 7560 3292 7624 3296
rect 7560 3236 7564 3292
rect 7564 3236 7620 3292
rect 7620 3236 7624 3292
rect 7560 3232 7624 3236
rect 7640 3292 7704 3296
rect 7640 3236 7644 3292
rect 7644 3236 7700 3292
rect 7700 3236 7704 3292
rect 7640 3232 7704 3236
rect 7720 3292 7784 3296
rect 7720 3236 7724 3292
rect 7724 3236 7780 3292
rect 7780 3236 7784 3292
rect 7720 3232 7784 3236
rect 2584 2748 2648 2752
rect 2584 2692 2588 2748
rect 2588 2692 2644 2748
rect 2644 2692 2648 2748
rect 2584 2688 2648 2692
rect 2664 2748 2728 2752
rect 2664 2692 2668 2748
rect 2668 2692 2724 2748
rect 2724 2692 2728 2748
rect 2664 2688 2728 2692
rect 2744 2748 2808 2752
rect 2744 2692 2748 2748
rect 2748 2692 2804 2748
rect 2804 2692 2808 2748
rect 2744 2688 2808 2692
rect 2824 2748 2888 2752
rect 2824 2692 2828 2748
rect 2828 2692 2884 2748
rect 2884 2692 2888 2748
rect 2824 2688 2888 2692
rect 5848 2748 5912 2752
rect 5848 2692 5852 2748
rect 5852 2692 5908 2748
rect 5908 2692 5912 2748
rect 5848 2688 5912 2692
rect 5928 2748 5992 2752
rect 5928 2692 5932 2748
rect 5932 2692 5988 2748
rect 5988 2692 5992 2748
rect 5928 2688 5992 2692
rect 6008 2748 6072 2752
rect 6008 2692 6012 2748
rect 6012 2692 6068 2748
rect 6068 2692 6072 2748
rect 6008 2688 6072 2692
rect 6088 2748 6152 2752
rect 6088 2692 6092 2748
rect 6092 2692 6148 2748
rect 6148 2692 6152 2748
rect 6088 2688 6152 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 9272 2748 9336 2752
rect 9272 2692 9276 2748
rect 9276 2692 9332 2748
rect 9332 2692 9336 2748
rect 9272 2688 9336 2692
rect 9352 2748 9416 2752
rect 9352 2692 9356 2748
rect 9356 2692 9412 2748
rect 9412 2692 9416 2748
rect 9352 2688 9416 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 7480 2204 7544 2208
rect 7480 2148 7484 2204
rect 7484 2148 7540 2204
rect 7540 2148 7544 2204
rect 7480 2144 7544 2148
rect 7560 2204 7624 2208
rect 7560 2148 7564 2204
rect 7564 2148 7620 2204
rect 7620 2148 7624 2204
rect 7560 2144 7624 2148
rect 7640 2204 7704 2208
rect 7640 2148 7644 2204
rect 7644 2148 7700 2204
rect 7700 2148 7704 2204
rect 7640 2144 7704 2148
rect 7720 2204 7784 2208
rect 7720 2148 7724 2204
rect 7724 2148 7780 2204
rect 7780 2148 7784 2204
rect 7720 2144 7784 2148
<< metal4 >>
rect 2576 77824 2896 77840
rect 2576 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2576 76736 2896 77760
rect 2576 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2576 75648 2896 76672
rect 2576 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2083 74764 2149 74765
rect 2083 74700 2084 74764
rect 2148 74700 2149 74764
rect 2083 74699 2149 74700
rect 1899 72724 1965 72725
rect 1899 72660 1900 72724
rect 1964 72660 1965 72724
rect 1899 72659 1965 72660
rect 1531 72180 1597 72181
rect 1531 72116 1532 72180
rect 1596 72116 1597 72180
rect 1531 72115 1597 72116
rect 1534 70413 1594 72115
rect 1531 70412 1597 70413
rect 1531 70348 1532 70412
rect 1596 70348 1597 70412
rect 1531 70347 1597 70348
rect 1902 70277 1962 72659
rect 1899 70276 1965 70277
rect 1899 70212 1900 70276
rect 1964 70212 1965 70276
rect 1899 70211 1965 70212
rect 1347 70004 1413 70005
rect 1347 69940 1348 70004
rect 1412 69940 1413 70004
rect 1347 69939 1413 69940
rect 1350 60349 1410 69939
rect 1531 66332 1597 66333
rect 1531 66268 1532 66332
rect 1596 66268 1597 66332
rect 1531 66267 1597 66268
rect 1347 60348 1413 60349
rect 1347 60284 1348 60348
rect 1412 60284 1413 60348
rect 1347 60283 1413 60284
rect 979 57900 1045 57901
rect 979 57836 980 57900
rect 1044 57836 1045 57900
rect 979 57835 1045 57836
rect 982 57762 1042 57835
rect 430 57702 1042 57762
rect 1163 57764 1229 57765
rect 243 53548 309 53549
rect 243 53484 244 53548
rect 308 53484 309 53548
rect 243 53483 309 53484
rect 246 39949 306 53483
rect 430 50149 490 57702
rect 1163 57700 1164 57764
rect 1228 57700 1229 57764
rect 1163 57699 1229 57700
rect 1166 57221 1226 57699
rect 1347 57492 1413 57493
rect 1347 57428 1348 57492
rect 1412 57428 1413 57492
rect 1347 57427 1413 57428
rect 1163 57220 1229 57221
rect 1163 57156 1164 57220
rect 1228 57156 1229 57220
rect 1163 57155 1229 57156
rect 1350 57085 1410 57427
rect 1347 57084 1413 57085
rect 1347 57020 1348 57084
rect 1412 57020 1413 57084
rect 1347 57019 1413 57020
rect 795 56948 861 56949
rect 795 56884 796 56948
rect 860 56884 861 56948
rect 795 56883 861 56884
rect 611 50998 677 50999
rect 611 50934 612 50998
rect 676 50934 677 50998
rect 611 50933 677 50934
rect 427 50148 493 50149
rect 427 50084 428 50148
rect 492 50084 493 50148
rect 427 50083 493 50084
rect 427 46748 493 46749
rect 427 46684 428 46748
rect 492 46684 493 46748
rect 427 46683 493 46684
rect 430 39949 490 46683
rect 614 45831 674 50933
rect 611 45830 677 45831
rect 611 45766 612 45830
rect 676 45766 677 45830
rect 611 45765 677 45766
rect 798 43349 858 56883
rect 1163 56812 1229 56813
rect 1163 56748 1164 56812
rect 1228 56748 1229 56812
rect 1163 56747 1229 56748
rect 979 52596 1045 52597
rect 979 52532 980 52596
rect 1044 52532 1045 52596
rect 979 52531 1045 52532
rect 795 43348 861 43349
rect 795 43284 796 43348
rect 860 43284 861 43348
rect 795 43283 861 43284
rect 243 39948 309 39949
rect 243 39884 244 39948
rect 308 39884 309 39948
rect 243 39883 309 39884
rect 427 39948 493 39949
rect 427 39884 428 39948
rect 492 39884 493 39948
rect 427 39883 493 39884
rect 982 31109 1042 52531
rect 1166 51509 1226 56747
rect 1347 54908 1413 54909
rect 1347 54844 1348 54908
rect 1412 54844 1413 54908
rect 1347 54843 1413 54844
rect 1163 51508 1229 51509
rect 1163 51444 1164 51508
rect 1228 51444 1229 51508
rect 1163 51443 1229 51444
rect 1163 49740 1229 49741
rect 1163 49676 1164 49740
rect 1228 49676 1229 49740
rect 1163 49675 1229 49676
rect 979 31108 1045 31109
rect 979 31044 980 31108
rect 1044 31044 1045 31108
rect 979 31043 1045 31044
rect 1166 30293 1226 49675
rect 1350 48109 1410 54843
rect 1534 50421 1594 66267
rect 1715 64972 1781 64973
rect 1715 64908 1716 64972
rect 1780 64908 1781 64972
rect 1715 64907 1781 64908
rect 1531 50420 1597 50421
rect 1531 50356 1532 50420
rect 1596 50356 1597 50420
rect 1531 50355 1597 50356
rect 1531 50148 1597 50149
rect 1531 50084 1532 50148
rect 1596 50084 1597 50148
rect 1531 50083 1597 50084
rect 1534 48517 1594 50083
rect 1718 49605 1778 64907
rect 1899 62660 1965 62661
rect 1899 62596 1900 62660
rect 1964 62596 1965 62660
rect 1899 62595 1965 62596
rect 1902 55589 1962 62595
rect 2086 60213 2146 74699
rect 2576 74560 2896 75584
rect 2576 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2576 73472 2896 74496
rect 2576 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2576 72384 2896 73408
rect 2576 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2576 71296 2896 72320
rect 2576 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2267 70684 2333 70685
rect 2267 70620 2268 70684
rect 2332 70620 2333 70684
rect 2267 70619 2333 70620
rect 2270 70277 2330 70619
rect 2267 70276 2333 70277
rect 2267 70212 2268 70276
rect 2332 70212 2333 70276
rect 2267 70211 2333 70212
rect 2576 70208 2896 71232
rect 2576 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2267 70140 2333 70141
rect 2267 70076 2268 70140
rect 2332 70076 2333 70140
rect 2267 70075 2333 70076
rect 2270 62933 2330 70075
rect 2576 69120 2896 70144
rect 2576 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2576 68032 2896 69056
rect 2576 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2576 66944 2896 67968
rect 2576 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2576 65856 2896 66880
rect 4208 77280 4528 77840
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 76192 4528 77216
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 75104 4528 76128
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 74016 4528 75040
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 72928 4528 73952
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 71840 4528 72864
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 70752 4528 71776
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 69664 4528 70688
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 68576 4528 69600
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 67488 4528 68512
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 66400 4528 67424
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 3739 66060 3805 66061
rect 3739 65996 3740 66060
rect 3804 65996 3805 66060
rect 3739 65995 3805 65996
rect 2576 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2576 64768 2896 65792
rect 3555 65108 3621 65109
rect 3555 65044 3556 65108
rect 3620 65044 3621 65108
rect 3555 65043 3621 65044
rect 2576 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2576 63680 2896 64704
rect 3003 63884 3069 63885
rect 3003 63820 3004 63884
rect 3068 63820 3069 63884
rect 3003 63819 3069 63820
rect 2576 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2267 62932 2333 62933
rect 2267 62868 2268 62932
rect 2332 62868 2333 62932
rect 2267 62867 2333 62868
rect 2576 62592 2896 63616
rect 2576 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2576 61504 2896 62528
rect 2576 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2267 61164 2333 61165
rect 2267 61100 2268 61164
rect 2332 61100 2333 61164
rect 2267 61099 2333 61100
rect 2270 60485 2330 61099
rect 2267 60484 2333 60485
rect 2267 60420 2268 60484
rect 2332 60420 2333 60484
rect 2267 60419 2333 60420
rect 2576 60416 2896 61440
rect 2576 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2267 60348 2333 60349
rect 2267 60284 2268 60348
rect 2332 60284 2333 60348
rect 2267 60283 2333 60284
rect 2083 60212 2149 60213
rect 2083 60148 2084 60212
rect 2148 60148 2149 60212
rect 2083 60147 2149 60148
rect 2083 60076 2149 60077
rect 2083 60012 2084 60076
rect 2148 60012 2149 60076
rect 2083 60011 2149 60012
rect 2086 58037 2146 60011
rect 2083 58036 2149 58037
rect 2083 57972 2084 58036
rect 2148 57972 2149 58036
rect 2083 57971 2149 57972
rect 2083 57628 2149 57629
rect 2083 57564 2084 57628
rect 2148 57564 2149 57628
rect 2083 57563 2149 57564
rect 2086 56541 2146 57563
rect 2270 56677 2330 60283
rect 2576 59328 2896 60352
rect 2576 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2576 58240 2896 59264
rect 2576 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2576 57152 2896 58176
rect 2576 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2267 56676 2333 56677
rect 2267 56612 2268 56676
rect 2332 56612 2333 56676
rect 2267 56611 2333 56612
rect 2083 56540 2149 56541
rect 2083 56476 2084 56540
rect 2148 56476 2149 56540
rect 2083 56475 2149 56476
rect 1899 55588 1965 55589
rect 1899 55524 1900 55588
rect 1964 55524 1965 55588
rect 1899 55523 1965 55524
rect 2086 54909 2146 56475
rect 2576 56064 2896 57088
rect 3006 56405 3066 63819
rect 3187 61708 3253 61709
rect 3187 61644 3188 61708
rect 3252 61644 3253 61708
rect 3187 61643 3253 61644
rect 3190 60893 3250 61643
rect 3187 60892 3253 60893
rect 3187 60828 3188 60892
rect 3252 60828 3253 60892
rect 3187 60827 3253 60828
rect 3190 58445 3250 60827
rect 3371 59940 3437 59941
rect 3371 59876 3372 59940
rect 3436 59876 3437 59940
rect 3371 59875 3437 59876
rect 3187 58444 3253 58445
rect 3187 58380 3188 58444
rect 3252 58380 3253 58444
rect 3187 58379 3253 58380
rect 3187 57628 3253 57629
rect 3187 57564 3188 57628
rect 3252 57564 3253 57628
rect 3187 57563 3253 57564
rect 3003 56404 3069 56405
rect 3003 56340 3004 56404
rect 3068 56340 3069 56404
rect 3003 56339 3069 56340
rect 2576 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2267 55316 2333 55317
rect 2267 55252 2268 55316
rect 2332 55252 2333 55316
rect 2267 55251 2333 55252
rect 1899 54908 1965 54909
rect 1899 54844 1900 54908
rect 1964 54844 1965 54908
rect 1899 54843 1965 54844
rect 2083 54908 2149 54909
rect 2083 54844 2084 54908
rect 2148 54844 2149 54908
rect 2083 54843 2149 54844
rect 1902 51373 1962 54843
rect 2270 54770 2330 55251
rect 2086 54710 2330 54770
rect 2576 54976 2896 56000
rect 2576 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2086 53141 2146 54710
rect 2267 54500 2333 54501
rect 2267 54436 2268 54500
rect 2332 54436 2333 54500
rect 2267 54435 2333 54436
rect 2083 53140 2149 53141
rect 2083 53076 2084 53140
rect 2148 53076 2149 53140
rect 2083 53075 2149 53076
rect 2086 52053 2146 53075
rect 2270 52730 2330 54435
rect 2576 53888 2896 54912
rect 3190 54501 3250 57563
rect 3187 54500 3253 54501
rect 3187 54436 3188 54500
rect 3252 54436 3253 54500
rect 3187 54435 3253 54436
rect 3187 54092 3253 54093
rect 3187 54028 3188 54092
rect 3252 54028 3253 54092
rect 3187 54027 3253 54028
rect 2576 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2576 52800 2896 53824
rect 2576 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2270 52670 2514 52730
rect 2267 52188 2333 52189
rect 2267 52124 2268 52188
rect 2332 52124 2333 52188
rect 2267 52123 2333 52124
rect 2083 52052 2149 52053
rect 2083 51988 2084 52052
rect 2148 51988 2149 52052
rect 2083 51987 2149 51988
rect 2083 51916 2149 51917
rect 2083 51852 2084 51916
rect 2148 51852 2149 51916
rect 2083 51851 2149 51852
rect 1899 51372 1965 51373
rect 1899 51308 1900 51372
rect 1964 51308 1965 51372
rect 1899 51307 1965 51308
rect 1899 51236 1965 51237
rect 1899 51172 1900 51236
rect 1964 51172 1965 51236
rect 1899 51171 1965 51172
rect 1715 49604 1781 49605
rect 1715 49540 1716 49604
rect 1780 49540 1781 49604
rect 1715 49539 1781 49540
rect 1715 49196 1781 49197
rect 1715 49132 1716 49196
rect 1780 49132 1781 49196
rect 1715 49131 1781 49132
rect 1531 48516 1597 48517
rect 1531 48452 1532 48516
rect 1596 48452 1597 48516
rect 1531 48451 1597 48452
rect 1347 48108 1413 48109
rect 1347 48044 1348 48108
rect 1412 48044 1413 48108
rect 1347 48043 1413 48044
rect 1531 47972 1597 47973
rect 1531 47908 1532 47972
rect 1596 47908 1597 47972
rect 1531 47907 1597 47908
rect 1534 46749 1594 47907
rect 1531 46748 1597 46749
rect 1531 46684 1532 46748
rect 1596 46684 1597 46748
rect 1531 46683 1597 46684
rect 1718 45525 1778 49131
rect 1902 48517 1962 51171
rect 1899 48516 1965 48517
rect 1899 48452 1900 48516
rect 1964 48452 1965 48516
rect 1899 48451 1965 48452
rect 1899 48108 1965 48109
rect 1899 48044 1900 48108
rect 1964 48044 1965 48108
rect 1899 48043 1965 48044
rect 1347 45524 1413 45525
rect 1347 45460 1348 45524
rect 1412 45460 1413 45524
rect 1347 45459 1413 45460
rect 1715 45524 1781 45525
rect 1715 45460 1716 45524
rect 1780 45460 1781 45524
rect 1715 45459 1781 45460
rect 1350 30565 1410 45459
rect 1531 44572 1597 44573
rect 1531 44508 1532 44572
rect 1596 44508 1597 44572
rect 1531 44507 1597 44508
rect 1534 40901 1594 44507
rect 1715 43484 1781 43485
rect 1715 43420 1716 43484
rect 1780 43420 1781 43484
rect 1715 43419 1781 43420
rect 1531 40900 1597 40901
rect 1531 40836 1532 40900
rect 1596 40836 1597 40900
rect 1718 40898 1778 43419
rect 1902 42533 1962 48043
rect 1899 42532 1965 42533
rect 1899 42468 1900 42532
rect 1964 42468 1965 42532
rect 1899 42467 1965 42468
rect 1899 42124 1965 42125
rect 1899 42060 1900 42124
rect 1964 42060 1965 42124
rect 1899 42059 1965 42060
rect 1902 41173 1962 42059
rect 1899 41172 1965 41173
rect 1899 41108 1900 41172
rect 1964 41108 1965 41172
rect 1899 41107 1965 41108
rect 1718 40838 1962 40898
rect 1531 40835 1597 40836
rect 1715 40764 1781 40765
rect 1715 40700 1716 40764
rect 1780 40700 1781 40764
rect 1715 40699 1781 40700
rect 1531 37772 1597 37773
rect 1531 37708 1532 37772
rect 1596 37708 1597 37772
rect 1531 37707 1597 37708
rect 1534 30701 1594 37707
rect 1718 34917 1778 40699
rect 1902 38181 1962 40838
rect 1899 38180 1965 38181
rect 1899 38116 1900 38180
rect 1964 38116 1965 38180
rect 1899 38115 1965 38116
rect 1715 34916 1781 34917
rect 1715 34852 1716 34916
rect 1780 34852 1781 34916
rect 1715 34851 1781 34852
rect 1899 32196 1965 32197
rect 1899 32132 1900 32196
rect 1964 32132 1965 32196
rect 1899 32131 1965 32132
rect 1902 31381 1962 32131
rect 1899 31380 1965 31381
rect 1899 31316 1900 31380
rect 1964 31316 1965 31380
rect 1899 31315 1965 31316
rect 1531 30700 1597 30701
rect 1531 30636 1532 30700
rect 1596 30636 1597 30700
rect 1531 30635 1597 30636
rect 1347 30564 1413 30565
rect 1347 30500 1348 30564
rect 1412 30500 1413 30564
rect 1347 30499 1413 30500
rect 1163 30292 1229 30293
rect 1163 30228 1164 30292
rect 1228 30228 1229 30292
rect 1163 30227 1229 30228
rect 1531 30020 1597 30021
rect 1531 29956 1532 30020
rect 1596 29956 1597 30020
rect 1531 29955 1597 29956
rect 1534 28117 1594 29955
rect 2086 29885 2146 51851
rect 2270 50965 2330 52123
rect 2267 50964 2333 50965
rect 2267 50900 2268 50964
rect 2332 50900 2333 50964
rect 2267 50899 2333 50900
rect 2267 50012 2333 50013
rect 2267 49948 2268 50012
rect 2332 49948 2333 50012
rect 2267 49947 2333 49948
rect 2270 42397 2330 49947
rect 2267 42396 2333 42397
rect 2267 42332 2268 42396
rect 2332 42332 2333 42396
rect 2267 42331 2333 42332
rect 2454 41430 2514 52670
rect 2270 41370 2514 41430
rect 2576 51712 2896 52736
rect 2576 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2576 50624 2896 51648
rect 3003 51508 3069 51509
rect 3003 51444 3004 51508
rect 3068 51444 3069 51508
rect 3003 51443 3069 51444
rect 2576 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2576 49536 2896 50560
rect 2576 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2576 48448 2896 49472
rect 2576 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2576 47360 2896 48384
rect 2576 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2576 46272 2896 47296
rect 3006 46885 3066 51443
rect 3190 47157 3250 54027
rect 3374 49194 3434 59875
rect 3558 59261 3618 65043
rect 3555 59260 3621 59261
rect 3555 59196 3556 59260
rect 3620 59196 3621 59260
rect 3555 59195 3621 59196
rect 3555 59124 3621 59125
rect 3555 59060 3556 59124
rect 3620 59060 3621 59124
rect 3555 59059 3621 59060
rect 3558 49197 3618 59059
rect 3742 58037 3802 65995
rect 4208 65312 4528 66336
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 64224 4528 65248
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 63136 4528 64160
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 62048 4528 63072
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 60960 4528 61984
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 3923 60892 3989 60893
rect 3923 60828 3924 60892
rect 3988 60828 3989 60892
rect 3923 60827 3989 60828
rect 3926 60621 3986 60827
rect 3923 60620 3989 60621
rect 3923 60556 3924 60620
rect 3988 60556 3989 60620
rect 3923 60555 3989 60556
rect 4208 59872 4528 60896
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 58784 4528 59808
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 3739 58036 3805 58037
rect 3739 57972 3740 58036
rect 3804 57972 3805 58036
rect 3739 57971 3805 57972
rect 3739 57764 3805 57765
rect 3739 57700 3740 57764
rect 3804 57700 3805 57764
rect 3739 57699 3805 57700
rect 3742 54090 3802 57699
rect 4208 57696 4528 58720
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 56608 4528 57632
rect 5840 77824 6160 77840
rect 5840 77760 5848 77824
rect 5912 77760 5928 77824
rect 5992 77760 6008 77824
rect 6072 77760 6088 77824
rect 6152 77760 6160 77824
rect 5840 76736 6160 77760
rect 5840 76672 5848 76736
rect 5912 76672 5928 76736
rect 5992 76672 6008 76736
rect 6072 76672 6088 76736
rect 6152 76672 6160 76736
rect 5840 75648 6160 76672
rect 5840 75584 5848 75648
rect 5912 75584 5928 75648
rect 5992 75584 6008 75648
rect 6072 75584 6088 75648
rect 6152 75584 6160 75648
rect 5840 74560 6160 75584
rect 5840 74496 5848 74560
rect 5912 74496 5928 74560
rect 5992 74496 6008 74560
rect 6072 74496 6088 74560
rect 6152 74496 6160 74560
rect 5840 73472 6160 74496
rect 5840 73408 5848 73472
rect 5912 73408 5928 73472
rect 5992 73408 6008 73472
rect 6072 73408 6088 73472
rect 6152 73408 6160 73472
rect 5840 72384 6160 73408
rect 5840 72320 5848 72384
rect 5912 72320 5928 72384
rect 5992 72320 6008 72384
rect 6072 72320 6088 72384
rect 6152 72320 6160 72384
rect 5840 71296 6160 72320
rect 5840 71232 5848 71296
rect 5912 71232 5928 71296
rect 5992 71232 6008 71296
rect 6072 71232 6088 71296
rect 6152 71232 6160 71296
rect 5840 70208 6160 71232
rect 5840 70144 5848 70208
rect 5912 70144 5928 70208
rect 5992 70144 6008 70208
rect 6072 70144 6088 70208
rect 6152 70144 6160 70208
rect 5840 69120 6160 70144
rect 5840 69056 5848 69120
rect 5912 69056 5928 69120
rect 5992 69056 6008 69120
rect 6072 69056 6088 69120
rect 6152 69056 6160 69120
rect 5840 68032 6160 69056
rect 5840 67968 5848 68032
rect 5912 67968 5928 68032
rect 5992 67968 6008 68032
rect 6072 67968 6088 68032
rect 6152 67968 6160 68032
rect 5840 66944 6160 67968
rect 5840 66880 5848 66944
rect 5912 66880 5928 66944
rect 5992 66880 6008 66944
rect 6072 66880 6088 66944
rect 6152 66880 6160 66944
rect 5840 65856 6160 66880
rect 5840 65792 5848 65856
rect 5912 65792 5928 65856
rect 5992 65792 6008 65856
rect 6072 65792 6088 65856
rect 6152 65792 6160 65856
rect 5840 64768 6160 65792
rect 5840 64704 5848 64768
rect 5912 64704 5928 64768
rect 5992 64704 6008 64768
rect 6072 64704 6088 64768
rect 6152 64704 6160 64768
rect 5840 63680 6160 64704
rect 5840 63616 5848 63680
rect 5912 63616 5928 63680
rect 5992 63616 6008 63680
rect 6072 63616 6088 63680
rect 6152 63616 6160 63680
rect 5840 62592 6160 63616
rect 5840 62528 5848 62592
rect 5912 62528 5928 62592
rect 5992 62528 6008 62592
rect 6072 62528 6088 62592
rect 6152 62528 6160 62592
rect 5840 61504 6160 62528
rect 5840 61440 5848 61504
rect 5912 61440 5928 61504
rect 5992 61440 6008 61504
rect 6072 61440 6088 61504
rect 6152 61440 6160 61504
rect 5840 60416 6160 61440
rect 5840 60352 5848 60416
rect 5912 60352 5928 60416
rect 5992 60352 6008 60416
rect 6072 60352 6088 60416
rect 6152 60352 6160 60416
rect 5840 59328 6160 60352
rect 5840 59264 5848 59328
rect 5912 59264 5928 59328
rect 5992 59264 6008 59328
rect 6072 59264 6088 59328
rect 6152 59264 6160 59328
rect 5840 58240 6160 59264
rect 5840 58176 5848 58240
rect 5912 58176 5928 58240
rect 5992 58176 6008 58240
rect 6072 58176 6088 58240
rect 6152 58176 6160 58240
rect 5579 57356 5645 57357
rect 5579 57292 5580 57356
rect 5644 57292 5645 57356
rect 5579 57291 5645 57292
rect 5395 56812 5461 56813
rect 5395 56748 5396 56812
rect 5460 56748 5461 56812
rect 5395 56747 5461 56748
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 3923 55860 3989 55861
rect 3923 55796 3924 55860
rect 3988 55796 3989 55860
rect 3923 55795 3989 55796
rect 3926 54365 3986 55795
rect 4208 55520 4528 56544
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 54432 4528 55456
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 3923 54364 3989 54365
rect 3923 54300 3924 54364
rect 3988 54300 3989 54364
rect 3923 54299 3989 54300
rect 3742 54030 3986 54090
rect 3739 50420 3805 50421
rect 3739 50356 3740 50420
rect 3804 50356 3805 50420
rect 3739 50355 3805 50356
rect 3555 49196 3621 49197
rect 3374 49134 3480 49194
rect 3420 48514 3480 49134
rect 3555 49132 3556 49196
rect 3620 49132 3621 49196
rect 3555 49131 3621 49132
rect 3555 48652 3621 48653
rect 3555 48588 3556 48652
rect 3620 48588 3621 48652
rect 3555 48587 3621 48588
rect 3374 48454 3480 48514
rect 3187 47156 3253 47157
rect 3187 47092 3188 47156
rect 3252 47092 3253 47156
rect 3187 47091 3253 47092
rect 3003 46884 3069 46885
rect 3003 46820 3004 46884
rect 3068 46820 3069 46884
rect 3003 46819 3069 46820
rect 3187 46748 3253 46749
rect 3187 46684 3188 46748
rect 3252 46684 3253 46748
rect 3187 46683 3253 46684
rect 2576 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2576 45184 2896 46208
rect 3003 45524 3069 45525
rect 3003 45460 3004 45524
rect 3068 45460 3069 45524
rect 3003 45459 3069 45460
rect 2576 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2576 44096 2896 45120
rect 2576 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2576 43008 2896 44032
rect 2576 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2576 41920 2896 42944
rect 2576 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2270 40085 2330 41370
rect 2576 40832 2896 41856
rect 3006 41581 3066 45459
rect 3190 44570 3250 46683
rect 3374 44845 3434 48454
rect 3558 46749 3618 48587
rect 3555 46748 3621 46749
rect 3555 46684 3556 46748
rect 3620 46684 3621 46748
rect 3555 46683 3621 46684
rect 3555 46612 3621 46613
rect 3555 46548 3556 46612
rect 3620 46548 3621 46612
rect 3555 46547 3621 46548
rect 3371 44844 3437 44845
rect 3371 44780 3372 44844
rect 3436 44780 3437 44844
rect 3371 44779 3437 44780
rect 3190 44510 3434 44570
rect 3187 44300 3253 44301
rect 3187 44236 3188 44300
rect 3252 44236 3253 44300
rect 3187 44235 3253 44236
rect 3003 41580 3069 41581
rect 3003 41516 3004 41580
rect 3068 41516 3069 41580
rect 3003 41515 3069 41516
rect 3003 41036 3069 41037
rect 3003 40972 3004 41036
rect 3068 40972 3069 41036
rect 3003 40971 3069 40972
rect 2576 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2267 40084 2333 40085
rect 2267 40020 2268 40084
rect 2332 40020 2333 40084
rect 2267 40019 2333 40020
rect 2576 39744 2896 40768
rect 2576 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2267 39132 2333 39133
rect 2267 39068 2268 39132
rect 2332 39068 2333 39132
rect 2267 39067 2333 39068
rect 2083 29884 2149 29885
rect 2083 29820 2084 29884
rect 2148 29820 2149 29884
rect 2083 29819 2149 29820
rect 2270 29341 2330 39067
rect 2576 38656 2896 39680
rect 3006 39133 3066 40971
rect 3190 40085 3250 44235
rect 3374 43077 3434 44510
rect 3371 43076 3437 43077
rect 3371 43012 3372 43076
rect 3436 43012 3437 43076
rect 3371 43011 3437 43012
rect 3371 42804 3437 42805
rect 3371 42740 3372 42804
rect 3436 42740 3437 42804
rect 3371 42739 3437 42740
rect 3187 40084 3253 40085
rect 3187 40020 3188 40084
rect 3252 40020 3253 40084
rect 3187 40019 3253 40020
rect 3003 39132 3069 39133
rect 3003 39068 3004 39132
rect 3068 39068 3069 39132
rect 3003 39067 3069 39068
rect 3187 38996 3253 38997
rect 3187 38932 3188 38996
rect 3252 38932 3253 38996
rect 3187 38931 3253 38932
rect 3003 38860 3069 38861
rect 3003 38796 3004 38860
rect 3068 38796 3069 38860
rect 3003 38795 3069 38796
rect 2576 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2576 37568 2896 38592
rect 2576 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2576 36480 2896 37504
rect 2576 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2576 35392 2896 36416
rect 2576 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2576 34304 2896 35328
rect 2576 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2576 33216 2896 34240
rect 2576 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2576 32128 2896 33152
rect 2576 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2576 31040 2896 32064
rect 3006 31517 3066 38795
rect 3190 37909 3250 38931
rect 3187 37908 3253 37909
rect 3187 37844 3188 37908
rect 3252 37844 3253 37908
rect 3187 37843 3253 37844
rect 3190 32197 3250 37843
rect 3187 32196 3253 32197
rect 3187 32132 3188 32196
rect 3252 32132 3253 32196
rect 3187 32131 3253 32132
rect 3187 32060 3253 32061
rect 3187 31996 3188 32060
rect 3252 31996 3253 32060
rect 3187 31995 3253 31996
rect 3003 31516 3069 31517
rect 3003 31452 3004 31516
rect 3068 31452 3069 31516
rect 3003 31451 3069 31452
rect 3003 31380 3069 31381
rect 3003 31316 3004 31380
rect 3068 31316 3069 31380
rect 3003 31315 3069 31316
rect 2576 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2576 29952 2896 30976
rect 2576 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2267 29340 2333 29341
rect 2267 29276 2268 29340
rect 2332 29276 2333 29340
rect 2267 29275 2333 29276
rect 1899 28932 1965 28933
rect 1899 28868 1900 28932
rect 1964 28868 1965 28932
rect 1899 28867 1965 28868
rect 2083 28932 2149 28933
rect 2083 28868 2084 28932
rect 2148 28868 2149 28932
rect 2083 28867 2149 28868
rect 1902 28253 1962 28867
rect 1899 28252 1965 28253
rect 1899 28188 1900 28252
rect 1964 28188 1965 28252
rect 1899 28187 1965 28188
rect 1531 28116 1597 28117
rect 1531 28052 1532 28116
rect 1596 28052 1597 28116
rect 1531 28051 1597 28052
rect 2086 27981 2146 28867
rect 2576 28864 2896 29888
rect 2576 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2267 28524 2333 28525
rect 2267 28460 2268 28524
rect 2332 28460 2333 28524
rect 2267 28459 2333 28460
rect 2083 27980 2149 27981
rect 2083 27916 2084 27980
rect 2148 27916 2149 27980
rect 2083 27915 2149 27916
rect 2270 24173 2330 28459
rect 2576 27776 2896 28800
rect 3006 28661 3066 31315
rect 3003 28660 3069 28661
rect 3003 28596 3004 28660
rect 3068 28596 3069 28660
rect 3003 28595 3069 28596
rect 2576 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2576 26688 2896 27712
rect 2576 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2576 25600 2896 26624
rect 3190 26349 3250 31995
rect 3374 30429 3434 42739
rect 3558 42261 3618 46547
rect 3742 44981 3802 50355
rect 3926 49333 3986 54030
rect 4208 53344 4528 54368
rect 5211 53684 5277 53685
rect 5211 53620 5212 53684
rect 5276 53620 5277 53684
rect 5211 53619 5277 53620
rect 4659 53548 4725 53549
rect 4659 53484 4660 53548
rect 4724 53484 4725 53548
rect 4659 53483 4725 53484
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 52256 4528 53280
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 51168 4528 52192
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 50080 4528 51104
rect 4662 50829 4722 53483
rect 5027 53140 5093 53141
rect 5027 53076 5028 53140
rect 5092 53076 5093 53140
rect 5027 53075 5093 53076
rect 4843 51236 4909 51237
rect 4843 51172 4844 51236
rect 4908 51172 4909 51236
rect 4843 51171 4909 51172
rect 4846 50965 4906 51171
rect 5030 51101 5090 53075
rect 5027 51100 5093 51101
rect 5027 51036 5028 51100
rect 5092 51036 5093 51100
rect 5027 51035 5093 51036
rect 4843 50964 4909 50965
rect 4843 50900 4844 50964
rect 4908 50900 4909 50964
rect 4843 50899 4909 50900
rect 4659 50828 4725 50829
rect 4659 50764 4660 50828
rect 4724 50764 4725 50828
rect 4659 50763 4725 50764
rect 5214 50285 5274 53619
rect 5211 50284 5277 50285
rect 5211 50220 5212 50284
rect 5276 50220 5277 50284
rect 5211 50219 5277 50220
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 3923 49332 3989 49333
rect 3923 49268 3924 49332
rect 3988 49268 3989 49332
rect 3923 49267 3989 49268
rect 3923 49196 3989 49197
rect 3923 49132 3924 49196
rect 3988 49132 3989 49196
rect 3923 49131 3989 49132
rect 3739 44980 3805 44981
rect 3739 44916 3740 44980
rect 3804 44916 3805 44980
rect 3739 44915 3805 44916
rect 3739 44844 3805 44845
rect 3739 44780 3740 44844
rect 3804 44780 3805 44844
rect 3739 44779 3805 44780
rect 3555 42260 3621 42261
rect 3555 42196 3556 42260
rect 3620 42196 3621 42260
rect 3555 42195 3621 42196
rect 3555 39948 3621 39949
rect 3555 39884 3556 39948
rect 3620 39884 3621 39948
rect 3555 39883 3621 39884
rect 3558 38450 3618 39883
rect 3742 38997 3802 44779
rect 3739 38996 3805 38997
rect 3739 38932 3740 38996
rect 3804 38932 3805 38996
rect 3739 38931 3805 38932
rect 3558 38390 3802 38450
rect 3555 33012 3621 33013
rect 3555 32948 3556 33012
rect 3620 32948 3621 33012
rect 3555 32947 3621 32948
rect 3371 30428 3437 30429
rect 3371 30364 3372 30428
rect 3436 30364 3437 30428
rect 3371 30363 3437 30364
rect 3558 27981 3618 32947
rect 3742 32197 3802 38390
rect 3739 32196 3805 32197
rect 3739 32132 3740 32196
rect 3804 32132 3805 32196
rect 3739 32131 3805 32132
rect 3739 32060 3805 32061
rect 3739 31996 3740 32060
rect 3804 31996 3805 32060
rect 3739 31995 3805 31996
rect 3742 31517 3802 31995
rect 3739 31516 3805 31517
rect 3739 31452 3740 31516
rect 3804 31452 3805 31516
rect 3739 31451 3805 31452
rect 3739 30972 3805 30973
rect 3739 30908 3740 30972
rect 3804 30908 3805 30972
rect 3739 30907 3805 30908
rect 3555 27980 3621 27981
rect 3555 27916 3556 27980
rect 3620 27916 3621 27980
rect 3555 27915 3621 27916
rect 3187 26348 3253 26349
rect 3187 26284 3188 26348
rect 3252 26284 3253 26348
rect 3187 26283 3253 26284
rect 3558 25805 3618 27915
rect 3742 27437 3802 30907
rect 3739 27436 3805 27437
rect 3739 27372 3740 27436
rect 3804 27372 3805 27436
rect 3739 27371 3805 27372
rect 3555 25804 3621 25805
rect 3555 25740 3556 25804
rect 3620 25740 3621 25804
rect 3555 25739 3621 25740
rect 2576 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2576 24512 2896 25536
rect 2576 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2267 24172 2333 24173
rect 2267 24108 2268 24172
rect 2332 24108 2333 24172
rect 2267 24107 2333 24108
rect 2576 23424 2896 24448
rect 2576 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2576 22336 2896 23360
rect 2576 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2576 21248 2896 22272
rect 2576 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2576 20160 2896 21184
rect 2576 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2576 19072 2896 20096
rect 2576 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2576 17984 2896 19008
rect 2576 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2576 16896 2896 17920
rect 3003 17100 3069 17101
rect 3003 17036 3004 17100
rect 3068 17036 3069 17100
rect 3003 17035 3069 17036
rect 2576 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2576 15808 2896 16832
rect 2576 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2576 14720 2896 15744
rect 2576 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2576 13632 2896 14656
rect 2576 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2576 12544 2896 13568
rect 2576 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2576 11456 2896 12480
rect 3006 11797 3066 17035
rect 3371 15740 3437 15741
rect 3371 15676 3372 15740
rect 3436 15676 3437 15740
rect 3371 15675 3437 15676
rect 3003 11796 3069 11797
rect 3003 11732 3004 11796
rect 3068 11732 3069 11796
rect 3003 11731 3069 11732
rect 3374 11525 3434 15675
rect 3555 14108 3621 14109
rect 3555 14044 3556 14108
rect 3620 14044 3621 14108
rect 3555 14043 3621 14044
rect 3558 12477 3618 14043
rect 3555 12476 3621 12477
rect 3555 12412 3556 12476
rect 3620 12412 3621 12476
rect 3555 12411 3621 12412
rect 3371 11524 3437 11525
rect 3371 11460 3372 11524
rect 3436 11460 3437 11524
rect 3371 11459 3437 11460
rect 2576 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2576 10368 2896 11392
rect 2576 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2576 9280 2896 10304
rect 3926 10301 3986 49131
rect 4208 48992 4528 50016
rect 4659 49468 4725 49469
rect 4659 49404 4660 49468
rect 4724 49404 4725 49468
rect 4659 49403 4725 49404
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 47904 4528 48928
rect 4662 48381 4722 49403
rect 5211 49196 5277 49197
rect 5211 49132 5212 49196
rect 5276 49132 5277 49196
rect 5211 49131 5277 49132
rect 4659 48380 4725 48381
rect 4659 48316 4660 48380
rect 4724 48316 4725 48380
rect 4659 48315 4725 48316
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 46816 4528 47840
rect 4659 47020 4725 47021
rect 4659 46956 4660 47020
rect 4724 46956 4725 47020
rect 4659 46955 4725 46956
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4662 42805 4722 46955
rect 5027 46476 5093 46477
rect 5027 46412 5028 46476
rect 5092 46412 5093 46476
rect 5027 46411 5093 46412
rect 4843 45796 4909 45797
rect 4843 45732 4844 45796
rect 4908 45732 4909 45796
rect 4843 45731 4909 45732
rect 4659 42804 4725 42805
rect 4659 42740 4660 42804
rect 4724 42740 4725 42804
rect 4659 42739 4725 42740
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4659 41580 4725 41581
rect 4659 41516 4660 41580
rect 4724 41516 4725 41580
rect 4659 41515 4725 41516
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4662 37365 4722 41515
rect 4659 37364 4725 37365
rect 4659 37300 4660 37364
rect 4724 37300 4725 37364
rect 4659 37299 4725 37300
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4659 36820 4725 36821
rect 4659 36756 4660 36820
rect 4724 36756 4725 36820
rect 4659 36755 4725 36756
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 3923 10300 3989 10301
rect 3923 10236 3924 10300
rect 3988 10236 3989 10300
rect 3923 10235 3989 10236
rect 2576 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2576 8192 2896 9216
rect 2576 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2576 7104 2896 8128
rect 2576 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2576 6016 2896 7040
rect 2576 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2576 4928 2896 5952
rect 2576 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2576 3840 2896 4864
rect 2576 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2576 2752 2896 3776
rect 2576 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2576 2128 2896 2688
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4662 5949 4722 36755
rect 4659 5948 4725 5949
rect 4659 5884 4660 5948
rect 4724 5884 4725 5948
rect 4659 5883 4725 5884
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4846 5269 4906 45731
rect 5030 6765 5090 46411
rect 5214 42125 5274 49131
rect 5398 48109 5458 56747
rect 5395 48108 5461 48109
rect 5395 48044 5396 48108
rect 5460 48044 5461 48108
rect 5395 48043 5461 48044
rect 5395 47564 5461 47565
rect 5395 47500 5396 47564
rect 5460 47500 5461 47564
rect 5395 47499 5461 47500
rect 5211 42124 5277 42125
rect 5211 42060 5212 42124
rect 5276 42060 5277 42124
rect 5211 42059 5277 42060
rect 5211 41988 5277 41989
rect 5211 41924 5212 41988
rect 5276 41924 5277 41988
rect 5211 41923 5277 41924
rect 5214 38861 5274 41923
rect 5211 38860 5277 38861
rect 5211 38796 5212 38860
rect 5276 38796 5277 38860
rect 5211 38795 5277 38796
rect 5211 38316 5277 38317
rect 5211 38252 5212 38316
rect 5276 38252 5277 38316
rect 5211 38251 5277 38252
rect 5214 36410 5274 38251
rect 5398 36821 5458 47499
rect 5395 36820 5461 36821
rect 5395 36756 5396 36820
rect 5460 36756 5461 36820
rect 5395 36755 5461 36756
rect 5214 36350 5458 36410
rect 5211 36140 5277 36141
rect 5211 36076 5212 36140
rect 5276 36076 5277 36140
rect 5211 36075 5277 36076
rect 5214 32469 5274 36075
rect 5211 32468 5277 32469
rect 5211 32404 5212 32468
rect 5276 32404 5277 32468
rect 5211 32403 5277 32404
rect 5211 32060 5277 32061
rect 5211 31996 5212 32060
rect 5276 31996 5277 32060
rect 5211 31995 5277 31996
rect 5214 27029 5274 31995
rect 5398 31789 5458 36350
rect 5395 31788 5461 31789
rect 5395 31724 5396 31788
rect 5460 31724 5461 31788
rect 5395 31723 5461 31724
rect 5582 28117 5642 57291
rect 5840 57152 6160 58176
rect 5840 57088 5848 57152
rect 5912 57088 5928 57152
rect 5992 57088 6008 57152
rect 6072 57088 6088 57152
rect 6152 57088 6160 57152
rect 5840 56064 6160 57088
rect 5840 56000 5848 56064
rect 5912 56000 5928 56064
rect 5992 56000 6008 56064
rect 6072 56000 6088 56064
rect 6152 56000 6160 56064
rect 5840 54976 6160 56000
rect 7472 77280 7792 77840
rect 7472 77216 7480 77280
rect 7544 77216 7560 77280
rect 7624 77216 7640 77280
rect 7704 77216 7720 77280
rect 7784 77216 7792 77280
rect 7472 76192 7792 77216
rect 7472 76128 7480 76192
rect 7544 76128 7560 76192
rect 7624 76128 7640 76192
rect 7704 76128 7720 76192
rect 7784 76128 7792 76192
rect 7472 75104 7792 76128
rect 7472 75040 7480 75104
rect 7544 75040 7560 75104
rect 7624 75040 7640 75104
rect 7704 75040 7720 75104
rect 7784 75040 7792 75104
rect 7472 74016 7792 75040
rect 7472 73952 7480 74016
rect 7544 73952 7560 74016
rect 7624 73952 7640 74016
rect 7704 73952 7720 74016
rect 7784 73952 7792 74016
rect 7472 72928 7792 73952
rect 7472 72864 7480 72928
rect 7544 72864 7560 72928
rect 7624 72864 7640 72928
rect 7704 72864 7720 72928
rect 7784 72864 7792 72928
rect 7472 71840 7792 72864
rect 7472 71776 7480 71840
rect 7544 71776 7560 71840
rect 7624 71776 7640 71840
rect 7704 71776 7720 71840
rect 7784 71776 7792 71840
rect 7472 70752 7792 71776
rect 7472 70688 7480 70752
rect 7544 70688 7560 70752
rect 7624 70688 7640 70752
rect 7704 70688 7720 70752
rect 7784 70688 7792 70752
rect 7472 69664 7792 70688
rect 7472 69600 7480 69664
rect 7544 69600 7560 69664
rect 7624 69600 7640 69664
rect 7704 69600 7720 69664
rect 7784 69600 7792 69664
rect 7472 68576 7792 69600
rect 7472 68512 7480 68576
rect 7544 68512 7560 68576
rect 7624 68512 7640 68576
rect 7704 68512 7720 68576
rect 7784 68512 7792 68576
rect 7472 67488 7792 68512
rect 7472 67424 7480 67488
rect 7544 67424 7560 67488
rect 7624 67424 7640 67488
rect 7704 67424 7720 67488
rect 7784 67424 7792 67488
rect 7472 66400 7792 67424
rect 7472 66336 7480 66400
rect 7544 66336 7560 66400
rect 7624 66336 7640 66400
rect 7704 66336 7720 66400
rect 7784 66336 7792 66400
rect 7472 65312 7792 66336
rect 7472 65248 7480 65312
rect 7544 65248 7560 65312
rect 7624 65248 7640 65312
rect 7704 65248 7720 65312
rect 7784 65248 7792 65312
rect 7472 64224 7792 65248
rect 7472 64160 7480 64224
rect 7544 64160 7560 64224
rect 7624 64160 7640 64224
rect 7704 64160 7720 64224
rect 7784 64160 7792 64224
rect 7472 63136 7792 64160
rect 7472 63072 7480 63136
rect 7544 63072 7560 63136
rect 7624 63072 7640 63136
rect 7704 63072 7720 63136
rect 7784 63072 7792 63136
rect 7472 62048 7792 63072
rect 7472 61984 7480 62048
rect 7544 61984 7560 62048
rect 7624 61984 7640 62048
rect 7704 61984 7720 62048
rect 7784 61984 7792 62048
rect 7472 60960 7792 61984
rect 7472 60896 7480 60960
rect 7544 60896 7560 60960
rect 7624 60896 7640 60960
rect 7704 60896 7720 60960
rect 7784 60896 7792 60960
rect 7472 59872 7792 60896
rect 7472 59808 7480 59872
rect 7544 59808 7560 59872
rect 7624 59808 7640 59872
rect 7704 59808 7720 59872
rect 7784 59808 7792 59872
rect 7472 58784 7792 59808
rect 7472 58720 7480 58784
rect 7544 58720 7560 58784
rect 7624 58720 7640 58784
rect 7704 58720 7720 58784
rect 7784 58720 7792 58784
rect 7472 57696 7792 58720
rect 7472 57632 7480 57696
rect 7544 57632 7560 57696
rect 7624 57632 7640 57696
rect 7704 57632 7720 57696
rect 7784 57632 7792 57696
rect 7472 56608 7792 57632
rect 7472 56544 7480 56608
rect 7544 56544 7560 56608
rect 7624 56544 7640 56608
rect 7704 56544 7720 56608
rect 7784 56544 7792 56608
rect 7472 55520 7792 56544
rect 7472 55456 7480 55520
rect 7544 55456 7560 55520
rect 7624 55456 7640 55520
rect 7704 55456 7720 55520
rect 7784 55456 7792 55520
rect 6315 55316 6381 55317
rect 6315 55252 6316 55316
rect 6380 55252 6381 55316
rect 6315 55251 6381 55252
rect 5840 54912 5848 54976
rect 5912 54912 5928 54976
rect 5992 54912 6008 54976
rect 6072 54912 6088 54976
rect 6152 54912 6160 54976
rect 5840 53888 6160 54912
rect 5840 53824 5848 53888
rect 5912 53824 5928 53888
rect 5992 53824 6008 53888
rect 6072 53824 6088 53888
rect 6152 53824 6160 53888
rect 5840 52800 6160 53824
rect 5840 52736 5848 52800
rect 5912 52736 5928 52800
rect 5992 52736 6008 52800
rect 6072 52736 6088 52800
rect 6152 52736 6160 52800
rect 5840 51712 6160 52736
rect 5840 51648 5848 51712
rect 5912 51648 5928 51712
rect 5992 51648 6008 51712
rect 6072 51648 6088 51712
rect 6152 51648 6160 51712
rect 5840 50624 6160 51648
rect 5840 50560 5848 50624
rect 5912 50560 5928 50624
rect 5992 50560 6008 50624
rect 6072 50560 6088 50624
rect 6152 50560 6160 50624
rect 5840 49536 6160 50560
rect 5840 49472 5848 49536
rect 5912 49472 5928 49536
rect 5992 49472 6008 49536
rect 6072 49472 6088 49536
rect 6152 49472 6160 49536
rect 5840 48448 6160 49472
rect 5840 48384 5848 48448
rect 5912 48384 5928 48448
rect 5992 48384 6008 48448
rect 6072 48384 6088 48448
rect 6152 48384 6160 48448
rect 5840 47360 6160 48384
rect 5840 47296 5848 47360
rect 5912 47296 5928 47360
rect 5992 47296 6008 47360
rect 6072 47296 6088 47360
rect 6152 47296 6160 47360
rect 5840 46272 6160 47296
rect 5840 46208 5848 46272
rect 5912 46208 5928 46272
rect 5992 46208 6008 46272
rect 6072 46208 6088 46272
rect 6152 46208 6160 46272
rect 5840 45184 6160 46208
rect 5840 45120 5848 45184
rect 5912 45120 5928 45184
rect 5992 45120 6008 45184
rect 6072 45120 6088 45184
rect 6152 45120 6160 45184
rect 5840 44096 6160 45120
rect 5840 44032 5848 44096
rect 5912 44032 5928 44096
rect 5992 44032 6008 44096
rect 6072 44032 6088 44096
rect 6152 44032 6160 44096
rect 5840 43008 6160 44032
rect 5840 42944 5848 43008
rect 5912 42944 5928 43008
rect 5992 42944 6008 43008
rect 6072 42944 6088 43008
rect 6152 42944 6160 43008
rect 5840 41920 6160 42944
rect 5840 41856 5848 41920
rect 5912 41856 5928 41920
rect 5992 41856 6008 41920
rect 6072 41856 6088 41920
rect 6152 41856 6160 41920
rect 5840 40832 6160 41856
rect 5840 40768 5848 40832
rect 5912 40768 5928 40832
rect 5992 40768 6008 40832
rect 6072 40768 6088 40832
rect 6152 40768 6160 40832
rect 5840 39744 6160 40768
rect 5840 39680 5848 39744
rect 5912 39680 5928 39744
rect 5992 39680 6008 39744
rect 6072 39680 6088 39744
rect 6152 39680 6160 39744
rect 5840 38656 6160 39680
rect 5840 38592 5848 38656
rect 5912 38592 5928 38656
rect 5992 38592 6008 38656
rect 6072 38592 6088 38656
rect 6152 38592 6160 38656
rect 5840 37568 6160 38592
rect 5840 37504 5848 37568
rect 5912 37504 5928 37568
rect 5992 37504 6008 37568
rect 6072 37504 6088 37568
rect 6152 37504 6160 37568
rect 5840 36480 6160 37504
rect 5840 36416 5848 36480
rect 5912 36416 5928 36480
rect 5992 36416 6008 36480
rect 6072 36416 6088 36480
rect 6152 36416 6160 36480
rect 5840 35392 6160 36416
rect 5840 35328 5848 35392
rect 5912 35328 5928 35392
rect 5992 35328 6008 35392
rect 6072 35328 6088 35392
rect 6152 35328 6160 35392
rect 5840 34304 6160 35328
rect 5840 34240 5848 34304
rect 5912 34240 5928 34304
rect 5992 34240 6008 34304
rect 6072 34240 6088 34304
rect 6152 34240 6160 34304
rect 5840 33216 6160 34240
rect 5840 33152 5848 33216
rect 5912 33152 5928 33216
rect 5992 33152 6008 33216
rect 6072 33152 6088 33216
rect 6152 33152 6160 33216
rect 5840 32128 6160 33152
rect 5840 32064 5848 32128
rect 5912 32064 5928 32128
rect 5992 32064 6008 32128
rect 6072 32064 6088 32128
rect 6152 32064 6160 32128
rect 5840 31040 6160 32064
rect 5840 30976 5848 31040
rect 5912 30976 5928 31040
rect 5992 30976 6008 31040
rect 6072 30976 6088 31040
rect 6152 30976 6160 31040
rect 5840 29952 6160 30976
rect 5840 29888 5848 29952
rect 5912 29888 5928 29952
rect 5992 29888 6008 29952
rect 6072 29888 6088 29952
rect 6152 29888 6160 29952
rect 5840 28864 6160 29888
rect 5840 28800 5848 28864
rect 5912 28800 5928 28864
rect 5992 28800 6008 28864
rect 6072 28800 6088 28864
rect 6152 28800 6160 28864
rect 5579 28116 5645 28117
rect 5579 28052 5580 28116
rect 5644 28052 5645 28116
rect 5579 28051 5645 28052
rect 5840 27776 6160 28800
rect 5840 27712 5848 27776
rect 5912 27712 5928 27776
rect 5992 27712 6008 27776
rect 6072 27712 6088 27776
rect 6152 27712 6160 27776
rect 5211 27028 5277 27029
rect 5211 26964 5212 27028
rect 5276 26964 5277 27028
rect 5211 26963 5277 26964
rect 5840 26688 6160 27712
rect 6318 26893 6378 55251
rect 7472 54432 7792 55456
rect 7472 54368 7480 54432
rect 7544 54368 7560 54432
rect 7624 54368 7640 54432
rect 7704 54368 7720 54432
rect 7784 54368 7792 54432
rect 7472 53344 7792 54368
rect 7472 53280 7480 53344
rect 7544 53280 7560 53344
rect 7624 53280 7640 53344
rect 7704 53280 7720 53344
rect 7784 53280 7792 53344
rect 7472 52256 7792 53280
rect 7472 52192 7480 52256
rect 7544 52192 7560 52256
rect 7624 52192 7640 52256
rect 7704 52192 7720 52256
rect 7784 52192 7792 52256
rect 7472 51168 7792 52192
rect 7472 51104 7480 51168
rect 7544 51104 7560 51168
rect 7624 51104 7640 51168
rect 7704 51104 7720 51168
rect 7784 51104 7792 51168
rect 7472 50080 7792 51104
rect 7472 50016 7480 50080
rect 7544 50016 7560 50080
rect 7624 50016 7640 50080
rect 7704 50016 7720 50080
rect 7784 50016 7792 50080
rect 7472 48992 7792 50016
rect 7472 48928 7480 48992
rect 7544 48928 7560 48992
rect 7624 48928 7640 48992
rect 7704 48928 7720 48992
rect 7784 48928 7792 48992
rect 7472 47904 7792 48928
rect 7472 47840 7480 47904
rect 7544 47840 7560 47904
rect 7624 47840 7640 47904
rect 7704 47840 7720 47904
rect 7784 47840 7792 47904
rect 7472 46816 7792 47840
rect 7472 46752 7480 46816
rect 7544 46752 7560 46816
rect 7624 46752 7640 46816
rect 7704 46752 7720 46816
rect 7784 46752 7792 46816
rect 7472 45728 7792 46752
rect 7472 45664 7480 45728
rect 7544 45664 7560 45728
rect 7624 45664 7640 45728
rect 7704 45664 7720 45728
rect 7784 45664 7792 45728
rect 7472 44640 7792 45664
rect 7472 44576 7480 44640
rect 7544 44576 7560 44640
rect 7624 44576 7640 44640
rect 7704 44576 7720 44640
rect 7784 44576 7792 44640
rect 7472 43552 7792 44576
rect 7472 43488 7480 43552
rect 7544 43488 7560 43552
rect 7624 43488 7640 43552
rect 7704 43488 7720 43552
rect 7784 43488 7792 43552
rect 7472 42464 7792 43488
rect 7472 42400 7480 42464
rect 7544 42400 7560 42464
rect 7624 42400 7640 42464
rect 7704 42400 7720 42464
rect 7784 42400 7792 42464
rect 7472 41376 7792 42400
rect 7472 41312 7480 41376
rect 7544 41312 7560 41376
rect 7624 41312 7640 41376
rect 7704 41312 7720 41376
rect 7784 41312 7792 41376
rect 7472 40288 7792 41312
rect 7472 40224 7480 40288
rect 7544 40224 7560 40288
rect 7624 40224 7640 40288
rect 7704 40224 7720 40288
rect 7784 40224 7792 40288
rect 7472 39200 7792 40224
rect 7472 39136 7480 39200
rect 7544 39136 7560 39200
rect 7624 39136 7640 39200
rect 7704 39136 7720 39200
rect 7784 39136 7792 39200
rect 7472 38112 7792 39136
rect 7472 38048 7480 38112
rect 7544 38048 7560 38112
rect 7624 38048 7640 38112
rect 7704 38048 7720 38112
rect 7784 38048 7792 38112
rect 7472 37024 7792 38048
rect 7472 36960 7480 37024
rect 7544 36960 7560 37024
rect 7624 36960 7640 37024
rect 7704 36960 7720 37024
rect 7784 36960 7792 37024
rect 7472 35936 7792 36960
rect 7472 35872 7480 35936
rect 7544 35872 7560 35936
rect 7624 35872 7640 35936
rect 7704 35872 7720 35936
rect 7784 35872 7792 35936
rect 7472 34848 7792 35872
rect 7472 34784 7480 34848
rect 7544 34784 7560 34848
rect 7624 34784 7640 34848
rect 7704 34784 7720 34848
rect 7784 34784 7792 34848
rect 7472 33760 7792 34784
rect 7472 33696 7480 33760
rect 7544 33696 7560 33760
rect 7624 33696 7640 33760
rect 7704 33696 7720 33760
rect 7784 33696 7792 33760
rect 7472 32672 7792 33696
rect 7472 32608 7480 32672
rect 7544 32608 7560 32672
rect 7624 32608 7640 32672
rect 7704 32608 7720 32672
rect 7784 32608 7792 32672
rect 7472 31584 7792 32608
rect 7472 31520 7480 31584
rect 7544 31520 7560 31584
rect 7624 31520 7640 31584
rect 7704 31520 7720 31584
rect 7784 31520 7792 31584
rect 7472 30496 7792 31520
rect 7472 30432 7480 30496
rect 7544 30432 7560 30496
rect 7624 30432 7640 30496
rect 7704 30432 7720 30496
rect 7784 30432 7792 30496
rect 7472 29408 7792 30432
rect 7472 29344 7480 29408
rect 7544 29344 7560 29408
rect 7624 29344 7640 29408
rect 7704 29344 7720 29408
rect 7784 29344 7792 29408
rect 7472 28320 7792 29344
rect 7472 28256 7480 28320
rect 7544 28256 7560 28320
rect 7624 28256 7640 28320
rect 7704 28256 7720 28320
rect 7784 28256 7792 28320
rect 7472 27232 7792 28256
rect 7472 27168 7480 27232
rect 7544 27168 7560 27232
rect 7624 27168 7640 27232
rect 7704 27168 7720 27232
rect 7784 27168 7792 27232
rect 6315 26892 6381 26893
rect 6315 26828 6316 26892
rect 6380 26828 6381 26892
rect 6315 26827 6381 26828
rect 5840 26624 5848 26688
rect 5912 26624 5928 26688
rect 5992 26624 6008 26688
rect 6072 26624 6088 26688
rect 6152 26624 6160 26688
rect 5840 25600 6160 26624
rect 5840 25536 5848 25600
rect 5912 25536 5928 25600
rect 5992 25536 6008 25600
rect 6072 25536 6088 25600
rect 6152 25536 6160 25600
rect 5840 24512 6160 25536
rect 5840 24448 5848 24512
rect 5912 24448 5928 24512
rect 5992 24448 6008 24512
rect 6072 24448 6088 24512
rect 6152 24448 6160 24512
rect 5840 23424 6160 24448
rect 5840 23360 5848 23424
rect 5912 23360 5928 23424
rect 5992 23360 6008 23424
rect 6072 23360 6088 23424
rect 6152 23360 6160 23424
rect 5840 22336 6160 23360
rect 5840 22272 5848 22336
rect 5912 22272 5928 22336
rect 5992 22272 6008 22336
rect 6072 22272 6088 22336
rect 6152 22272 6160 22336
rect 5840 21248 6160 22272
rect 5840 21184 5848 21248
rect 5912 21184 5928 21248
rect 5992 21184 6008 21248
rect 6072 21184 6088 21248
rect 6152 21184 6160 21248
rect 5840 20160 6160 21184
rect 5840 20096 5848 20160
rect 5912 20096 5928 20160
rect 5992 20096 6008 20160
rect 6072 20096 6088 20160
rect 6152 20096 6160 20160
rect 5840 19072 6160 20096
rect 5840 19008 5848 19072
rect 5912 19008 5928 19072
rect 5992 19008 6008 19072
rect 6072 19008 6088 19072
rect 6152 19008 6160 19072
rect 5840 17984 6160 19008
rect 5840 17920 5848 17984
rect 5912 17920 5928 17984
rect 5992 17920 6008 17984
rect 6072 17920 6088 17984
rect 6152 17920 6160 17984
rect 5840 16896 6160 17920
rect 5840 16832 5848 16896
rect 5912 16832 5928 16896
rect 5992 16832 6008 16896
rect 6072 16832 6088 16896
rect 6152 16832 6160 16896
rect 5840 15808 6160 16832
rect 5840 15744 5848 15808
rect 5912 15744 5928 15808
rect 5992 15744 6008 15808
rect 6072 15744 6088 15808
rect 6152 15744 6160 15808
rect 5840 14720 6160 15744
rect 5840 14656 5848 14720
rect 5912 14656 5928 14720
rect 5992 14656 6008 14720
rect 6072 14656 6088 14720
rect 6152 14656 6160 14720
rect 5840 13632 6160 14656
rect 5840 13568 5848 13632
rect 5912 13568 5928 13632
rect 5992 13568 6008 13632
rect 6072 13568 6088 13632
rect 6152 13568 6160 13632
rect 5840 12544 6160 13568
rect 5840 12480 5848 12544
rect 5912 12480 5928 12544
rect 5992 12480 6008 12544
rect 6072 12480 6088 12544
rect 6152 12480 6160 12544
rect 5840 11456 6160 12480
rect 5840 11392 5848 11456
rect 5912 11392 5928 11456
rect 5992 11392 6008 11456
rect 6072 11392 6088 11456
rect 6152 11392 6160 11456
rect 5840 10368 6160 11392
rect 5840 10304 5848 10368
rect 5912 10304 5928 10368
rect 5992 10304 6008 10368
rect 6072 10304 6088 10368
rect 6152 10304 6160 10368
rect 5840 9280 6160 10304
rect 5840 9216 5848 9280
rect 5912 9216 5928 9280
rect 5992 9216 6008 9280
rect 6072 9216 6088 9280
rect 6152 9216 6160 9280
rect 5840 8192 6160 9216
rect 5840 8128 5848 8192
rect 5912 8128 5928 8192
rect 5992 8128 6008 8192
rect 6072 8128 6088 8192
rect 6152 8128 6160 8192
rect 5840 7104 6160 8128
rect 5840 7040 5848 7104
rect 5912 7040 5928 7104
rect 5992 7040 6008 7104
rect 6072 7040 6088 7104
rect 6152 7040 6160 7104
rect 5027 6764 5093 6765
rect 5027 6700 5028 6764
rect 5092 6700 5093 6764
rect 5027 6699 5093 6700
rect 5840 6016 6160 7040
rect 5840 5952 5848 6016
rect 5912 5952 5928 6016
rect 5992 5952 6008 6016
rect 6072 5952 6088 6016
rect 6152 5952 6160 6016
rect 4843 5268 4909 5269
rect 4843 5204 4844 5268
rect 4908 5204 4909 5268
rect 4843 5203 4909 5204
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 5840 4928 6160 5952
rect 5840 4864 5848 4928
rect 5912 4864 5928 4928
rect 5992 4864 6008 4928
rect 6072 4864 6088 4928
rect 6152 4864 6160 4928
rect 5840 3840 6160 4864
rect 5840 3776 5848 3840
rect 5912 3776 5928 3840
rect 5992 3776 6008 3840
rect 6072 3776 6088 3840
rect 6152 3776 6160 3840
rect 5840 2752 6160 3776
rect 5840 2688 5848 2752
rect 5912 2688 5928 2752
rect 5992 2688 6008 2752
rect 6072 2688 6088 2752
rect 6152 2688 6160 2752
rect 5840 2128 6160 2688
rect 7472 26144 7792 27168
rect 7472 26080 7480 26144
rect 7544 26080 7560 26144
rect 7624 26080 7640 26144
rect 7704 26080 7720 26144
rect 7784 26080 7792 26144
rect 7472 25056 7792 26080
rect 7472 24992 7480 25056
rect 7544 24992 7560 25056
rect 7624 24992 7640 25056
rect 7704 24992 7720 25056
rect 7784 24992 7792 25056
rect 7472 23968 7792 24992
rect 7472 23904 7480 23968
rect 7544 23904 7560 23968
rect 7624 23904 7640 23968
rect 7704 23904 7720 23968
rect 7784 23904 7792 23968
rect 7472 22880 7792 23904
rect 7472 22816 7480 22880
rect 7544 22816 7560 22880
rect 7624 22816 7640 22880
rect 7704 22816 7720 22880
rect 7784 22816 7792 22880
rect 7472 21792 7792 22816
rect 7472 21728 7480 21792
rect 7544 21728 7560 21792
rect 7624 21728 7640 21792
rect 7704 21728 7720 21792
rect 7784 21728 7792 21792
rect 7472 20704 7792 21728
rect 7472 20640 7480 20704
rect 7544 20640 7560 20704
rect 7624 20640 7640 20704
rect 7704 20640 7720 20704
rect 7784 20640 7792 20704
rect 7472 19616 7792 20640
rect 7472 19552 7480 19616
rect 7544 19552 7560 19616
rect 7624 19552 7640 19616
rect 7704 19552 7720 19616
rect 7784 19552 7792 19616
rect 7472 18528 7792 19552
rect 7472 18464 7480 18528
rect 7544 18464 7560 18528
rect 7624 18464 7640 18528
rect 7704 18464 7720 18528
rect 7784 18464 7792 18528
rect 7472 17440 7792 18464
rect 7472 17376 7480 17440
rect 7544 17376 7560 17440
rect 7624 17376 7640 17440
rect 7704 17376 7720 17440
rect 7784 17376 7792 17440
rect 7472 16352 7792 17376
rect 7472 16288 7480 16352
rect 7544 16288 7560 16352
rect 7624 16288 7640 16352
rect 7704 16288 7720 16352
rect 7784 16288 7792 16352
rect 7472 15264 7792 16288
rect 7472 15200 7480 15264
rect 7544 15200 7560 15264
rect 7624 15200 7640 15264
rect 7704 15200 7720 15264
rect 7784 15200 7792 15264
rect 7472 14176 7792 15200
rect 7472 14112 7480 14176
rect 7544 14112 7560 14176
rect 7624 14112 7640 14176
rect 7704 14112 7720 14176
rect 7784 14112 7792 14176
rect 7472 13088 7792 14112
rect 7472 13024 7480 13088
rect 7544 13024 7560 13088
rect 7624 13024 7640 13088
rect 7704 13024 7720 13088
rect 7784 13024 7792 13088
rect 7472 12000 7792 13024
rect 7472 11936 7480 12000
rect 7544 11936 7560 12000
rect 7624 11936 7640 12000
rect 7704 11936 7720 12000
rect 7784 11936 7792 12000
rect 7472 10912 7792 11936
rect 7472 10848 7480 10912
rect 7544 10848 7560 10912
rect 7624 10848 7640 10912
rect 7704 10848 7720 10912
rect 7784 10848 7792 10912
rect 7472 9824 7792 10848
rect 7472 9760 7480 9824
rect 7544 9760 7560 9824
rect 7624 9760 7640 9824
rect 7704 9760 7720 9824
rect 7784 9760 7792 9824
rect 7472 8736 7792 9760
rect 7472 8672 7480 8736
rect 7544 8672 7560 8736
rect 7624 8672 7640 8736
rect 7704 8672 7720 8736
rect 7784 8672 7792 8736
rect 7472 7648 7792 8672
rect 7472 7584 7480 7648
rect 7544 7584 7560 7648
rect 7624 7584 7640 7648
rect 7704 7584 7720 7648
rect 7784 7584 7792 7648
rect 7472 6560 7792 7584
rect 7472 6496 7480 6560
rect 7544 6496 7560 6560
rect 7624 6496 7640 6560
rect 7704 6496 7720 6560
rect 7784 6496 7792 6560
rect 7472 5472 7792 6496
rect 7472 5408 7480 5472
rect 7544 5408 7560 5472
rect 7624 5408 7640 5472
rect 7704 5408 7720 5472
rect 7784 5408 7792 5472
rect 7472 4384 7792 5408
rect 7472 4320 7480 4384
rect 7544 4320 7560 4384
rect 7624 4320 7640 4384
rect 7704 4320 7720 4384
rect 7784 4320 7792 4384
rect 7472 3296 7792 4320
rect 7472 3232 7480 3296
rect 7544 3232 7560 3296
rect 7624 3232 7640 3296
rect 7704 3232 7720 3296
rect 7784 3232 7792 3296
rect 7472 2208 7792 3232
rect 7472 2144 7480 2208
rect 7544 2144 7560 2208
rect 7624 2144 7640 2208
rect 7704 2144 7720 2208
rect 7784 2144 7792 2208
rect 7472 2128 7792 2144
rect 9104 77824 9424 77840
rect 9104 77760 9112 77824
rect 9176 77760 9192 77824
rect 9256 77760 9272 77824
rect 9336 77760 9352 77824
rect 9416 77760 9424 77824
rect 9104 76736 9424 77760
rect 9104 76672 9112 76736
rect 9176 76672 9192 76736
rect 9256 76672 9272 76736
rect 9336 76672 9352 76736
rect 9416 76672 9424 76736
rect 9104 75648 9424 76672
rect 9104 75584 9112 75648
rect 9176 75584 9192 75648
rect 9256 75584 9272 75648
rect 9336 75584 9352 75648
rect 9416 75584 9424 75648
rect 9104 74560 9424 75584
rect 9104 74496 9112 74560
rect 9176 74496 9192 74560
rect 9256 74496 9272 74560
rect 9336 74496 9352 74560
rect 9416 74496 9424 74560
rect 9104 73472 9424 74496
rect 9104 73408 9112 73472
rect 9176 73408 9192 73472
rect 9256 73408 9272 73472
rect 9336 73408 9352 73472
rect 9416 73408 9424 73472
rect 9104 72384 9424 73408
rect 9104 72320 9112 72384
rect 9176 72320 9192 72384
rect 9256 72320 9272 72384
rect 9336 72320 9352 72384
rect 9416 72320 9424 72384
rect 9104 71296 9424 72320
rect 9104 71232 9112 71296
rect 9176 71232 9192 71296
rect 9256 71232 9272 71296
rect 9336 71232 9352 71296
rect 9416 71232 9424 71296
rect 9104 70208 9424 71232
rect 9104 70144 9112 70208
rect 9176 70144 9192 70208
rect 9256 70144 9272 70208
rect 9336 70144 9352 70208
rect 9416 70144 9424 70208
rect 9104 69120 9424 70144
rect 9104 69056 9112 69120
rect 9176 69056 9192 69120
rect 9256 69056 9272 69120
rect 9336 69056 9352 69120
rect 9416 69056 9424 69120
rect 9104 68032 9424 69056
rect 9104 67968 9112 68032
rect 9176 67968 9192 68032
rect 9256 67968 9272 68032
rect 9336 67968 9352 68032
rect 9416 67968 9424 68032
rect 9104 66944 9424 67968
rect 9104 66880 9112 66944
rect 9176 66880 9192 66944
rect 9256 66880 9272 66944
rect 9336 66880 9352 66944
rect 9416 66880 9424 66944
rect 9104 65856 9424 66880
rect 9104 65792 9112 65856
rect 9176 65792 9192 65856
rect 9256 65792 9272 65856
rect 9336 65792 9352 65856
rect 9416 65792 9424 65856
rect 9104 64768 9424 65792
rect 9104 64704 9112 64768
rect 9176 64704 9192 64768
rect 9256 64704 9272 64768
rect 9336 64704 9352 64768
rect 9416 64704 9424 64768
rect 9104 63680 9424 64704
rect 9104 63616 9112 63680
rect 9176 63616 9192 63680
rect 9256 63616 9272 63680
rect 9336 63616 9352 63680
rect 9416 63616 9424 63680
rect 9104 62592 9424 63616
rect 9104 62528 9112 62592
rect 9176 62528 9192 62592
rect 9256 62528 9272 62592
rect 9336 62528 9352 62592
rect 9416 62528 9424 62592
rect 9104 61504 9424 62528
rect 9104 61440 9112 61504
rect 9176 61440 9192 61504
rect 9256 61440 9272 61504
rect 9336 61440 9352 61504
rect 9416 61440 9424 61504
rect 9104 60416 9424 61440
rect 9104 60352 9112 60416
rect 9176 60352 9192 60416
rect 9256 60352 9272 60416
rect 9336 60352 9352 60416
rect 9416 60352 9424 60416
rect 9104 59328 9424 60352
rect 9104 59264 9112 59328
rect 9176 59264 9192 59328
rect 9256 59264 9272 59328
rect 9336 59264 9352 59328
rect 9416 59264 9424 59328
rect 9104 58240 9424 59264
rect 9104 58176 9112 58240
rect 9176 58176 9192 58240
rect 9256 58176 9272 58240
rect 9336 58176 9352 58240
rect 9416 58176 9424 58240
rect 9104 57152 9424 58176
rect 9104 57088 9112 57152
rect 9176 57088 9192 57152
rect 9256 57088 9272 57152
rect 9336 57088 9352 57152
rect 9416 57088 9424 57152
rect 9104 56064 9424 57088
rect 9104 56000 9112 56064
rect 9176 56000 9192 56064
rect 9256 56000 9272 56064
rect 9336 56000 9352 56064
rect 9416 56000 9424 56064
rect 9104 54976 9424 56000
rect 9104 54912 9112 54976
rect 9176 54912 9192 54976
rect 9256 54912 9272 54976
rect 9336 54912 9352 54976
rect 9416 54912 9424 54976
rect 9104 53888 9424 54912
rect 9104 53824 9112 53888
rect 9176 53824 9192 53888
rect 9256 53824 9272 53888
rect 9336 53824 9352 53888
rect 9416 53824 9424 53888
rect 9104 52800 9424 53824
rect 9104 52736 9112 52800
rect 9176 52736 9192 52800
rect 9256 52736 9272 52800
rect 9336 52736 9352 52800
rect 9416 52736 9424 52800
rect 9104 51712 9424 52736
rect 9104 51648 9112 51712
rect 9176 51648 9192 51712
rect 9256 51648 9272 51712
rect 9336 51648 9352 51712
rect 9416 51648 9424 51712
rect 9104 50624 9424 51648
rect 9104 50560 9112 50624
rect 9176 50560 9192 50624
rect 9256 50560 9272 50624
rect 9336 50560 9352 50624
rect 9416 50560 9424 50624
rect 9104 49536 9424 50560
rect 9104 49472 9112 49536
rect 9176 49472 9192 49536
rect 9256 49472 9272 49536
rect 9336 49472 9352 49536
rect 9416 49472 9424 49536
rect 9104 48448 9424 49472
rect 9104 48384 9112 48448
rect 9176 48384 9192 48448
rect 9256 48384 9272 48448
rect 9336 48384 9352 48448
rect 9416 48384 9424 48448
rect 9104 47360 9424 48384
rect 9104 47296 9112 47360
rect 9176 47296 9192 47360
rect 9256 47296 9272 47360
rect 9336 47296 9352 47360
rect 9416 47296 9424 47360
rect 9104 46272 9424 47296
rect 9104 46208 9112 46272
rect 9176 46208 9192 46272
rect 9256 46208 9272 46272
rect 9336 46208 9352 46272
rect 9416 46208 9424 46272
rect 9104 45184 9424 46208
rect 9104 45120 9112 45184
rect 9176 45120 9192 45184
rect 9256 45120 9272 45184
rect 9336 45120 9352 45184
rect 9416 45120 9424 45184
rect 9104 44096 9424 45120
rect 9104 44032 9112 44096
rect 9176 44032 9192 44096
rect 9256 44032 9272 44096
rect 9336 44032 9352 44096
rect 9416 44032 9424 44096
rect 9104 43008 9424 44032
rect 9104 42944 9112 43008
rect 9176 42944 9192 43008
rect 9256 42944 9272 43008
rect 9336 42944 9352 43008
rect 9416 42944 9424 43008
rect 9104 41920 9424 42944
rect 9104 41856 9112 41920
rect 9176 41856 9192 41920
rect 9256 41856 9272 41920
rect 9336 41856 9352 41920
rect 9416 41856 9424 41920
rect 9104 40832 9424 41856
rect 9104 40768 9112 40832
rect 9176 40768 9192 40832
rect 9256 40768 9272 40832
rect 9336 40768 9352 40832
rect 9416 40768 9424 40832
rect 9104 39744 9424 40768
rect 9104 39680 9112 39744
rect 9176 39680 9192 39744
rect 9256 39680 9272 39744
rect 9336 39680 9352 39744
rect 9416 39680 9424 39744
rect 9104 38656 9424 39680
rect 9104 38592 9112 38656
rect 9176 38592 9192 38656
rect 9256 38592 9272 38656
rect 9336 38592 9352 38656
rect 9416 38592 9424 38656
rect 9104 37568 9424 38592
rect 9104 37504 9112 37568
rect 9176 37504 9192 37568
rect 9256 37504 9272 37568
rect 9336 37504 9352 37568
rect 9416 37504 9424 37568
rect 9104 36480 9424 37504
rect 9104 36416 9112 36480
rect 9176 36416 9192 36480
rect 9256 36416 9272 36480
rect 9336 36416 9352 36480
rect 9416 36416 9424 36480
rect 9104 35392 9424 36416
rect 9104 35328 9112 35392
rect 9176 35328 9192 35392
rect 9256 35328 9272 35392
rect 9336 35328 9352 35392
rect 9416 35328 9424 35392
rect 9104 34304 9424 35328
rect 9104 34240 9112 34304
rect 9176 34240 9192 34304
rect 9256 34240 9272 34304
rect 9336 34240 9352 34304
rect 9416 34240 9424 34304
rect 9104 33216 9424 34240
rect 9104 33152 9112 33216
rect 9176 33152 9192 33216
rect 9256 33152 9272 33216
rect 9336 33152 9352 33216
rect 9416 33152 9424 33216
rect 9104 32128 9424 33152
rect 9104 32064 9112 32128
rect 9176 32064 9192 32128
rect 9256 32064 9272 32128
rect 9336 32064 9352 32128
rect 9416 32064 9424 32128
rect 9104 31040 9424 32064
rect 9104 30976 9112 31040
rect 9176 30976 9192 31040
rect 9256 30976 9272 31040
rect 9336 30976 9352 31040
rect 9416 30976 9424 31040
rect 9104 29952 9424 30976
rect 9104 29888 9112 29952
rect 9176 29888 9192 29952
rect 9256 29888 9272 29952
rect 9336 29888 9352 29952
rect 9416 29888 9424 29952
rect 9104 28864 9424 29888
rect 9104 28800 9112 28864
rect 9176 28800 9192 28864
rect 9256 28800 9272 28864
rect 9336 28800 9352 28864
rect 9416 28800 9424 28864
rect 9104 27776 9424 28800
rect 9104 27712 9112 27776
rect 9176 27712 9192 27776
rect 9256 27712 9272 27776
rect 9336 27712 9352 27776
rect 9416 27712 9424 27776
rect 9104 26688 9424 27712
rect 9104 26624 9112 26688
rect 9176 26624 9192 26688
rect 9256 26624 9272 26688
rect 9336 26624 9352 26688
rect 9416 26624 9424 26688
rect 9104 25600 9424 26624
rect 9104 25536 9112 25600
rect 9176 25536 9192 25600
rect 9256 25536 9272 25600
rect 9336 25536 9352 25600
rect 9416 25536 9424 25600
rect 9104 24512 9424 25536
rect 9104 24448 9112 24512
rect 9176 24448 9192 24512
rect 9256 24448 9272 24512
rect 9336 24448 9352 24512
rect 9416 24448 9424 24512
rect 9104 23424 9424 24448
rect 9104 23360 9112 23424
rect 9176 23360 9192 23424
rect 9256 23360 9272 23424
rect 9336 23360 9352 23424
rect 9416 23360 9424 23424
rect 9104 22336 9424 23360
rect 9104 22272 9112 22336
rect 9176 22272 9192 22336
rect 9256 22272 9272 22336
rect 9336 22272 9352 22336
rect 9416 22272 9424 22336
rect 9104 21248 9424 22272
rect 9104 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9272 21248
rect 9336 21184 9352 21248
rect 9416 21184 9424 21248
rect 9104 20160 9424 21184
rect 9104 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9272 20160
rect 9336 20096 9352 20160
rect 9416 20096 9424 20160
rect 9104 19072 9424 20096
rect 9104 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9272 19072
rect 9336 19008 9352 19072
rect 9416 19008 9424 19072
rect 9104 17984 9424 19008
rect 9104 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9272 17984
rect 9336 17920 9352 17984
rect 9416 17920 9424 17984
rect 9104 16896 9424 17920
rect 9104 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9272 16896
rect 9336 16832 9352 16896
rect 9416 16832 9424 16896
rect 9104 15808 9424 16832
rect 9104 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9272 15808
rect 9336 15744 9352 15808
rect 9416 15744 9424 15808
rect 9104 14720 9424 15744
rect 9104 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9272 14720
rect 9336 14656 9352 14720
rect 9416 14656 9424 14720
rect 9104 13632 9424 14656
rect 9104 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9272 13632
rect 9336 13568 9352 13632
rect 9416 13568 9424 13632
rect 9104 12544 9424 13568
rect 9104 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9272 12544
rect 9336 12480 9352 12544
rect 9416 12480 9424 12544
rect 9104 11456 9424 12480
rect 9104 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9272 11456
rect 9336 11392 9352 11456
rect 9416 11392 9424 11456
rect 9104 10368 9424 11392
rect 9104 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9272 10368
rect 9336 10304 9352 10368
rect 9416 10304 9424 10368
rect 9104 9280 9424 10304
rect 9104 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9272 9280
rect 9336 9216 9352 9280
rect 9416 9216 9424 9280
rect 9104 8192 9424 9216
rect 9104 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9272 8192
rect 9336 8128 9352 8192
rect 9416 8128 9424 8192
rect 9104 7104 9424 8128
rect 9104 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9272 7104
rect 9336 7040 9352 7104
rect 9416 7040 9424 7104
rect 9104 6016 9424 7040
rect 9104 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9272 6016
rect 9336 5952 9352 6016
rect 9416 5952 9424 6016
rect 9104 4928 9424 5952
rect 9104 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9272 4928
rect 9336 4864 9352 4928
rect 9416 4864 9424 4928
rect 9104 3840 9424 4864
rect 9104 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9272 3840
rect 9336 3776 9352 3840
rect 9416 3776 9424 3840
rect 9104 2752 9424 3776
rect 9104 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9272 2752
rect 9336 2688 9352 2752
rect 9416 2688 9424 2752
rect 9104 2128 9424 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4324 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1644511149
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91
timestamp 1644511149
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6
timestamp 1644511149
transform 1 0 1656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 1644511149
transform 1 0 2944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1644511149
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_91
timestamp 1644511149
transform 1 0 9476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_99
timestamp 1644511149
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6
timestamp 1644511149
transform 1 0 1656 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_12
timestamp 1644511149
transform 1 0 2208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_16
timestamp 1644511149
transform 1 0 2576 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1644511149
transform 1 0 4692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_51
timestamp 1644511149
transform 1 0 5796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_63
timestamp 1644511149
transform 1 0 6900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1644511149
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1644511149
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1644511149
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_21
timestamp 1644511149
transform 1 0 3036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1644511149
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_46
timestamp 1644511149
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1644511149
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1644511149
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1644511149
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_34
timestamp 1644511149
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1644511149
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_99
timestamp 1644511149
transform 1 0 10212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1644511149
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_21
timestamp 1644511149
transform 1 0 3036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_28
timestamp 1644511149
transform 1 0 3680 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_34
timestamp 1644511149
transform 1 0 4232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_38
timestamp 1644511149
transform 1 0 4600 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1644511149
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 1644511149
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_91
timestamp 1644511149
transform 1 0 9476 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1644511149
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1644511149
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1644511149
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1644511149
transform 1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1644511149
transform 1 0 4692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_51
timestamp 1644511149
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_63
timestamp 1644511149
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1644511149
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1644511149
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1644511149
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_10
timestamp 1644511149
transform 1 0 2024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_18
timestamp 1644511149
transform 1 0 2760 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_29
timestamp 1644511149
transform 1 0 3772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_41
timestamp 1644511149
transform 1 0 4876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1644511149
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1644511149
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1644511149
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1644511149
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_37
timestamp 1644511149
transform 1 0 4508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_49
timestamp 1644511149
transform 1 0 5612 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_61
timestamp 1644511149
transform 1 0 6716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_73
timestamp 1644511149
transform 1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1644511149
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1644511149
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_99
timestamp 1644511149
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_14
timestamp 1644511149
transform 1 0 2392 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_22
timestamp 1644511149
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1644511149
transform 1 0 3864 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_37
timestamp 1644511149
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1644511149
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1644511149
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1644511149
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1644511149
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1644511149
transform 1 0 4048 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1644511149
transform 1 0 5152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1644511149
transform 1 0 6256 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1644511149
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1644511149
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_13
timestamp 1644511149
transform 1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_21
timestamp 1644511149
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_33
timestamp 1644511149
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_45
timestamp 1644511149
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1644511149
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1644511149
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1644511149
transform 1 0 4048 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1644511149
transform 1 0 5152 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1644511149
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1644511149
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1644511149
transform 1 0 9660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_99
timestamp 1644511149
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1644511149
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1644511149
transform 1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_28
timestamp 1644511149
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_35
timestamp 1644511149
transform 1 0 4324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1644511149
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_99
timestamp 1644511149
transform 1 0 10212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1644511149
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1644511149
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_33
timestamp 1644511149
transform 1 0 4140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_45
timestamp 1644511149
transform 1 0 5244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_57
timestamp 1644511149
transform 1 0 6348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_69
timestamp 1644511149
transform 1 0 7452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_81
timestamp 1644511149
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1644511149
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1644511149
transform 1 0 3036 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_28
timestamp 1644511149
transform 1 0 3680 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_40
timestamp 1644511149
transform 1 0 4784 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1644511149
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1644511149
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp 1644511149
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1644511149
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1644511149
transform 1 0 9660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_99
timestamp 1644511149
transform 1 0 10212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1644511149
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_22
timestamp 1644511149
transform 1 0 3128 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_29
timestamp 1644511149
transform 1 0 3772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_41
timestamp 1644511149
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1644511149
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_99
timestamp 1644511149
transform 1 0 10212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_13
timestamp 1644511149
transform 1 0 2300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1644511149
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1644511149
transform 1 0 9660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_99
timestamp 1644511149
transform 1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_9
timestamp 1644511149
transform 1 0 1932 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_22
timestamp 1644511149
transform 1 0 3128 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_29
timestamp 1644511149
transform 1 0 3772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_41
timestamp 1644511149
transform 1 0 4876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1644511149
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1644511149
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_6
timestamp 1644511149
transform 1 0 1656 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_14
timestamp 1644511149
transform 1 0 2392 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1644511149
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1644511149
transform 1 0 4048 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1644511149
transform 1 0 5152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1644511149
transform 1 0 6256 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1644511149
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_92
timestamp 1644511149
transform 1 0 9568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99
timestamp 1644511149
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_6
timestamp 1644511149
transform 1 0 1656 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_14
timestamp 1644511149
transform 1 0 2392 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_19
timestamp 1644511149
transform 1 0 2852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_26
timestamp 1644511149
transform 1 0 3496 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_38
timestamp 1644511149
transform 1 0 4600 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1644511149
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_87
timestamp 1644511149
transform 1 0 9108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_91
timestamp 1644511149
transform 1 0 9476 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1644511149
transform 1 0 10212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_9
timestamp 1644511149
transform 1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_18
timestamp 1644511149
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1644511149
transform 1 0 4048 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1644511149
transform 1 0 5152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1644511149
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1644511149
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1644511149
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1644511149
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1644511149
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_12
timestamp 1644511149
transform 1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_19
timestamp 1644511149
transform 1 0 2852 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_31
timestamp 1644511149
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_43
timestamp 1644511149
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_99
timestamp 1644511149
transform 1 0 10212 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_12
timestamp 1644511149
transform 1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1644511149
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1644511149
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_99
timestamp 1644511149
transform 1 0 10212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_13
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_20
timestamp 1644511149
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_32
timestamp 1644511149
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_44
timestamp 1644511149
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 1644511149
transform 1 0 9108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_91
timestamp 1644511149
transform 1 0 9476 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1644511149
transform 1 0 10212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_6
timestamp 1644511149
transform 1 0 1656 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1644511149
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1644511149
transform 1 0 4048 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1644511149
transform 1 0 5152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1644511149
transform 1 0 6256 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1644511149
transform 1 0 7360 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1644511149
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1644511149
transform 1 0 10212 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_28
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_40
timestamp 1644511149
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_99
timestamp 1644511149
transform 1 0 10212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_6
timestamp 1644511149
transform 1 0 1656 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_10
timestamp 1644511149
transform 1 0 2024 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_34
timestamp 1644511149
transform 1 0 4232 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_46
timestamp 1644511149
transform 1 0 5336 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_58
timestamp 1644511149
transform 1 0 6440 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_70
timestamp 1644511149
transform 1 0 7544 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1644511149
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1644511149
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_99
timestamp 1644511149
transform 1 0 10212 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_11
timestamp 1644511149
transform 1 0 2116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_22
timestamp 1644511149
transform 1 0 3128 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_29
timestamp 1644511149
transform 1 0 3772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_41
timestamp 1644511149
transform 1 0 4876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1644511149
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_99
timestamp 1644511149
transform 1 0 10212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_13
timestamp 1644511149
transform 1 0 2300 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1644511149
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1644511149
transform 1 0 4048 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1644511149
transform 1 0 5152 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1644511149
transform 1 0 6256 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1644511149
transform 1 0 7360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1644511149
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1644511149
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_99
timestamp 1644511149
transform 1 0 10212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_13
timestamp 1644511149
transform 1 0 2300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_21
timestamp 1644511149
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_33
timestamp 1644511149
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1644511149
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1644511149
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_87
timestamp 1644511149
transform 1 0 9108 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_91
timestamp 1644511149
transform 1 0 9476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_98
timestamp 1644511149
transform 1 0 10120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_102
timestamp 1644511149
transform 1 0 10488 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_13
timestamp 1644511149
transform 1 0 2300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_22
timestamp 1644511149
transform 1 0 3128 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1644511149
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1644511149
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_13
timestamp 1644511149
transform 1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_99
timestamp 1644511149
transform 1 0 10212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_13
timestamp 1644511149
transform 1 0 2300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1644511149
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_13
timestamp 1644511149
transform 1 0 2300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1644511149
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_29
timestamp 1644511149
transform 1 0 3772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_41
timestamp 1644511149
transform 1 0 4876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1644511149
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_99
timestamp 1644511149
transform 1 0 10212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1644511149
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1644511149
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_93
timestamp 1644511149
transform 1 0 9660 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1644511149
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_11
timestamp 1644511149
transform 1 0 2116 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1644511149
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_29
timestamp 1644511149
transform 1 0 3772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_41
timestamp 1644511149
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1644511149
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_99
timestamp 1644511149
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_13
timestamp 1644511149
transform 1 0 2300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1644511149
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_37
timestamp 1644511149
transform 1 0 4508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_45
timestamp 1644511149
transform 1 0 5244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_57
timestamp 1644511149
transform 1 0 6348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_69
timestamp 1644511149
transform 1 0 7452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_81
timestamp 1644511149
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_13
timestamp 1644511149
transform 1 0 2300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_22
timestamp 1644511149
transform 1 0 3128 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_28
timestamp 1644511149
transform 1 0 3680 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_46
timestamp 1644511149
transform 1 0 5336 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1644511149
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_99
timestamp 1644511149
transform 1 0 10212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1644511149
transform 1 0 2116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1644511149
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_39
timestamp 1644511149
transform 1 0 4692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_51
timestamp 1644511149
transform 1 0 5796 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_63
timestamp 1644511149
transform 1 0 6900 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_75
timestamp 1644511149
transform 1 0 8004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_93
timestamp 1644511149
transform 1 0 9660 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1644511149
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_10
timestamp 1644511149
transform 1 0 2024 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_19
timestamp 1644511149
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_31
timestamp 1644511149
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_43
timestamp 1644511149
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_101
timestamp 1644511149
transform 1 0 10396 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1644511149
transform 1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_19
timestamp 1644511149
transform 1 0 2852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_33
timestamp 1644511149
transform 1 0 4140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_45
timestamp 1644511149
transform 1 0 5244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_57
timestamp 1644511149
transform 1 0 6348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_69
timestamp 1644511149
transform 1 0 7452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1644511149
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_93
timestamp 1644511149
transform 1 0 9660 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1644511149
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_11
timestamp 1644511149
transform 1 0 2116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_19
timestamp 1644511149
transform 1 0 2852 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_99
timestamp 1644511149
transform 1 0 10212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_11
timestamp 1644511149
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1644511149
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_7
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_16
timestamp 1644511149
transform 1 0 2576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_24
timestamp 1644511149
transform 1 0 3312 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_36
timestamp 1644511149
transform 1 0 4416 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_48
timestamp 1644511149
transform 1 0 5520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_99
timestamp 1644511149
transform 1 0 10212 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_13
timestamp 1644511149
transform 1 0 2300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1644511149
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_93
timestamp 1644511149
transform 1 0 9660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_99
timestamp 1644511149
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_12
timestamp 1644511149
transform 1 0 2208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_20
timestamp 1644511149
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_32
timestamp 1644511149
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_44
timestamp 1644511149
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_99
timestamp 1644511149
transform 1 0 10212 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_10
timestamp 1644511149
transform 1 0 2024 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1644511149
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1644511149
transform 1 0 4048 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_44
timestamp 1644511149
transform 1 0 5152 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_56
timestamp 1644511149
transform 1 0 6256 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_68
timestamp 1644511149
transform 1 0 7360 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1644511149
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_11
timestamp 1644511149
transform 1 0 2116 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_19
timestamp 1644511149
transform 1 0 2852 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_99
timestamp 1644511149
transform 1 0 10212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_11
timestamp 1644511149
transform 1 0 2116 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_22
timestamp 1644511149
transform 1 0 3128 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_93
timestamp 1644511149
transform 1 0 9660 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_99
timestamp 1644511149
transform 1 0 10212 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_11
timestamp 1644511149
transform 1 0 2116 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_19
timestamp 1644511149
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_31
timestamp 1644511149
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_43
timestamp 1644511149
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_101
timestamp 1644511149
transform 1 0 10396 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_7
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_16
timestamp 1644511149
transform 1 0 2576 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_93
timestamp 1644511149
transform 1 0 9660 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_99
timestamp 1644511149
transform 1 0 10212 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_13
timestamp 1644511149
transform 1 0 2300 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_21
timestamp 1644511149
transform 1 0 3036 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_29
timestamp 1644511149
transform 1 0 3772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_41
timestamp 1644511149
transform 1 0 4876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1644511149
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_99
timestamp 1644511149
transform 1 0 10212 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_8
timestamp 1644511149
transform 1 0 1840 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1644511149
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_33
timestamp 1644511149
transform 1 0 4140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_45
timestamp 1644511149
transform 1 0 5244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_57
timestamp 1644511149
transform 1 0 6348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_69
timestamp 1644511149
transform 1 0 7452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_81
timestamp 1644511149
transform 1 0 8556 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_93
timestamp 1644511149
transform 1 0 9660 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_99
timestamp 1644511149
transform 1 0 10212 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_8
timestamp 1644511149
transform 1 0 1840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_17
timestamp 1644511149
transform 1 0 2668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_25
timestamp 1644511149
transform 1 0 3404 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_33
timestamp 1644511149
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1644511149
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1644511149
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_101
timestamp 1644511149
transform 1 0 10396 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_9
timestamp 1644511149
transform 1 0 1932 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_14
timestamp 1644511149
transform 1 0 2392 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_23
timestamp 1644511149
transform 1 0 3220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_33
timestamp 1644511149
transform 1 0 4140 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_93
timestamp 1644511149
transform 1 0 9660 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_99
timestamp 1644511149
transform 1 0 10212 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_12
timestamp 1644511149
transform 1 0 2208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_21
timestamp 1644511149
transform 1 0 3036 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_30
timestamp 1644511149
transform 1 0 3864 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_37
timestamp 1644511149
transform 1 0 4508 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_45
timestamp 1644511149
transform 1 0 5244 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_99
timestamp 1644511149
transform 1 0 10212 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_11
timestamp 1644511149
transform 1 0 2116 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_19
timestamp 1644511149
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_47
timestamp 1644511149
transform 1 0 5428 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_59
timestamp 1644511149
transform 1 0 6532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_71
timestamp 1644511149
transform 1 0 7636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_7
timestamp 1644511149
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_23
timestamp 1644511149
transform 1 0 3220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_32
timestamp 1644511149
transform 1 0 4048 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_44
timestamp 1644511149
transform 1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_99
timestamp 1644511149
transform 1 0 10212 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_7
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1644511149
transform 1 0 4048 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_44
timestamp 1644511149
transform 1 0 5152 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_56
timestamp 1644511149
transform 1 0 6256 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_68
timestamp 1644511149
transform 1 0 7360 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1644511149
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_93
timestamp 1644511149
transform 1 0 9660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_99
timestamp 1644511149
transform 1 0 10212 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_7
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_21
timestamp 1644511149
transform 1 0 3036 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_29
timestamp 1644511149
transform 1 0 3772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_36
timestamp 1644511149
transform 1 0 4416 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_48
timestamp 1644511149
transform 1 0 5520 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_62
timestamp 1644511149
transform 1 0 6808 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_74
timestamp 1644511149
transform 1 0 7912 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_86
timestamp 1644511149
transform 1 0 9016 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_98
timestamp 1644511149
transform 1 0 10120 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_102
timestamp 1644511149
transform 1 0 10488 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_11
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_33
timestamp 1644511149
transform 1 0 4140 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_40
timestamp 1644511149
transform 1 0 4784 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_52
timestamp 1644511149
transform 1 0 5888 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_64
timestamp 1644511149
transform 1 0 6992 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_76
timestamp 1644511149
transform 1 0 8096 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_93
timestamp 1644511149
transform 1 0 9660 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_99
timestamp 1644511149
transform 1 0 10212 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_9
timestamp 1644511149
transform 1 0 1932 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_23
timestamp 1644511149
transform 1 0 3220 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_35
timestamp 1644511149
transform 1 0 4324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1644511149
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_60
timestamp 1644511149
transform 1 0 6624 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_67
timestamp 1644511149
transform 1 0 7268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_79
timestamp 1644511149
transform 1 0 8372 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_91
timestamp 1644511149
transform 1 0 9476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_99
timestamp 1644511149
transform 1 0 10212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_9
timestamp 1644511149
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_18
timestamp 1644511149
transform 1 0 2760 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1644511149
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_33
timestamp 1644511149
transform 1 0 4140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_45
timestamp 1644511149
transform 1 0 5244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_69
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 1644511149
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_93
timestamp 1644511149
transform 1 0 9660 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_99
timestamp 1644511149
transform 1 0 10212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_9
timestamp 1644511149
transform 1 0 1932 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_18
timestamp 1644511149
transform 1 0 2760 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_26
timestamp 1644511149
transform 1 0 3496 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_38
timestamp 1644511149
transform 1 0 4600 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_44
timestamp 1644511149
transform 1 0 5152 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_101
timestamp 1644511149
transform 1 0 10396 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_14
timestamp 1644511149
transform 1 0 2392 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1644511149
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_46
timestamp 1644511149
transform 1 0 5336 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_58
timestamp 1644511149
transform 1 0 6440 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_70
timestamp 1644511149
transform 1 0 7544 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1644511149
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_93
timestamp 1644511149
transform 1 0 9660 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_99
timestamp 1644511149
transform 1 0 10212 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_14
timestamp 1644511149
transform 1 0 2392 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_22
timestamp 1644511149
transform 1 0 3128 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_30
timestamp 1644511149
transform 1 0 3864 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_42
timestamp 1644511149
transform 1 0 4968 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1644511149
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_62
timestamp 1644511149
transform 1 0 6808 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_74
timestamp 1644511149
transform 1 0 7912 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_86
timestamp 1644511149
transform 1 0 9016 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_94
timestamp 1644511149
transform 1 0 9752 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_99
timestamp 1644511149
transform 1 0 10212 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_7
timestamp 1644511149
transform 1 0 1748 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_23
timestamp 1644511149
transform 1 0 3220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_33
timestamp 1644511149
transform 1 0 4140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_50
timestamp 1644511149
transform 1 0 5704 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_58
timestamp 1644511149
transform 1 0 6440 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_63
timestamp 1644511149
transform 1 0 6900 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_75
timestamp 1644511149
transform 1 0 8004 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_93
timestamp 1644511149
transform 1 0 9660 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_98
timestamp 1644511149
transform 1 0 10120 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_102
timestamp 1644511149
transform 1 0 10488 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_9
timestamp 1644511149
transform 1 0 1932 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_25
timestamp 1644511149
transform 1 0 3404 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_33
timestamp 1644511149
transform 1 0 4140 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_45
timestamp 1644511149
transform 1 0 5244 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_53
timestamp 1644511149
transform 1 0 5980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_87
timestamp 1644511149
transform 1 0 9108 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_91
timestamp 1644511149
transform 1 0 9476 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_99
timestamp 1644511149
transform 1 0 10212 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_7
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_21
timestamp 1644511149
transform 1 0 3036 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_33
timestamp 1644511149
transform 1 0 4140 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_45
timestamp 1644511149
transform 1 0 5244 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_57
timestamp 1644511149
transform 1 0 6348 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_69
timestamp 1644511149
transform 1 0 7452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_81
timestamp 1644511149
transform 1 0 8556 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_91
timestamp 1644511149
transform 1 0 9476 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_99
timestamp 1644511149
transform 1 0 10212 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_10
timestamp 1644511149
transform 1 0 2024 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_14
timestamp 1644511149
transform 1 0 2392 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_20
timestamp 1644511149
transform 1 0 2944 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_28
timestamp 1644511149
transform 1 0 3680 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_40
timestamp 1644511149
transform 1 0 4784 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_47
timestamp 1644511149
transform 1 0 5428 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_99
timestamp 1644511149
transform 1 0 10212 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_10
timestamp 1644511149
transform 1 0 2024 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_37
timestamp 1644511149
transform 1 0 4508 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_44
timestamp 1644511149
transform 1 0 5152 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_56
timestamp 1644511149
transform 1 0 6256 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_68
timestamp 1644511149
transform 1 0 7360 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_80
timestamp 1644511149
transform 1 0 8464 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_93
timestamp 1644511149
transform 1 0 9660 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_99
timestamp 1644511149
transform 1 0 10212 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_15
timestamp 1644511149
transform 1 0 2484 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_99
timestamp 1644511149
transform 1 0 10212 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_12
timestamp 1644511149
transform 1 0 2208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_20
timestamp 1644511149
transform 1 0 2944 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_33
timestamp 1644511149
transform 1 0 4140 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_45
timestamp 1644511149
transform 1 0 5244 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_59
timestamp 1644511149
transform 1 0 6532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_71
timestamp 1644511149
transform 1 0 7636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_93
timestamp 1644511149
transform 1 0 9660 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_99
timestamp 1644511149
transform 1 0 10212 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_14
timestamp 1644511149
transform 1 0 2392 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_25
timestamp 1644511149
transform 1 0 3404 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1644511149
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1644511149
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_99
timestamp 1644511149
transform 1 0 10212 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_9
timestamp 1644511149
transform 1 0 1932 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_18
timestamp 1644511149
transform 1 0 2760 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_26
timestamp 1644511149
transform 1 0 3496 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_33
timestamp 1644511149
transform 1 0 4140 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_42
timestamp 1644511149
transform 1 0 4968 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_54
timestamp 1644511149
transform 1 0 6072 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_66
timestamp 1644511149
transform 1 0 7176 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_78
timestamp 1644511149
transform 1 0 8280 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_93
timestamp 1644511149
transform 1 0 9660 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_99
timestamp 1644511149
transform 1 0 10212 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_16
timestamp 1644511149
transform 1 0 2576 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_24
timestamp 1644511149
transform 1 0 3312 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_36
timestamp 1644511149
transform 1 0 4416 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_48
timestamp 1644511149
transform 1 0 5520 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_60
timestamp 1644511149
transform 1 0 6624 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_72
timestamp 1644511149
transform 1 0 7728 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_84
timestamp 1644511149
transform 1 0 8832 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_92
timestamp 1644511149
transform 1 0 9568 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_99
timestamp 1644511149
transform 1 0 10212 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_14
timestamp 1644511149
transform 1 0 2392 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_22
timestamp 1644511149
transform 1 0 3128 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_47
timestamp 1644511149
transform 1 0 5428 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_56
timestamp 1644511149
transform 1 0 6256 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_63
timestamp 1644511149
transform 1 0 6900 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_75
timestamp 1644511149
transform 1 0 8004 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_93
timestamp 1644511149
transform 1 0 9660 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_99
timestamp 1644511149
transform 1 0 10212 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_7
timestamp 1644511149
transform 1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_15
timestamp 1644511149
transform 1 0 2484 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_23
timestamp 1644511149
transform 1 0 3220 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_35
timestamp 1644511149
transform 1 0 4324 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_47
timestamp 1644511149
transform 1 0 5428 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_60
timestamp 1644511149
transform 1 0 6624 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_72
timestamp 1644511149
transform 1 0 7728 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_84
timestamp 1644511149
transform 1 0 8832 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_96
timestamp 1644511149
transform 1 0 9936 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_102
timestamp 1644511149
transform 1 0 10488 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_9
timestamp 1644511149
transform 1 0 1932 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_23
timestamp 1644511149
transform 1 0 3220 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_93
timestamp 1644511149
transform 1 0 9660 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_99
timestamp 1644511149
transform 1 0 10212 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_19
timestamp 1644511149
transform 1 0 2852 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1644511149
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1644511149
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1644511149
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_62
timestamp 1644511149
transform 1 0 6808 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_70
timestamp 1644511149
transform 1 0 7544 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_76
timestamp 1644511149
transform 1 0 8096 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_88
timestamp 1644511149
transform 1 0 9200 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_94
timestamp 1644511149
transform 1 0 9752 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_99
timestamp 1644511149
transform 1 0 10212 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_10
timestamp 1644511149
transform 1 0 2024 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_19
timestamp 1644511149
transform 1 0 2852 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_33
timestamp 1644511149
transform 1 0 4140 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_42
timestamp 1644511149
transform 1 0 4968 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_65
timestamp 1644511149
transform 1 0 7084 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_71
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_75
timestamp 1644511149
transform 1 0 8004 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_99
timestamp 1644511149
transform 1 0 10212 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_7
timestamp 1644511149
transform 1 0 1748 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_15
timestamp 1644511149
transform 1 0 2484 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_26
timestamp 1644511149
transform 1 0 3496 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_38
timestamp 1644511149
transform 1 0 4600 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_50
timestamp 1644511149
transform 1 0 5704 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1644511149
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1644511149
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_93
timestamp 1644511149
transform 1 0 9660 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_99
timestamp 1644511149
transform 1 0 10212 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_7
timestamp 1644511149
transform 1 0 1748 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_13
timestamp 1644511149
transform 1 0 2300 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_24
timestamp 1644511149
transform 1 0 3312 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1644511149
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1644511149
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1644511149
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1644511149
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1644511149
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_91
timestamp 1644511149
transform 1 0 9476 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_99
timestamp 1644511149
transform 1 0 10212 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_10
timestamp 1644511149
transform 1 0 2024 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_85_23
timestamp 1644511149
transform 1 0 3220 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_31
timestamp 1644511149
transform 1 0 3956 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_43
timestamp 1644511149
transform 1 0 5060 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1644511149
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1644511149
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_81
timestamp 1644511149
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_93
timestamp 1644511149
transform 1 0 9660 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_99
timestamp 1644511149
transform 1 0 10212 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_10
timestamp 1644511149
transform 1 0 2024 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_19
timestamp 1644511149
transform 1 0 2852 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1644511149
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_33
timestamp 1644511149
transform 1 0 4140 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_45
timestamp 1644511149
transform 1 0 5244 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_57
timestamp 1644511149
transform 1 0 6348 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_69
timestamp 1644511149
transform 1 0 7452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_81
timestamp 1644511149
transform 1 0 8556 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_86_85
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_93
timestamp 1644511149
transform 1 0 9660 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_99
timestamp 1644511149
transform 1 0 10212 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_10
timestamp 1644511149
transform 1 0 2024 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_18
timestamp 1644511149
transform 1 0 2760 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_25
timestamp 1644511149
transform 1 0 3404 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_37
timestamp 1644511149
transform 1 0 4508 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_49
timestamp 1644511149
transform 1 0 5612 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1644511149
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1644511149
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1644511149
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1644511149
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_93
timestamp 1644511149
transform 1 0 9660 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_99
timestamp 1644511149
transform 1 0 10212 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_10
timestamp 1644511149
transform 1 0 2024 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_18
timestamp 1644511149
transform 1 0 2760 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1644511149
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_88_29
timestamp 1644511149
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_41
timestamp 1644511149
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_53
timestamp 1644511149
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_65
timestamp 1644511149
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1644511149
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1644511149
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_85
timestamp 1644511149
transform 1 0 8924 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_93
timestamp 1644511149
transform 1 0 9660 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_99
timestamp 1644511149
transform 1 0 10212 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_7
timestamp 1644511149
transform 1 0 1748 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1644511149
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1644511149
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_39
timestamp 1644511149
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1644511149
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1644511149
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1644511149
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1644511149
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1644511149
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_93
timestamp 1644511149
transform 1 0 9660 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_99
timestamp 1644511149
transform 1 0 10212 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_7
timestamp 1644511149
transform 1 0 1748 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_13
timestamp 1644511149
transform 1 0 2300 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_19
timestamp 1644511149
transform 1 0 2852 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1644511149
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1644511149
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_41
timestamp 1644511149
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_53
timestamp 1644511149
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_65
timestamp 1644511149
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1644511149
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1644511149
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_85
timestamp 1644511149
transform 1 0 8924 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_93
timestamp 1644511149
transform 1 0 9660 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_99
timestamp 1644511149
transform 1 0 10212 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_7
timestamp 1644511149
transform 1 0 1748 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_11
timestamp 1644511149
transform 1 0 2116 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_15
timestamp 1644511149
transform 1 0 2484 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_24
timestamp 1644511149
transform 1 0 3312 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_33
timestamp 1644511149
transform 1 0 4140 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_45
timestamp 1644511149
transform 1 0 5244 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_53
timestamp 1644511149
transform 1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1644511149
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1644511149
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1644511149
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_93
timestamp 1644511149
transform 1 0 9660 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_99
timestamp 1644511149
transform 1 0 10212 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_7
timestamp 1644511149
transform 1 0 1748 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1644511149
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1644511149
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1644511149
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_41
timestamp 1644511149
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_53
timestamp 1644511149
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_65
timestamp 1644511149
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1644511149
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1644511149
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_85
timestamp 1644511149
transform 1 0 8924 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_93
timestamp 1644511149
transform 1 0 9660 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_99
timestamp 1644511149
transform 1 0 10212 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_7
timestamp 1644511149
transform 1 0 1748 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_16
timestamp 1644511149
transform 1 0 2576 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_20
timestamp 1644511149
transform 1 0 2944 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_26
timestamp 1644511149
transform 1 0 3496 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_38
timestamp 1644511149
transform 1 0 4600 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_50
timestamp 1644511149
transform 1 0 5704 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1644511149
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1644511149
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_81
timestamp 1644511149
transform 1 0 8556 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_87
timestamp 1644511149
transform 1 0 9108 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_91
timestamp 1644511149
transform 1 0 9476 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_99
timestamp 1644511149
transform 1 0 10212 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_7
timestamp 1644511149
transform 1 0 1748 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_19
timestamp 1644511149
transform 1 0 2852 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1644511149
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1644511149
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1644511149
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_53
timestamp 1644511149
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1644511149
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1644511149
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1644511149
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_85
timestamp 1644511149
transform 1 0 8924 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_93
timestamp 1644511149
transform 1 0 9660 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_99
timestamp 1644511149
transform 1 0 10212 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_7
timestamp 1644511149
transform 1 0 1748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_15
timestamp 1644511149
transform 1 0 2484 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_22
timestamp 1644511149
transform 1 0 3128 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_34
timestamp 1644511149
transform 1 0 4232 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_46
timestamp 1644511149
transform 1 0 5336 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1644511149
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1644511149
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1644511149
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_81
timestamp 1644511149
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_93
timestamp 1644511149
transform 1 0 9660 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_99
timestamp 1644511149
transform 1 0 10212 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_10
timestamp 1644511149
transform 1 0 2024 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_18
timestamp 1644511149
transform 1 0 2760 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_26
timestamp 1644511149
transform 1 0 3496 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1644511149
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1644511149
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1644511149
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1644511149
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1644511149
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1644511149
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_85
timestamp 1644511149
transform 1 0 8924 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_96_93
timestamp 1644511149
transform 1 0 9660 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_99
timestamp 1644511149
transform 1 0 10212 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_11
timestamp 1644511149
transform 1 0 2116 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_19
timestamp 1644511149
transform 1 0 2852 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1644511149
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1644511149
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1644511149
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1644511149
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1644511149
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1644511149
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_81
timestamp 1644511149
transform 1 0 8556 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_97_99
timestamp 1644511149
transform 1 0 10212 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_7
timestamp 1644511149
transform 1 0 1748 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_13
timestamp 1644511149
transform 1 0 2300 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_19
timestamp 1644511149
transform 1 0 2852 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1644511149
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_34
timestamp 1644511149
transform 1 0 4232 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_42
timestamp 1644511149
transform 1 0 4968 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_54
timestamp 1644511149
transform 1 0 6072 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_66
timestamp 1644511149
transform 1 0 7176 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_78
timestamp 1644511149
transform 1 0 8280 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_85
timestamp 1644511149
transform 1 0 8924 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_99
timestamp 1644511149
transform 1 0 10212 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_3
timestamp 1644511149
transform 1 0 1380 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_12
timestamp 1644511149
transform 1 0 2208 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_22
timestamp 1644511149
transform 1 0 3128 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_31
timestamp 1644511149
transform 1 0 3956 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_43
timestamp 1644511149
transform 1 0 5060 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1644511149
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_57
timestamp 1644511149
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_69
timestamp 1644511149
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_81
timestamp 1644511149
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_93
timestamp 1644511149
transform 1 0 9660 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_99
timestamp 1644511149
transform 1 0 10212 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_11
timestamp 1644511149
transform 1 0 2116 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_15
timestamp 1644511149
transform 1 0 2484 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_21
timestamp 1644511149
transform 1 0 3036 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1644511149
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_32
timestamp 1644511149
transform 1 0 4048 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_44
timestamp 1644511149
transform 1 0 5152 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_56
timestamp 1644511149
transform 1 0 6256 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_68
timestamp 1644511149
transform 1 0 7360 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_80
timestamp 1644511149
transform 1 0 8464 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_85
timestamp 1644511149
transform 1 0 8924 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_99
timestamp 1644511149
transform 1 0 10212 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_7
timestamp 1644511149
transform 1 0 1748 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_15
timestamp 1644511149
transform 1 0 2484 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_23
timestamp 1644511149
transform 1 0 3220 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_30
timestamp 1644511149
transform 1 0 3864 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_42
timestamp 1644511149
transform 1 0 4968 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_54
timestamp 1644511149
transform 1 0 6072 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1644511149
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1644511149
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_81
timestamp 1644511149
transform 1 0 8556 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_99
timestamp 1644511149
transform 1 0 10212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_102_11
timestamp 1644511149
transform 1 0 2116 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_102_23
timestamp 1644511149
transform 1 0 3220 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1644511149
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_29
timestamp 1644511149
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_41
timestamp 1644511149
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_53
timestamp 1644511149
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_65
timestamp 1644511149
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1644511149
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1644511149
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_85
timestamp 1644511149
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_97
timestamp 1644511149
transform 1 0 10028 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_103_3
timestamp 1644511149
transform 1 0 1380 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_7
timestamp 1644511149
transform 1 0 1748 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_16
timestamp 1644511149
transform 1 0 2576 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_28
timestamp 1644511149
transform 1 0 3680 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_40
timestamp 1644511149
transform 1 0 4784 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_52
timestamp 1644511149
transform 1 0 5888 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_57
timestamp 1644511149
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_69
timestamp 1644511149
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_81
timestamp 1644511149
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_103_93
timestamp 1644511149
transform 1 0 9660 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_103_99
timestamp 1644511149
transform 1 0 10212 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_7
timestamp 1644511149
transform 1 0 1748 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_15
timestamp 1644511149
transform 1 0 2484 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_23
timestamp 1644511149
transform 1 0 3220 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1644511149
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_29
timestamp 1644511149
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_41
timestamp 1644511149
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_53
timestamp 1644511149
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_65
timestamp 1644511149
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1644511149
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1644511149
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_85
timestamp 1644511149
transform 1 0 8924 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_104_93
timestamp 1644511149
transform 1 0 9660 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_104_99
timestamp 1644511149
transform 1 0 10212 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_7
timestamp 1644511149
transform 1 0 1748 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_19
timestamp 1644511149
transform 1 0 2852 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_31
timestamp 1644511149
transform 1 0 3956 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_43
timestamp 1644511149
transform 1 0 5060 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1644511149
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_57
timestamp 1644511149
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_69
timestamp 1644511149
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_81
timestamp 1644511149
transform 1 0 8556 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_105_99
timestamp 1644511149
transform 1 0 10212 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_7
timestamp 1644511149
transform 1 0 1748 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_15
timestamp 1644511149
transform 1 0 2484 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_22
timestamp 1644511149
transform 1 0 3128 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1644511149
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1644511149
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_53
timestamp 1644511149
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_65
timestamp 1644511149
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1644511149
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1644511149
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_85
timestamp 1644511149
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_97
timestamp 1644511149
transform 1 0 10028 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_107_11
timestamp 1644511149
transform 1 0 2116 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_19
timestamp 1644511149
transform 1 0 2852 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_31
timestamp 1644511149
transform 1 0 3956 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_43
timestamp 1644511149
transform 1 0 5060 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1644511149
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_57
timestamp 1644511149
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_69
timestamp 1644511149
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_81
timestamp 1644511149
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_107_93
timestamp 1644511149
transform 1 0 9660 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_99
timestamp 1644511149
transform 1 0 10212 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_7
timestamp 1644511149
transform 1 0 1748 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_108_15
timestamp 1644511149
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1644511149
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_29
timestamp 1644511149
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_41
timestamp 1644511149
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_53
timestamp 1644511149
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_65
timestamp 1644511149
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1644511149
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1644511149
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_85
timestamp 1644511149
transform 1 0 8924 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_108_93
timestamp 1644511149
transform 1 0 9660 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_99
timestamp 1644511149
transform 1 0 10212 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_109_11
timestamp 1644511149
transform 1 0 2116 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_23
timestamp 1644511149
transform 1 0 3220 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_35
timestamp 1644511149
transform 1 0 4324 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_47
timestamp 1644511149
transform 1 0 5428 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1644511149
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_57
timestamp 1644511149
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_69
timestamp 1644511149
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_81
timestamp 1644511149
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_93
timestamp 1644511149
transform 1 0 9660 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_101
timestamp 1644511149
transform 1 0 10396 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_110_7
timestamp 1644511149
transform 1 0 1748 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_15
timestamp 1644511149
transform 1 0 2484 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_23
timestamp 1644511149
transform 1 0 3220 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1644511149
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_29
timestamp 1644511149
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_41
timestamp 1644511149
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_53
timestamp 1644511149
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_65
timestamp 1644511149
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1644511149
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1644511149
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_85
timestamp 1644511149
transform 1 0 8924 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_110_93
timestamp 1644511149
transform 1 0 9660 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_110_99
timestamp 1644511149
transform 1 0 10212 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_111_11
timestamp 1644511149
transform 1 0 2116 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_111_22
timestamp 1644511149
transform 1 0 3128 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_30
timestamp 1644511149
transform 1 0 3864 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_42
timestamp 1644511149
transform 1 0 4968 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_54
timestamp 1644511149
transform 1 0 6072 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_111_57
timestamp 1644511149
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_69
timestamp 1644511149
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_81
timestamp 1644511149
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_93
timestamp 1644511149
transform 1 0 9660 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_111_99
timestamp 1644511149
transform 1 0 10212 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_112_3
timestamp 1644511149
transform 1 0 1380 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_112_17
timestamp 1644511149
transform 1 0 2668 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_112_25
timestamp 1644511149
transform 1 0 3404 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_33
timestamp 1644511149
transform 1 0 4140 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_45
timestamp 1644511149
transform 1 0 5244 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_57
timestamp 1644511149
transform 1 0 6348 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_69
timestamp 1644511149
transform 1 0 7452 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_112_81
timestamp 1644511149
transform 1 0 8556 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_112_85
timestamp 1644511149
transform 1 0 8924 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_99
timestamp 1644511149
transform 1 0 10212 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_113_3
timestamp 1644511149
transform 1 0 1380 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_113_17
timestamp 1644511149
transform 1 0 2668 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_29
timestamp 1644511149
transform 1 0 3772 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_41
timestamp 1644511149
transform 1 0 4876 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_113_53
timestamp 1644511149
transform 1 0 5980 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_113_57
timestamp 1644511149
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_69
timestamp 1644511149
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_81
timestamp 1644511149
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_93
timestamp 1644511149
transform 1 0 9660 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_113_101
timestamp 1644511149
transform 1 0 10396 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_114_3
timestamp 1644511149
transform 1 0 1380 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_114_17
timestamp 1644511149
transform 1 0 2668 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_114_25
timestamp 1644511149
transform 1 0 3404 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_114_29
timestamp 1644511149
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_41
timestamp 1644511149
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_53
timestamp 1644511149
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_65
timestamp 1644511149
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1644511149
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1644511149
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_85
timestamp 1644511149
transform 1 0 8924 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_114_93
timestamp 1644511149
transform 1 0 9660 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_114_99
timestamp 1644511149
transform 1 0 10212 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_7
timestamp 1644511149
transform 1 0 1748 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_15
timestamp 1644511149
transform 1 0 2484 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_23
timestamp 1644511149
transform 1 0 3220 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_115_31
timestamp 1644511149
transform 1 0 3956 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_43
timestamp 1644511149
transform 1 0 5060 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1644511149
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_57
timestamp 1644511149
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_69
timestamp 1644511149
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_81
timestamp 1644511149
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_115_93
timestamp 1644511149
transform 1 0 9660 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_115_99
timestamp 1644511149
transform 1 0 10212 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_13
timestamp 1644511149
transform 1 0 2300 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_23
timestamp 1644511149
transform 1 0 3220 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1644511149
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_33
timestamp 1644511149
transform 1 0 4140 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_45
timestamp 1644511149
transform 1 0 5244 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_57
timestamp 1644511149
transform 1 0 6348 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_69
timestamp 1644511149
transform 1 0 7452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_116_81
timestamp 1644511149
transform 1 0 8556 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_85
timestamp 1644511149
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_97
timestamp 1644511149
transform 1 0 10028 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_117_13
timestamp 1644511149
transform 1 0 2300 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_117_25
timestamp 1644511149
transform 1 0 3404 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_37
timestamp 1644511149
transform 1 0 4508 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_49
timestamp 1644511149
transform 1 0 5612 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_55
timestamp 1644511149
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_57
timestamp 1644511149
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_69
timestamp 1644511149
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_81
timestamp 1644511149
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_93
timestamp 1644511149
transform 1 0 9660 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_117_99
timestamp 1644511149
transform 1 0 10212 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_13
timestamp 1644511149
transform 1 0 2300 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_17
timestamp 1644511149
transform 1 0 2668 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_118_24
timestamp 1644511149
transform 1 0 3312 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_118_29
timestamp 1644511149
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_41
timestamp 1644511149
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_53
timestamp 1644511149
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_65
timestamp 1644511149
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1644511149
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1644511149
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_85
timestamp 1644511149
transform 1 0 8924 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_93
timestamp 1644511149
transform 1 0 9660 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_118_99
timestamp 1644511149
transform 1 0 10212 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_13
timestamp 1644511149
transform 1 0 2300 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_119_25
timestamp 1644511149
transform 1 0 3404 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_37
timestamp 1644511149
transform 1 0 4508 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_49
timestamp 1644511149
transform 1 0 5612 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1644511149
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_57
timestamp 1644511149
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_69
timestamp 1644511149
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_81
timestamp 1644511149
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_93
timestamp 1644511149
transform 1 0 9660 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_99
timestamp 1644511149
transform 1 0 10212 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_120_6
timestamp 1644511149
transform 1 0 1656 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_120_20
timestamp 1644511149
transform 1 0 2944 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_120_29
timestamp 1644511149
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_41
timestamp 1644511149
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_53
timestamp 1644511149
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_65
timestamp 1644511149
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1644511149
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1644511149
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_85
timestamp 1644511149
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_97
timestamp 1644511149
transform 1 0 10028 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_121_11
timestamp 1644511149
transform 1 0 2116 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_18
timestamp 1644511149
transform 1 0 2760 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_30
timestamp 1644511149
transform 1 0 3864 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_42
timestamp 1644511149
transform 1 0 4968 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_121_54
timestamp 1644511149
transform 1 0 6072 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_121_57
timestamp 1644511149
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_69
timestamp 1644511149
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_81
timestamp 1644511149
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_121_93
timestamp 1644511149
transform 1 0 9660 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_121_99
timestamp 1644511149
transform 1 0 10212 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_122_11
timestamp 1644511149
transform 1 0 2116 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_122_18
timestamp 1644511149
transform 1 0 2760 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_122_26
timestamp 1644511149
transform 1 0 3496 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_122_29
timestamp 1644511149
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_41
timestamp 1644511149
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_53
timestamp 1644511149
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_65
timestamp 1644511149
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1644511149
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1644511149
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_85
timestamp 1644511149
transform 1 0 8924 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_93
timestamp 1644511149
transform 1 0 9660 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_99
timestamp 1644511149
transform 1 0 10212 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_6
timestamp 1644511149
transform 1 0 1656 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_123_13
timestamp 1644511149
transform 1 0 2300 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_25
timestamp 1644511149
transform 1 0 3404 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_37
timestamp 1644511149
transform 1 0 4508 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_49
timestamp 1644511149
transform 1 0 5612 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1644511149
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_57
timestamp 1644511149
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_69
timestamp 1644511149
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_81
timestamp 1644511149
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_93
timestamp 1644511149
transform 1 0 9660 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_123_101
timestamp 1644511149
transform 1 0 10396 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_124_6
timestamp 1644511149
transform 1 0 1656 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_124_13
timestamp 1644511149
transform 1 0 2300 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_124_25
timestamp 1644511149
transform 1 0 3404 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_124_29
timestamp 1644511149
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_41
timestamp 1644511149
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_53
timestamp 1644511149
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_65
timestamp 1644511149
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1644511149
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1644511149
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_85
timestamp 1644511149
transform 1 0 8924 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_124_93
timestamp 1644511149
transform 1 0 9660 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_124_99
timestamp 1644511149
transform 1 0 10212 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_125_11
timestamp 1644511149
transform 1 0 2116 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_23
timestamp 1644511149
transform 1 0 3220 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_35
timestamp 1644511149
transform 1 0 4324 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_47
timestamp 1644511149
transform 1 0 5428 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1644511149
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_57
timestamp 1644511149
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_69
timestamp 1644511149
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_81
timestamp 1644511149
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_125_93
timestamp 1644511149
transform 1 0 9660 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_125_99
timestamp 1644511149
transform 1 0 10212 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_126_6
timestamp 1644511149
transform 1 0 1656 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_126_13
timestamp 1644511149
transform 1 0 2300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_126_25
timestamp 1644511149
transform 1 0 3404 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_126_29
timestamp 1644511149
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_41
timestamp 1644511149
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_53
timestamp 1644511149
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_65
timestamp 1644511149
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1644511149
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1644511149
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_85
timestamp 1644511149
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_97
timestamp 1644511149
transform 1 0 10028 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_127_11
timestamp 1644511149
transform 1 0 2116 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_127_23
timestamp 1644511149
transform 1 0 3220 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_35
timestamp 1644511149
transform 1 0 4324 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_47
timestamp 1644511149
transform 1 0 5428 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1644511149
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_57
timestamp 1644511149
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_69
timestamp 1644511149
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_81
timestamp 1644511149
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_93
timestamp 1644511149
transform 1 0 9660 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_127_99
timestamp 1644511149
transform 1 0 10212 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_128_6
timestamp 1644511149
transform 1 0 1656 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_128_18
timestamp 1644511149
transform 1 0 2760 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_128_26
timestamp 1644511149
transform 1 0 3496 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_128_29
timestamp 1644511149
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_41
timestamp 1644511149
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_53
timestamp 1644511149
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_65
timestamp 1644511149
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1644511149
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1644511149
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_85
timestamp 1644511149
transform 1 0 8924 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_128_93
timestamp 1644511149
transform 1 0 9660 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_128_99
timestamp 1644511149
transform 1 0 10212 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_129_6
timestamp 1644511149
transform 1 0 1656 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_129_13
timestamp 1644511149
transform 1 0 2300 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_129_20
timestamp 1644511149
transform 1 0 2944 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_32
timestamp 1644511149
transform 1 0 4048 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_44
timestamp 1644511149
transform 1 0 5152 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_57
timestamp 1644511149
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_69
timestamp 1644511149
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_81
timestamp 1644511149
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_129_93
timestamp 1644511149
transform 1 0 9660 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_129_99
timestamp 1644511149
transform 1 0 10212 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_130_11
timestamp 1644511149
transform 1 0 2116 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_130_23
timestamp 1644511149
transform 1 0 3220 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 1644511149
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_29
timestamp 1644511149
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_41
timestamp 1644511149
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_53
timestamp 1644511149
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_65
timestamp 1644511149
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1644511149
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1644511149
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_85
timestamp 1644511149
transform 1 0 8924 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_97
timestamp 1644511149
transform 1 0 10028 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_131_6
timestamp 1644511149
transform 1 0 1656 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_131_13
timestamp 1644511149
transform 1 0 2300 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_25
timestamp 1644511149
transform 1 0 3404 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_37
timestamp 1644511149
transform 1 0 4508 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_49
timestamp 1644511149
transform 1 0 5612 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_55
timestamp 1644511149
transform 1 0 6164 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_57
timestamp 1644511149
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_69
timestamp 1644511149
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_81
timestamp 1644511149
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_131_93
timestamp 1644511149
transform 1 0 9660 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_131_99
timestamp 1644511149
transform 1 0 10212 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_132_3
timestamp 1644511149
transform 1 0 1380 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_132_17
timestamp 1644511149
transform 1 0 2668 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_132_24
timestamp 1644511149
transform 1 0 3312 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_132_29
timestamp 1644511149
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_41
timestamp 1644511149
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_53
timestamp 1644511149
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_65
timestamp 1644511149
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1644511149
transform 1 0 8188 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1644511149
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_85
timestamp 1644511149
transform 1 0 8924 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_132_93
timestamp 1644511149
transform 1 0 9660 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_132_99
timestamp 1644511149
transform 1 0 10212 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_133_11
timestamp 1644511149
transform 1 0 2116 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_133_18
timestamp 1644511149
transform 1 0 2760 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_30
timestamp 1644511149
transform 1 0 3864 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_42
timestamp 1644511149
transform 1 0 4968 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_133_54
timestamp 1644511149
transform 1 0 6072 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_133_57
timestamp 1644511149
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_69
timestamp 1644511149
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_81
timestamp 1644511149
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_93
timestamp 1644511149
transform 1 0 9660 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_133_101
timestamp 1644511149
transform 1 0 10396 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_134_3
timestamp 1644511149
transform 1 0 1380 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_134_17
timestamp 1644511149
transform 1 0 2668 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_134_24
timestamp 1644511149
transform 1 0 3312 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_134_29
timestamp 1644511149
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_41
timestamp 1644511149
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_53
timestamp 1644511149
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_65
timestamp 1644511149
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1644511149
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1644511149
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_85
timestamp 1644511149
transform 1 0 8924 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_134_93
timestamp 1644511149
transform 1 0 9660 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_134_99
timestamp 1644511149
transform 1 0 10212 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_135_6
timestamp 1644511149
transform 1 0 1656 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_12
timestamp 1644511149
transform 1 0 2208 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_135_21
timestamp 1644511149
transform 1 0 3036 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_28
timestamp 1644511149
transform 1 0 3680 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_40
timestamp 1644511149
transform 1 0 4784 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_52
timestamp 1644511149
transform 1 0 5888 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_57
timestamp 1644511149
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_69
timestamp 1644511149
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_81
timestamp 1644511149
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_135_93
timestamp 1644511149
transform 1 0 9660 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_135_99
timestamp 1644511149
transform 1 0 10212 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_136_11
timestamp 1644511149
transform 1 0 2116 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_136_23
timestamp 1644511149
transform 1 0 3220 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 1644511149
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_29
timestamp 1644511149
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_41
timestamp 1644511149
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_53
timestamp 1644511149
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_65
timestamp 1644511149
transform 1 0 7084 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1644511149
transform 1 0 8188 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1644511149
transform 1 0 8740 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_85
timestamp 1644511149
transform 1 0 8924 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_136_93
timestamp 1644511149
transform 1 0 9660 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_136_99
timestamp 1644511149
transform 1 0 10212 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_7
timestamp 1644511149
transform 1 0 1748 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_14
timestamp 1644511149
transform 1 0 2392 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_21
timestamp 1644511149
transform 1 0 3036 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_28
timestamp 1644511149
transform 1 0 3680 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_137_35
timestamp 1644511149
transform 1 0 4324 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_47
timestamp 1644511149
transform 1 0 5428 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1644511149
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_57
timestamp 1644511149
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_69
timestamp 1644511149
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_81
timestamp 1644511149
transform 1 0 8556 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_87
timestamp 1644511149
transform 1 0 9108 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_137_91
timestamp 1644511149
transform 1 0 9476 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_99
timestamp 1644511149
transform 1 0 10212 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_13
timestamp 1644511149
transform 1 0 2300 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_138_20
timestamp 1644511149
transform 1 0 2944 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_138_32
timestamp 1644511149
transform 1 0 4048 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_138_39
timestamp 1644511149
transform 1 0 4692 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_138_51
timestamp 1644511149
transform 1 0 5796 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_55
timestamp 1644511149
transform 1 0 6164 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_57
timestamp 1644511149
transform 1 0 6348 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_69
timestamp 1644511149
transform 1 0 7452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1644511149
transform 1 0 8556 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_138_85
timestamp 1644511149
transform 1 0 8924 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_91
timestamp 1644511149
transform 1 0 9476 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_99
timestamp 1644511149
transform 1 0 10212 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 10856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 10856 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 10856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 10856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 10856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 10856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 10856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 10856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 10856 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 10856 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 10856 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 10856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 10856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 10856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 10856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 10856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 10856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 10856 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 10856 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 10856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 10856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 10856 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 10856 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 10856 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 10856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 10856 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 10856 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 10856 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 10856 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 10856 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 10856 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 10856 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 10856 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 10856 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 10856 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 10856 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 10856 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 10856 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 10856 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 10856 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 10856 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 10856 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 10856 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 10856 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 10856 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 10856 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 10856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 10856 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 10856 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 10856 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 10856 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 10856 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1644511149
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1644511149
transform -1 0 10856 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1644511149
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1644511149
transform -1 0 10856 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1644511149
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1644511149
transform -1 0 10856 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1644511149
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1644511149
transform -1 0 10856 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1644511149
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1644511149
transform -1 0 10856 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1644511149
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1644511149
transform -1 0 10856 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1644511149
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1644511149
transform -1 0 10856 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1644511149
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1644511149
transform -1 0 10856 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1644511149
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1644511149
transform -1 0 10856 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1644511149
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1644511149
transform -1 0 10856 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1644511149
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1644511149
transform -1 0 10856 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1644511149
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1644511149
transform -1 0 10856 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1644511149
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1644511149
transform -1 0 10856 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1644511149
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1644511149
transform -1 0 10856 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1644511149
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1644511149
transform -1 0 10856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1644511149
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1644511149
transform -1 0 10856 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1644511149
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1644511149
transform -1 0 10856 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1644511149
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1644511149
transform -1 0 10856 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1644511149
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1644511149
transform -1 0 10856 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1644511149
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1644511149
transform -1 0 10856 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1644511149
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1644511149
transform -1 0 10856 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1644511149
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1644511149
transform -1 0 10856 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1644511149
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1644511149
transform -1 0 10856 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1644511149
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1644511149
transform -1 0 10856 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1644511149
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1644511149
transform -1 0 10856 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1644511149
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1644511149
transform -1 0 10856 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1644511149
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1644511149
transform -1 0 10856 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1644511149
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1644511149
transform -1 0 10856 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1644511149
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1644511149
transform -1 0 10856 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1644511149
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1644511149
transform -1 0 10856 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1644511149
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1644511149
transform -1 0 10856 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1644511149
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1644511149
transform -1 0 10856 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1644511149
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1644511149
transform -1 0 10856 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1644511149
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1644511149
transform -1 0 10856 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1644511149
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1644511149
transform -1 0 10856 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1644511149
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1644511149
transform -1 0 10856 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1644511149
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1644511149
transform -1 0 10856 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1644511149
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1644511149
transform -1 0 10856 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1644511149
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1644511149
transform -1 0 10856 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1644511149
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1644511149
transform -1 0 10856 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1644511149
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1644511149
transform -1 0 10856 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1644511149
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1644511149
transform -1 0 10856 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1644511149
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1644511149
transform -1 0 10856 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1644511149
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1644511149
transform -1 0 10856 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1644511149
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1644511149
transform -1 0 10856 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1644511149
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1644511149
transform -1 0 10856 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1644511149
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1644511149
transform -1 0 10856 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1644511149
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1644511149
transform -1 0 10856 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1644511149
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1644511149
transform -1 0 10856 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1644511149
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1644511149
transform -1 0 10856 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1644511149
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1644511149
transform -1 0 10856 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1644511149
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1644511149
transform -1 0 10856 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__or4bb_1  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _096_
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _100_
timestamp 1644511149
transform 1 0 2668 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  _102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2852 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1656 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _106_
timestamp 1644511149
transform 1 0 1656 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1644511149
transform 1 0 2668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _108_
timestamp 1644511149
transform 1 0 2668 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1644511149
transform 1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _110_
timestamp 1644511149
transform 1 0 2668 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1644511149
transform 1 0 4140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _112_
timestamp 1644511149
transform 1 0 2668 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1644511149
transform 1 0 2668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _114_
timestamp 1644511149
transform 1 0 2116 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1644511149
transform 1 0 1932 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _116_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1644511149
transform 1 0 1472 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _118_
timestamp 1644511149
transform 1 0 1656 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _120_
timestamp 1644511149
transform 1 0 2116 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1644511149
transform 1 0 2944 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _122_
timestamp 1644511149
transform 1 0 1748 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1644511149
transform 1 0 1656 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _124_
timestamp 1644511149
transform 1 0 1748 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1644511149
transform 1 0 1748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _126_
timestamp 1644511149
transform 1 0 2208 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1644511149
transform 1 0 2024 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _128_
timestamp 1644511149
transform 1 0 2576 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _130_
timestamp 1644511149
transform 1 0 1472 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1472 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _132_
timestamp 1644511149
transform 1 0 2300 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _133_
timestamp 1644511149
transform 1 0 1472 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2760 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _135_
timestamp 1644511149
transform 1 0 2300 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1644511149
transform 1 0 3128 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _137_
timestamp 1644511149
transform 1 0 2024 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1644511149
transform 1 0 1564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _139_
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _140_
timestamp 1644511149
transform 1 0 2392 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _141_
timestamp 1644511149
transform 1 0 2024 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _142_
timestamp 1644511149
transform 1 0 2116 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _143_
timestamp 1644511149
transform 1 0 1748 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _144_
timestamp 1644511149
transform 1 0 1472 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _145_
timestamp 1644511149
transform 1 0 1472 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _146_
timestamp 1644511149
transform 1 0 1472 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _147_
timestamp 1644511149
transform 1 0 2300 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _148_
timestamp 1644511149
transform 1 0 1656 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _149_
timestamp 1644511149
transform 1 0 2024 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _150_
timestamp 1644511149
transform 1 0 1932 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _151_
timestamp 1644511149
transform 1 0 2392 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _152_
timestamp 1644511149
transform 1 0 2392 0 1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _153_
timestamp 1644511149
transform 1 0 1564 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _154_
timestamp 1644511149
transform 1 0 2576 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _155_
timestamp 1644511149
transform 1 0 1564 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1644511149
transform 1 0 1656 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _157_
timestamp 1644511149
transform 1 0 2392 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3128 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _159_
timestamp 1644511149
transform 1 0 2116 0 -1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1644511149
transform 1 0 2852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _161_
timestamp 1644511149
transform 1 0 2392 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1644511149
transform 1 0 2208 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _163_
timestamp 1644511149
transform 1 0 2392 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1644511149
transform 1 0 3588 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _165_
timestamp 1644511149
transform 1 0 2576 0 1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1644511149
transform 1 0 2852 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _167_
timestamp 1644511149
transform 1 0 1748 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1644511149
transform 1 0 3772 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _169_
timestamp 1644511149
transform 1 0 2576 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2116 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_4  _171_
timestamp 1644511149
transform 1 0 2668 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 -1 63104
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _173_
timestamp 1644511149
transform 1 0 1380 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _174_
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _175_
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _176_
timestamp 1644511149
transform 1 0 1380 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _178_
timestamp 1644511149
transform 1 0 1380 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _179_
timestamp 1644511149
transform 1 0 1380 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _180_
timestamp 1644511149
transform 1 0 1380 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _181_
timestamp 1644511149
transform 1 0 1380 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _182_
timestamp 1644511149
transform 1 0 1380 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _183_
timestamp 1644511149
transform 1 0 1380 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _184_
timestamp 1644511149
transform 1 0 1840 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _185_
timestamp 1644511149
transform 1 0 1932 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _186_
timestamp 1644511149
transform 1 0 1932 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _187_
timestamp 1644511149
transform 1 0 1932 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _188_
timestamp 1644511149
transform 1 0 2668 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _189_
timestamp 1644511149
transform 1 0 2760 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _190_
timestamp 1644511149
transform 1 0 2668 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _191_
timestamp 1644511149
transform 1 0 2208 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _192_
timestamp 1644511149
transform 1 0 2668 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _193_
timestamp 1644511149
transform 1 0 1380 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _194_
timestamp 1644511149
transform 1 0 1380 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _195_
timestamp 1644511149
transform 1 0 1380 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _196_
timestamp 1644511149
transform 1 0 1380 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _197_
timestamp 1644511149
transform 1 0 1380 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _198_
timestamp 1644511149
transform 1 0 2484 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _199_
timestamp 1644511149
transform 1 0 2024 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _200_
timestamp 1644511149
transform 1 0 1932 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _201_
timestamp 1644511149
transform 1 0 1932 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _202_
timestamp 1644511149
transform 1 0 2300 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _203_
timestamp 1644511149
transform 1 0 1380 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _204_
timestamp 1644511149
transform 1 0 1380 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _205_
timestamp 1644511149
transform 1 0 2484 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _206_
timestamp 1644511149
transform 1 0 2852 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _207_
timestamp 1644511149
transform 1 0 2760 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _208_
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _210_
timestamp 1644511149
transform 1 0 2576 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 1644511149
transform 1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _212_
timestamp 1644511149
transform 1 0 3404 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1644511149
transform 1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _214_
timestamp 1644511149
transform 1 0 4232 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1644511149
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _216_
timestamp 1644511149
transform 1 0 2392 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1644511149
transform 1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _218_
timestamp 1644511149
transform 1 0 3312 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1644511149
transform 1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _220_
timestamp 1644511149
transform 1 0 2668 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1644511149
transform 1 0 2852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _222_
timestamp 1644511149
transform 1 0 2576 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1644511149
transform 1 0 5060 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _224_
timestamp 1644511149
transform 1 0 2576 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _225_
timestamp 1644511149
transform 1 0 3772 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _226_
timestamp 1644511149
transform 1 0 2392 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _227_
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _228_
timestamp 1644511149
transform 1 0 2392 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _230_
timestamp 1644511149
transform 1 0 2576 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1644511149
transform 1 0 4232 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _232_
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _233_
timestamp 1644511149
transform 1 0 3772 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _234_
timestamp 1644511149
transform 1 0 2760 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _235_
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _236_
timestamp 1644511149
transform 1 0 2576 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 1644511149
transform 1 0 4508 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _238_
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _239_
timestamp 1644511149
transform 1 0 5060 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _241_
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1644511149
transform 1 0 6992 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _243_
timestamp 1644511149
transform 1 0 4968 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _245_
timestamp 1644511149
transform 1 0 5336 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1644511149
transform 1 0 9844 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _247_
timestamp 1644511149
transform 1 0 5244 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1644511149
transform 1 0 9200 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _249_
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1644511149
transform 1 0 6624 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _251_
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1644511149
transform 1 0 9200 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _253_
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1644511149
transform 1 0 9936 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _255_
timestamp 1644511149
transform 1 0 4692 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1644511149
transform 1 0 9936 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _257_
timestamp 1644511149
transform 1 0 4968 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _258_
timestamp 1644511149
transform 1 0 6256 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _259_
timestamp 1644511149
transform 1 0 4508 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _261_
timestamp 1644511149
transform 1 0 4968 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _263_
timestamp 1644511149
transform 1 0 5796 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1644511149
transform 1 0 6624 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _265_
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _266_
timestamp 1644511149
transform 1 0 7820 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _267_
timestamp 1644511149
transform 1 0 5520 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp 1644511149
transform 1 0 7728 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _269_
timestamp 1644511149
transform 1 0 4508 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _270_
timestamp 1644511149
transform 1 0 9936 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _271_
timestamp 1644511149
transform 1 0 2760 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 1644511149
transform 1 0 9200 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _273_
timestamp 1644511149
transform 1 0 2760 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1644511149
transform 1 0 9936 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _275_
timestamp 1644511149
transform 1 0 2852 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1644511149
transform 1 0 9936 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _277_
timestamp 1644511149
transform 1 0 3680 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _278_
timestamp 1644511149
transform 1 0 9936 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _279_
timestamp 1644511149
transform 1 0 3036 0 -1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp 1644511149
transform 1 0 9200 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _281_
timestamp 1644511149
transform 1 0 3496 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1644511149
transform 1 0 9936 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _283_
timestamp 1644511149
transform 1 0 3772 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 1644511149
transform 1 0 9936 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _285_
timestamp 1644511149
transform 1 0 2668 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _286_
timestamp 1644511149
transform 1 0 1840 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _287_
timestamp 1644511149
transform 1 0 1748 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _289_
timestamp 1644511149
transform 1 0 1564 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _290_
timestamp 1644511149
transform 1 0 2668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _291_
timestamp 1644511149
transform 1 0 1932 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _292_
timestamp 1644511149
transform 1 0 2392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _293_
timestamp 1644511149
transform 1 0 2576 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _294_
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _295_
timestamp 1644511149
transform 1 0 2668 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _296_
timestamp 1644511149
transform 1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _297__290 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9936 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _298__291
timestamp 1644511149
transform 1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _299__280
timestamp 1644511149
transform 1 0 9936 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _300__281
timestamp 1644511149
transform 1 0 9936 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _301__282
timestamp 1644511149
transform 1 0 9936 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _302__283
timestamp 1644511149
transform 1 0 9936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _303__284
timestamp 1644511149
transform 1 0 9936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _304__285
timestamp 1644511149
transform 1 0 9936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _305__286
timestamp 1644511149
transform 1 0 9936 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _306__287
timestamp 1644511149
transform 1 0 9936 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _307__288
timestamp 1644511149
transform 1 0 9936 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _308__289
timestamp 1644511149
transform 1 0 9936 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1644511149
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1644511149
transform 1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 1644511149
transform 1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1644511149
transform 1 0 4048 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1644511149
transform 1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp 1644511149
transform 1 0 2668 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1644511149
transform 1 0 3496 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp 1644511149
transform 1 0 2576 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1644511149
transform 1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _321_
timestamp 1644511149
transform 1 0 9200 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1644511149
transform 1 0 9936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1644511149
transform 1 0 9200 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1644511149
transform 1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp 1644511149
transform 1 0 9936 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1644511149
transform 1 0 9844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1644511149
transform 1 0 9200 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1644511149
transform 1 0 9936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _330_
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _331_
timestamp 1644511149
transform 1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _332_
timestamp 1644511149
transform 1 0 2668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _333_
timestamp 1644511149
transform 1 0 2668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _334_
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _335_
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _336_
timestamp 1644511149
transform 1 0 3404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _337_
timestamp 1644511149
transform 1 0 1656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _338_
timestamp 1644511149
transform 1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _339_
timestamp 1644511149
transform 1 0 3036 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _340_
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _341_
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1644511149
transform 1 0 9844 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1644511149
transform 1 0 9292 0 -1 55488
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 9936 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1644511149
transform 1 0 9292 0 1 63104
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 9936 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 9936 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 9936 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 9936 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 9936 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 9936 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 9936 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 9936 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1644511149
transform 1 0 9292 0 1 55488
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 9936 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 9936 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 9936 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 9936 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 9936 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 9936 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 9936 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 9936 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 9936 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 9200 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1644511149
transform 1 0 9292 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 9200 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1644511149
transform 1 0 9844 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1644511149
transform 1 0 9292 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 9936 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 9936 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1644511149
transform 1 0 9292 0 -1 59840
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 9936 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 9936 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 9936 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1644511149
transform 1 0 1380 0 1 77248
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1644511149
transform 1 0 1380 0 -1 66368
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 1380 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 1380 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 2024 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 1380 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 1380 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 2024 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 2668 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 1380 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 2024 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 2484 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1644511149
transform 1 0 1380 0 1 65280
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 3036 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 1380 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 3036 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 3404 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 2116 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform 1 0 2760 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform 1 0 2668 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform 1 0 3772 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1644511149
transform 1 0 3404 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform 1 0 4416 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1644511149
transform 1 0 1380 0 1 66368
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1644511149
transform 1 0 4048 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1644511149
transform 1 0 1380 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1644511149
transform 1 0 1380 0 -1 67456
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1644511149
transform 1 0 1380 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1644511149
transform 1 0 2484 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1644511149
transform 1 0 1380 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1644511149
transform 1 0 2484 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1644511149
transform 1 0 2024 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1644511149
transform 1 0 2024 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input68
timestamp 1644511149
transform 1 0 2668 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1644511149
transform 1 0 3496 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1644511149
transform 1 0 3220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1644511149
transform 1 0 2576 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1644511149
transform 1 0 2668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1644511149
transform 1 0 3404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1644511149
transform 1 0 4416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input94
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input95
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input96
timestamp 1644511149
transform 1 0 2760 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1644511149
transform 1 0 4140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1644511149
transform 1 0 3496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1644511149
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input101
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input102
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input103
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1644511149
transform 1 0 3404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input106
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input107
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1644511149
transform 1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input112
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input113
timestamp 1644511149
transform 1 0 3220 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input114
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1644511149
transform 1 0 2668 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1644511149
transform 1 0 2576 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input117
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 1644511149
transform 1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1644511149
transform 1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1644511149
transform 1 0 3220 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1644511149
transform 1 0 2852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input123
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input124
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1644511149
transform 1 0 3496 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input127
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input128
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input129
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input130
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input131
timestamp 1644511149
transform 1 0 2668 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1644511149
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1644511149
transform 1 0 2668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1644511149
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input137
timestamp 1644511149
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1644511149
transform 1 0 9844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1644511149
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1644511149
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1644511149
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1644511149
transform 1 0 9844 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1644511149
transform 1 0 9844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1644511149
transform 1 0 9844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1644511149
transform 1 0 9844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1644511149
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1644511149
transform 1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1644511149
transform 1 0 9844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1644511149
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1644511149
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1644511149
transform 1 0 9844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1644511149
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1644511149
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1644511149
transform 1 0 9844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1644511149
transform 1 0 9844 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1644511149
transform 1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1644511149
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1644511149
transform 1 0 9844 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1644511149
transform 1 0 9844 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1644511149
transform 1 0 9844 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1644511149
transform 1 0 9844 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1644511149
transform 1 0 9844 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1644511149
transform 1 0 9844 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1644511149
transform 1 0 9844 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1644511149
transform 1 0 9844 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1644511149
transform 1 0 9844 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1644511149
transform 1 0 9844 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1644511149
transform 1 0 9844 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1644511149
transform 1 0 9844 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1644511149
transform 1 0 9844 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1644511149
transform 1 0 9844 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1644511149
transform 1 0 9844 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1644511149
transform 1 0 9844 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1644511149
transform 1 0 9844 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1644511149
transform 1 0 9844 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1644511149
transform 1 0 9844 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1644511149
transform 1 0 9844 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1644511149
transform 1 0 9844 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1644511149
transform 1 0 9844 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1644511149
transform 1 0 9844 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1644511149
transform 1 0 9844 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1644511149
transform 1 0 9844 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1644511149
transform 1 0 9844 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1644511149
transform 1 0 9844 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1644511149
transform 1 0 9844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1644511149
transform 1 0 9844 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1644511149
transform 1 0 9844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1644511149
transform 1 0 9844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1644511149
transform 1 0 9844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1644511149
transform 1 0 9844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1644511149
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1644511149
transform 1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1644511149
transform 1 0 9844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1644511149
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1644511149
transform 1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1644511149
transform 1 0 1380 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1644511149
transform 1 0 3588 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1644511149
transform 1 0 2392 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1644511149
transform 1 0 1380 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1644511149
transform 1 0 2392 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1644511149
transform 1 0 1380 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1644511149
transform 1 0 2116 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1644511149
transform 1 0 1380 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1644511149
transform 1 0 1380 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1644511149
transform 1 0 1380 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1644511149
transform 1 0 1380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1644511149
transform 1 0 2116 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1644511149
transform 1 0 1380 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1644511149
transform 1 0 1380 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1644511149
transform 1 0 2116 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1644511149
transform 1 0 2852 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1644511149
transform 1 0 1380 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1644511149
transform 1 0 2116 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1644511149
transform 1 0 1380 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1644511149
transform 1 0 2116 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1644511149
transform 1 0 2484 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1644511149
transform 1 0 2116 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1644511149
transform 1 0 1380 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1644511149
transform 1 0 2116 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1644511149
transform 1 0 2852 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1644511149
transform 1 0 3496 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1644511149
transform 1 0 3772 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1644511149
transform 1 0 1380 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1644511149
transform 1 0 2116 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1644511149
transform 1 0 2852 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1644511149
transform 1 0 1380 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1644511149
transform 1 0 3588 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1644511149
transform 1 0 3772 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1644511149
transform 1 0 1380 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1644511149
transform 1 0 2116 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1644511149
transform 1 0 2392 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1644511149
transform 1 0 2484 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1644511149
transform 1 0 3220 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1644511149
transform 1 0 4600 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1644511149
transform 1 0 2852 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1644511149
transform 1 0 2852 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1644511149
transform 1 0 3220 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1644511149
transform 1 0 2116 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1644511149
transform 1 0 2760 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1644511149
transform 1 0 2852 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1644511149
transform 1 0 2944 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1644511149
transform 1 0 2760 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1644511149
transform 1 0 3496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1644511149
transform 1 0 2668 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1644511149
transform 1 0 3772 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1644511149
transform 1 0 3312 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1644511149
transform 1 0 2852 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1644511149
transform 1 0 2576 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1644511149
transform 1 0 3404 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1644511149
transform 1 0 3772 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1644511149
transform 1 0 3772 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1644511149
transform 1 0 4508 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1644511149
transform 1 0 2116 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1644511149
transform 1 0 2852 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1644511149
transform 1 0 2116 0 1 34816
box -38 -48 406 592
<< labels >>
rlabel metal4 s 2576 2128 2896 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 5840 2128 6160 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 9104 2128 9424 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 4208 2128 4528 77840 6 vssd1
port 1 nsew ground input
rlabel metal4 s 7472 2128 7792 77840 6 vssd1
port 1 nsew ground input
rlabel metal3 s 0 79568 800 79688 6 wb_clk_i
port 2 nsew signal input
rlabel metal2 s 5998 79200 6054 80000 6 wb_rst_i
port 3 nsew signal input
rlabel metal3 s 11200 79432 12000 79552 6 wbm_a_ack_i
port 4 nsew signal input
rlabel metal3 s 11200 5584 12000 5704 6 wbm_a_adr_o[0]
port 5 nsew signal tristate
rlabel metal3 s 11200 13336 12000 13456 6 wbm_a_adr_o[10]
port 6 nsew signal tristate
rlabel metal3 s 11200 14016 12000 14136 6 wbm_a_adr_o[11]
port 7 nsew signal tristate
rlabel metal3 s 11200 14832 12000 14952 6 wbm_a_adr_o[12]
port 8 nsew signal tristate
rlabel metal3 s 11200 15648 12000 15768 6 wbm_a_adr_o[13]
port 9 nsew signal tristate
rlabel metal3 s 11200 16328 12000 16448 6 wbm_a_adr_o[14]
port 10 nsew signal tristate
rlabel metal3 s 11200 17144 12000 17264 6 wbm_a_adr_o[15]
port 11 nsew signal tristate
rlabel metal3 s 11200 17960 12000 18080 6 wbm_a_adr_o[16]
port 12 nsew signal tristate
rlabel metal3 s 11200 18640 12000 18760 6 wbm_a_adr_o[17]
port 13 nsew signal tristate
rlabel metal3 s 11200 19456 12000 19576 6 wbm_a_adr_o[18]
port 14 nsew signal tristate
rlabel metal3 s 11200 20272 12000 20392 6 wbm_a_adr_o[19]
port 15 nsew signal tristate
rlabel metal3 s 11200 6400 12000 6520 6 wbm_a_adr_o[1]
port 16 nsew signal tristate
rlabel metal3 s 11200 20952 12000 21072 6 wbm_a_adr_o[20]
port 17 nsew signal tristate
rlabel metal3 s 11200 21768 12000 21888 6 wbm_a_adr_o[21]
port 18 nsew signal tristate
rlabel metal3 s 11200 22448 12000 22568 6 wbm_a_adr_o[22]
port 19 nsew signal tristate
rlabel metal3 s 11200 23264 12000 23384 6 wbm_a_adr_o[23]
port 20 nsew signal tristate
rlabel metal3 s 11200 24080 12000 24200 6 wbm_a_adr_o[24]
port 21 nsew signal tristate
rlabel metal3 s 11200 24760 12000 24880 6 wbm_a_adr_o[25]
port 22 nsew signal tristate
rlabel metal3 s 11200 25576 12000 25696 6 wbm_a_adr_o[26]
port 23 nsew signal tristate
rlabel metal3 s 11200 26392 12000 26512 6 wbm_a_adr_o[27]
port 24 nsew signal tristate
rlabel metal3 s 11200 27072 12000 27192 6 wbm_a_adr_o[28]
port 25 nsew signal tristate
rlabel metal3 s 11200 27888 12000 28008 6 wbm_a_adr_o[29]
port 26 nsew signal tristate
rlabel metal3 s 11200 7080 12000 7200 6 wbm_a_adr_o[2]
port 27 nsew signal tristate
rlabel metal3 s 11200 28704 12000 28824 6 wbm_a_adr_o[30]
port 28 nsew signal tristate
rlabel metal3 s 11200 29384 12000 29504 6 wbm_a_adr_o[31]
port 29 nsew signal tristate
rlabel metal3 s 11200 7896 12000 8016 6 wbm_a_adr_o[3]
port 30 nsew signal tristate
rlabel metal3 s 11200 8712 12000 8832 6 wbm_a_adr_o[4]
port 31 nsew signal tristate
rlabel metal3 s 11200 9392 12000 9512 6 wbm_a_adr_o[5]
port 32 nsew signal tristate
rlabel metal3 s 11200 10208 12000 10328 6 wbm_a_adr_o[6]
port 33 nsew signal tristate
rlabel metal3 s 11200 11024 12000 11144 6 wbm_a_adr_o[7]
port 34 nsew signal tristate
rlabel metal3 s 11200 11704 12000 11824 6 wbm_a_adr_o[8]
port 35 nsew signal tristate
rlabel metal3 s 11200 12520 12000 12640 6 wbm_a_adr_o[9]
port 36 nsew signal tristate
rlabel metal3 s 11200 960 12000 1080 6 wbm_a_cyc_o
port 37 nsew signal tristate
rlabel metal3 s 11200 54816 12000 54936 6 wbm_a_dat_i[0]
port 38 nsew signal input
rlabel metal3 s 11200 62432 12000 62552 6 wbm_a_dat_i[10]
port 39 nsew signal input
rlabel metal3 s 11200 63248 12000 63368 6 wbm_a_dat_i[11]
port 40 nsew signal input
rlabel metal3 s 11200 64064 12000 64184 6 wbm_a_dat_i[12]
port 41 nsew signal input
rlabel metal3 s 11200 64744 12000 64864 6 wbm_a_dat_i[13]
port 42 nsew signal input
rlabel metal3 s 11200 65560 12000 65680 6 wbm_a_dat_i[14]
port 43 nsew signal input
rlabel metal3 s 11200 66376 12000 66496 6 wbm_a_dat_i[15]
port 44 nsew signal input
rlabel metal3 s 11200 67056 12000 67176 6 wbm_a_dat_i[16]
port 45 nsew signal input
rlabel metal3 s 11200 67872 12000 67992 6 wbm_a_dat_i[17]
port 46 nsew signal input
rlabel metal3 s 11200 68688 12000 68808 6 wbm_a_dat_i[18]
port 47 nsew signal input
rlabel metal3 s 11200 69368 12000 69488 6 wbm_a_dat_i[19]
port 48 nsew signal input
rlabel metal3 s 11200 55632 12000 55752 6 wbm_a_dat_i[1]
port 49 nsew signal input
rlabel metal3 s 11200 70184 12000 70304 6 wbm_a_dat_i[20]
port 50 nsew signal input
rlabel metal3 s 11200 71000 12000 71120 6 wbm_a_dat_i[21]
port 51 nsew signal input
rlabel metal3 s 11200 71680 12000 71800 6 wbm_a_dat_i[22]
port 52 nsew signal input
rlabel metal3 s 11200 72496 12000 72616 6 wbm_a_dat_i[23]
port 53 nsew signal input
rlabel metal3 s 11200 73312 12000 73432 6 wbm_a_dat_i[24]
port 54 nsew signal input
rlabel metal3 s 11200 73992 12000 74112 6 wbm_a_dat_i[25]
port 55 nsew signal input
rlabel metal3 s 11200 74808 12000 74928 6 wbm_a_dat_i[26]
port 56 nsew signal input
rlabel metal3 s 11200 75624 12000 75744 6 wbm_a_dat_i[27]
port 57 nsew signal input
rlabel metal3 s 11200 76304 12000 76424 6 wbm_a_dat_i[28]
port 58 nsew signal input
rlabel metal3 s 11200 77120 12000 77240 6 wbm_a_dat_i[29]
port 59 nsew signal input
rlabel metal3 s 11200 56312 12000 56432 6 wbm_a_dat_i[2]
port 60 nsew signal input
rlabel metal3 s 11200 77936 12000 78056 6 wbm_a_dat_i[30]
port 61 nsew signal input
rlabel metal3 s 11200 78616 12000 78736 6 wbm_a_dat_i[31]
port 62 nsew signal input
rlabel metal3 s 11200 57128 12000 57248 6 wbm_a_dat_i[3]
port 63 nsew signal input
rlabel metal3 s 11200 57944 12000 58064 6 wbm_a_dat_i[4]
port 64 nsew signal input
rlabel metal3 s 11200 58624 12000 58744 6 wbm_a_dat_i[5]
port 65 nsew signal input
rlabel metal3 s 11200 59440 12000 59560 6 wbm_a_dat_i[6]
port 66 nsew signal input
rlabel metal3 s 11200 60256 12000 60376 6 wbm_a_dat_i[7]
port 67 nsew signal input
rlabel metal3 s 11200 60936 12000 61056 6 wbm_a_dat_i[8]
port 68 nsew signal input
rlabel metal3 s 11200 61752 12000 61872 6 wbm_a_dat_i[9]
port 69 nsew signal input
rlabel metal3 s 11200 30200 12000 30320 6 wbm_a_dat_o[0]
port 70 nsew signal tristate
rlabel metal3 s 11200 37952 12000 38072 6 wbm_a_dat_o[10]
port 71 nsew signal tristate
rlabel metal3 s 11200 38632 12000 38752 6 wbm_a_dat_o[11]
port 72 nsew signal tristate
rlabel metal3 s 11200 39448 12000 39568 6 wbm_a_dat_o[12]
port 73 nsew signal tristate
rlabel metal3 s 11200 40264 12000 40384 6 wbm_a_dat_o[13]
port 74 nsew signal tristate
rlabel metal3 s 11200 40944 12000 41064 6 wbm_a_dat_o[14]
port 75 nsew signal tristate
rlabel metal3 s 11200 41760 12000 41880 6 wbm_a_dat_o[15]
port 76 nsew signal tristate
rlabel metal3 s 11200 42440 12000 42560 6 wbm_a_dat_o[16]
port 77 nsew signal tristate
rlabel metal3 s 11200 43256 12000 43376 6 wbm_a_dat_o[17]
port 78 nsew signal tristate
rlabel metal3 s 11200 44072 12000 44192 6 wbm_a_dat_o[18]
port 79 nsew signal tristate
rlabel metal3 s 11200 44752 12000 44872 6 wbm_a_dat_o[19]
port 80 nsew signal tristate
rlabel metal3 s 11200 31016 12000 31136 6 wbm_a_dat_o[1]
port 81 nsew signal tristate
rlabel metal3 s 11200 45568 12000 45688 6 wbm_a_dat_o[20]
port 82 nsew signal tristate
rlabel metal3 s 11200 46384 12000 46504 6 wbm_a_dat_o[21]
port 83 nsew signal tristate
rlabel metal3 s 11200 47064 12000 47184 6 wbm_a_dat_o[22]
port 84 nsew signal tristate
rlabel metal3 s 11200 47880 12000 48000 6 wbm_a_dat_o[23]
port 85 nsew signal tristate
rlabel metal3 s 11200 48696 12000 48816 6 wbm_a_dat_o[24]
port 86 nsew signal tristate
rlabel metal3 s 11200 49376 12000 49496 6 wbm_a_dat_o[25]
port 87 nsew signal tristate
rlabel metal3 s 11200 50192 12000 50312 6 wbm_a_dat_o[26]
port 88 nsew signal tristate
rlabel metal3 s 11200 51008 12000 51128 6 wbm_a_dat_o[27]
port 89 nsew signal tristate
rlabel metal3 s 11200 51688 12000 51808 6 wbm_a_dat_o[28]
port 90 nsew signal tristate
rlabel metal3 s 11200 52504 12000 52624 6 wbm_a_dat_o[29]
port 91 nsew signal tristate
rlabel metal3 s 11200 31696 12000 31816 6 wbm_a_dat_o[2]
port 92 nsew signal tristate
rlabel metal3 s 11200 53320 12000 53440 6 wbm_a_dat_o[30]
port 93 nsew signal tristate
rlabel metal3 s 11200 54000 12000 54120 6 wbm_a_dat_o[31]
port 94 nsew signal tristate
rlabel metal3 s 11200 32512 12000 32632 6 wbm_a_dat_o[3]
port 95 nsew signal tristate
rlabel metal3 s 11200 33328 12000 33448 6 wbm_a_dat_o[4]
port 96 nsew signal tristate
rlabel metal3 s 11200 34008 12000 34128 6 wbm_a_dat_o[5]
port 97 nsew signal tristate
rlabel metal3 s 11200 34824 12000 34944 6 wbm_a_dat_o[6]
port 98 nsew signal tristate
rlabel metal3 s 11200 35640 12000 35760 6 wbm_a_dat_o[7]
port 99 nsew signal tristate
rlabel metal3 s 11200 36320 12000 36440 6 wbm_a_dat_o[8]
port 100 nsew signal tristate
rlabel metal3 s 11200 37136 12000 37256 6 wbm_a_dat_o[9]
port 101 nsew signal tristate
rlabel metal3 s 11200 2456 12000 2576 6 wbm_a_sel_o[0]
port 102 nsew signal tristate
rlabel metal3 s 11200 3272 12000 3392 6 wbm_a_sel_o[1]
port 103 nsew signal tristate
rlabel metal3 s 11200 4088 12000 4208 6 wbm_a_sel_o[2]
port 104 nsew signal tristate
rlabel metal3 s 11200 4768 12000 4888 6 wbm_a_sel_o[3]
port 105 nsew signal tristate
rlabel metal3 s 11200 280 12000 400 6 wbm_a_stb_o
port 106 nsew signal tristate
rlabel metal3 s 11200 1776 12000 1896 6 wbm_a_we_o
port 107 nsew signal tristate
rlabel metal3 s 0 79160 800 79280 6 wbm_b_ack_i
port 108 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 wbm_b_adr_o[0]
port 109 nsew signal tristate
rlabel metal3 s 0 51552 800 51672 6 wbm_b_adr_o[10]
port 110 nsew signal tristate
rlabel metal3 s 0 47744 800 47864 6 wbm_b_adr_o[1]
port 111 nsew signal tristate
rlabel metal3 s 0 48152 800 48272 6 wbm_b_adr_o[2]
port 112 nsew signal tristate
rlabel metal3 s 0 48560 800 48680 6 wbm_b_adr_o[3]
port 113 nsew signal tristate
rlabel metal3 s 0 48968 800 49088 6 wbm_b_adr_o[4]
port 114 nsew signal tristate
rlabel metal3 s 0 49376 800 49496 6 wbm_b_adr_o[5]
port 115 nsew signal tristate
rlabel metal3 s 0 49784 800 49904 6 wbm_b_adr_o[6]
port 116 nsew signal tristate
rlabel metal3 s 0 50328 800 50448 6 wbm_b_adr_o[7]
port 117 nsew signal tristate
rlabel metal3 s 0 50736 800 50856 6 wbm_b_adr_o[8]
port 118 nsew signal tristate
rlabel metal3 s 0 51144 800 51264 6 wbm_b_adr_o[9]
port 119 nsew signal tristate
rlabel metal3 s 0 44752 800 44872 6 wbm_b_cyc_o
port 120 nsew signal tristate
rlabel metal3 s 0 65560 800 65680 6 wbm_b_dat_i[0]
port 121 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 wbm_b_dat_i[10]
port 122 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 wbm_b_dat_i[11]
port 123 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 wbm_b_dat_i[12]
port 124 nsew signal input
rlabel metal3 s 0 71136 800 71256 6 wbm_b_dat_i[13]
port 125 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 wbm_b_dat_i[14]
port 126 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 wbm_b_dat_i[15]
port 127 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 wbm_b_dat_i[16]
port 128 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 wbm_b_dat_i[17]
port 129 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 wbm_b_dat_i[18]
port 130 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 wbm_b_dat_i[19]
port 131 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 wbm_b_dat_i[1]
port 132 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 wbm_b_dat_i[20]
port 133 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 wbm_b_dat_i[21]
port 134 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 wbm_b_dat_i[22]
port 135 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 wbm_b_dat_i[23]
port 136 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 wbm_b_dat_i[24]
port 137 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 wbm_b_dat_i[25]
port 138 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 wbm_b_dat_i[26]
port 139 nsew signal input
rlabel metal3 s 0 77120 800 77240 6 wbm_b_dat_i[27]
port 140 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 wbm_b_dat_i[28]
port 141 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 wbm_b_dat_i[29]
port 142 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 wbm_b_dat_i[2]
port 143 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 wbm_b_dat_i[30]
port 144 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 wbm_b_dat_i[31]
port 145 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 wbm_b_dat_i[3]
port 146 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 wbm_b_dat_i[4]
port 147 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 wbm_b_dat_i[5]
port 148 nsew signal input
rlabel metal3 s 0 68144 800 68264 6 wbm_b_dat_i[6]
port 149 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 wbm_b_dat_i[7]
port 150 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 wbm_b_dat_i[8]
port 151 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 wbm_b_dat_i[9]
port 152 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 wbm_b_dat_o[0]
port 153 nsew signal tristate
rlabel metal3 s 0 56176 800 56296 6 wbm_b_dat_o[10]
port 154 nsew signal tristate
rlabel metal3 s 0 56584 800 56704 6 wbm_b_dat_o[11]
port 155 nsew signal tristate
rlabel metal3 s 0 57128 800 57248 6 wbm_b_dat_o[12]
port 156 nsew signal tristate
rlabel metal3 s 0 57536 800 57656 6 wbm_b_dat_o[13]
port 157 nsew signal tristate
rlabel metal3 s 0 57944 800 58064 6 wbm_b_dat_o[14]
port 158 nsew signal tristate
rlabel metal3 s 0 58352 800 58472 6 wbm_b_dat_o[15]
port 159 nsew signal tristate
rlabel metal3 s 0 58760 800 58880 6 wbm_b_dat_o[16]
port 160 nsew signal tristate
rlabel metal3 s 0 59168 800 59288 6 wbm_b_dat_o[17]
port 161 nsew signal tristate
rlabel metal3 s 0 59576 800 59696 6 wbm_b_dat_o[18]
port 162 nsew signal tristate
rlabel metal3 s 0 60120 800 60240 6 wbm_b_dat_o[19]
port 163 nsew signal tristate
rlabel metal3 s 0 52368 800 52488 6 wbm_b_dat_o[1]
port 164 nsew signal tristate
rlabel metal3 s 0 60528 800 60648 6 wbm_b_dat_o[20]
port 165 nsew signal tristate
rlabel metal3 s 0 60936 800 61056 6 wbm_b_dat_o[21]
port 166 nsew signal tristate
rlabel metal3 s 0 61344 800 61464 6 wbm_b_dat_o[22]
port 167 nsew signal tristate
rlabel metal3 s 0 61752 800 61872 6 wbm_b_dat_o[23]
port 168 nsew signal tristate
rlabel metal3 s 0 62160 800 62280 6 wbm_b_dat_o[24]
port 169 nsew signal tristate
rlabel metal3 s 0 62568 800 62688 6 wbm_b_dat_o[25]
port 170 nsew signal tristate
rlabel metal3 s 0 62976 800 63096 6 wbm_b_dat_o[26]
port 171 nsew signal tristate
rlabel metal3 s 0 63520 800 63640 6 wbm_b_dat_o[27]
port 172 nsew signal tristate
rlabel metal3 s 0 63928 800 64048 6 wbm_b_dat_o[28]
port 173 nsew signal tristate
rlabel metal3 s 0 64336 800 64456 6 wbm_b_dat_o[29]
port 174 nsew signal tristate
rlabel metal3 s 0 52776 800 52896 6 wbm_b_dat_o[2]
port 175 nsew signal tristate
rlabel metal3 s 0 64744 800 64864 6 wbm_b_dat_o[30]
port 176 nsew signal tristate
rlabel metal3 s 0 65152 800 65272 6 wbm_b_dat_o[31]
port 177 nsew signal tristate
rlabel metal3 s 0 53184 800 53304 6 wbm_b_dat_o[3]
port 178 nsew signal tristate
rlabel metal3 s 0 53728 800 53848 6 wbm_b_dat_o[4]
port 179 nsew signal tristate
rlabel metal3 s 0 54136 800 54256 6 wbm_b_dat_o[5]
port 180 nsew signal tristate
rlabel metal3 s 0 54544 800 54664 6 wbm_b_dat_o[6]
port 181 nsew signal tristate
rlabel metal3 s 0 54952 800 55072 6 wbm_b_dat_o[7]
port 182 nsew signal tristate
rlabel metal3 s 0 55360 800 55480 6 wbm_b_dat_o[8]
port 183 nsew signal tristate
rlabel metal3 s 0 55768 800 55888 6 wbm_b_dat_o[9]
port 184 nsew signal tristate
rlabel metal3 s 0 45568 800 45688 6 wbm_b_sel_o[0]
port 185 nsew signal tristate
rlabel metal3 s 0 45976 800 46096 6 wbm_b_sel_o[1]
port 186 nsew signal tristate
rlabel metal3 s 0 46384 800 46504 6 wbm_b_sel_o[2]
port 187 nsew signal tristate
rlabel metal3 s 0 46928 800 47048 6 wbm_b_sel_o[3]
port 188 nsew signal tristate
rlabel metal3 s 0 44344 800 44464 6 wbm_b_stb_o
port 189 nsew signal tristate
rlabel metal3 s 0 45160 800 45280 6 wbm_b_we_o
port 190 nsew signal tristate
rlabel metal3 s 0 43936 800 44056 6 wbs_ack_o
port 191 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 wbs_adr_i[0]
port 192 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 wbs_adr_i[10]
port 193 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 wbs_adr_i[11]
port 194 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 wbs_adr_i[12]
port 195 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 wbs_adr_i[13]
port 196 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 wbs_adr_i[14]
port 197 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 wbs_adr_i[15]
port 198 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 wbs_adr_i[16]
port 199 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 wbs_adr_i[17]
port 200 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 wbs_adr_i[18]
port 201 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 wbs_adr_i[19]
port 202 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 wbs_adr_i[1]
port 203 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_adr_i[20]
port 204 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 wbs_adr_i[21]
port 205 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 wbs_adr_i[22]
port 206 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 wbs_adr_i[23]
port 207 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 wbs_adr_i[24]
port 208 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 wbs_adr_i[25]
port 209 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 wbs_adr_i[26]
port 210 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 wbs_adr_i[27]
port 211 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 wbs_adr_i[28]
port 212 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 wbs_adr_i[29]
port 213 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 wbs_adr_i[2]
port 214 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 wbs_adr_i[30]
port 215 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 wbs_adr_i[31]
port 216 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 wbs_adr_i[3]
port 217 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 wbs_adr_i[4]
port 218 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 wbs_adr_i[5]
port 219 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 wbs_adr_i[6]
port 220 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 wbs_adr_i[7]
port 221 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 wbs_adr_i[8]
port 222 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 wbs_adr_i[9]
port 223 nsew signal input
rlabel metal3 s 0 552 800 672 6 wbs_cyc_i
port 224 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 wbs_dat_i[0]
port 225 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 wbs_dat_i[10]
port 226 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 wbs_dat_i[11]
port 227 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 wbs_dat_i[12]
port 228 nsew signal input
rlabel metal3 s 0 22176 800 22296 6 wbs_dat_i[13]
port 229 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 wbs_dat_i[14]
port 230 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 wbs_dat_i[15]
port 231 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 wbs_dat_i[16]
port 232 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 wbs_dat_i[17]
port 233 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 wbs_dat_i[18]
port 234 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 wbs_dat_i[19]
port 235 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 wbs_dat_i[1]
port 236 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 wbs_dat_i[20]
port 237 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 wbs_dat_i[21]
port 238 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 wbs_dat_i[22]
port 239 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 wbs_dat_i[23]
port 240 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 wbs_dat_i[24]
port 241 nsew signal input
rlabel metal3 s 0 27344 800 27464 6 wbs_dat_i[25]
port 242 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 wbs_dat_i[26]
port 243 nsew signal input
rlabel metal3 s 0 28160 800 28280 6 wbs_dat_i[27]
port 244 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 wbs_dat_i[28]
port 245 nsew signal input
rlabel metal3 s 0 28976 800 29096 6 wbs_dat_i[29]
port 246 nsew signal input
rlabel metal3 s 0 17552 800 17672 6 wbs_dat_i[2]
port 247 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 wbs_dat_i[30]
port 248 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 wbs_dat_i[31]
port 249 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 wbs_dat_i[3]
port 250 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 wbs_dat_i[4]
port 251 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 wbs_dat_i[5]
port 252 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 wbs_dat_i[6]
port 253 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 wbs_dat_i[7]
port 254 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 wbs_dat_i[8]
port 255 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 wbs_dat_i[9]
port 256 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 wbs_dat_o[0]
port 257 nsew signal tristate
rlabel metal3 s 0 34552 800 34672 6 wbs_dat_o[10]
port 258 nsew signal tristate
rlabel metal3 s 0 34960 800 35080 6 wbs_dat_o[11]
port 259 nsew signal tristate
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_o[12]
port 260 nsew signal tristate
rlabel metal3 s 0 35776 800 35896 6 wbs_dat_o[13]
port 261 nsew signal tristate
rlabel metal3 s 0 36184 800 36304 6 wbs_dat_o[14]
port 262 nsew signal tristate
rlabel metal3 s 0 36592 800 36712 6 wbs_dat_o[15]
port 263 nsew signal tristate
rlabel metal3 s 0 37136 800 37256 6 wbs_dat_o[16]
port 264 nsew signal tristate
rlabel metal3 s 0 37544 800 37664 6 wbs_dat_o[17]
port 265 nsew signal tristate
rlabel metal3 s 0 37952 800 38072 6 wbs_dat_o[18]
port 266 nsew signal tristate
rlabel metal3 s 0 38360 800 38480 6 wbs_dat_o[19]
port 267 nsew signal tristate
rlabel metal3 s 0 30744 800 30864 6 wbs_dat_o[1]
port 268 nsew signal tristate
rlabel metal3 s 0 38768 800 38888 6 wbs_dat_o[20]
port 269 nsew signal tristate
rlabel metal3 s 0 39176 800 39296 6 wbs_dat_o[21]
port 270 nsew signal tristate
rlabel metal3 s 0 39584 800 39704 6 wbs_dat_o[22]
port 271 nsew signal tristate
rlabel metal3 s 0 40128 800 40248 6 wbs_dat_o[23]
port 272 nsew signal tristate
rlabel metal3 s 0 40536 800 40656 6 wbs_dat_o[24]
port 273 nsew signal tristate
rlabel metal3 s 0 40944 800 41064 6 wbs_dat_o[25]
port 274 nsew signal tristate
rlabel metal3 s 0 41352 800 41472 6 wbs_dat_o[26]
port 275 nsew signal tristate
rlabel metal3 s 0 41760 800 41880 6 wbs_dat_o[27]
port 276 nsew signal tristate
rlabel metal3 s 0 42168 800 42288 6 wbs_dat_o[28]
port 277 nsew signal tristate
rlabel metal3 s 0 42576 800 42696 6 wbs_dat_o[29]
port 278 nsew signal tristate
rlabel metal3 s 0 31152 800 31272 6 wbs_dat_o[2]
port 279 nsew signal tristate
rlabel metal3 s 0 42984 800 43104 6 wbs_dat_o[30]
port 280 nsew signal tristate
rlabel metal3 s 0 43528 800 43648 6 wbs_dat_o[31]
port 281 nsew signal tristate
rlabel metal3 s 0 31560 800 31680 6 wbs_dat_o[3]
port 282 nsew signal tristate
rlabel metal3 s 0 31968 800 32088 6 wbs_dat_o[4]
port 283 nsew signal tristate
rlabel metal3 s 0 32376 800 32496 6 wbs_dat_o[5]
port 284 nsew signal tristate
rlabel metal3 s 0 32784 800 32904 6 wbs_dat_o[6]
port 285 nsew signal tristate
rlabel metal3 s 0 33192 800 33312 6 wbs_dat_o[7]
port 286 nsew signal tristate
rlabel metal3 s 0 33736 800 33856 6 wbs_dat_o[8]
port 287 nsew signal tristate
rlabel metal3 s 0 34144 800 34264 6 wbs_dat_o[9]
port 288 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 wbs_sel_i[0]
port 289 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 wbs_sel_i[1]
port 290 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wbs_sel_i[2]
port 291 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 wbs_sel_i[3]
port 292 nsew signal input
rlabel metal3 s 0 144 800 264 6 wbs_stb_i
port 293 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wbs_we_i
port 294 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12000 80000
<< end >>
